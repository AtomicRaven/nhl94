GST@�                                                            \     �                                               R���      �  ��  5         ���2�������J�������������������        �g      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"��   " `  J  jF��     �j  
 ���
��
��    "�j��" " ��
  �                                                                               ����������������������������������      ��    bb? QQ0 5 118 44               		 


     
               ��� 4    �                 nn ))
         88:�����������������������������������������������������������������������������������������������������������������������������=  0b  4  11                                         �  �  �  �                  F  
          = �����������������������������������������������������������������������������                                ��  �   �  ��   @  #   �   �                                                                                '     )n)n
  
F    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE ; �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    	��AE=k�>�/������M��C�T@E=@R<ED_�Z3�T0 k� �t6�x6	E1 4#Q&�1D"3Q  �9    � !�;	��AE=c�>�/������M�C�H@E=8Q�4ED_�Z3�T0 k� ��8��8	E1 4#Q&�1D"3Q  ��?    � !�>	��AE=[�>�/������M�C�@AE=8Q�0DD_�Z3�T0 k� ��:��:	E1 4#Q&�1D"3Q  ��?    � !�A	��AE=O�>�.��������E�4AE=$Q�$CD_�Z3�T0 k� ��>��>	E1 4#Q&�1D"3Q  ��?    � !�D	ͼAE=K�>�.�|�����ۖE�,ACMQ�CE_�Z3�T0 k� ��@��@	E1 4#Q&�1D"3Q  ��?    � !�G	͸AE=C�^�.�t�����זE�$ACMQ�CE_�Z3�T0 k� ��B��B	E1 4#Q&�1D"3Q  ��?    � !�J	ͰAE-;�^�-p�����ӗE�$ACMQ�BE_�Z3�T0 k� ��E��E	E1 4#Q&�1D"3Q  ��?    � "�H�AE-/�^p-d����ǘE�ACM Q�AE_xZ3�T0 k� �E�E	E1 4#Q&�1D"3Q  ��8    � #�G�@E-+�^h,`�w�!����E�AE<�Q�AE_tZ3�T0 k� � B�B	E1 4#Q&�1D"3Q  ��8    � $�F�@E-'�^`,\�o�!����E�AE<�Q��@I�lZ3�T0 k� ��@��@	E1 4#Q&�1D"3Q  ��8    � %�E�@E-#�^X,X�g�!����E��AE<�Q	�@I�dZ3�T0 k� ��?��?	E1 4#Q&�1D"3Q  ��8    � &�D�@E-�^H+P�W�!����E��AE<�Q	�?I�XZ3�T0 k� ��=��=	E1 4#Q&�1D"3Q  ��8    � '�C�?E-�^@+L�O�!����E��AE<�Q	�?I�PZ3�T0 k� ��=��=	E1 4#Q&�1D"3Q  ��8    � (�B�x?E-��8+H�G�!����E��@E<�P	�>I�HZ3�T0 k� ��<��<	E1 4#Q&�1D"3Q  ��8    � (�A�p>E-��,+D�?�!����E��@E<�P	�>I�D	Z3�T0 k� ��<��<	E1 4#Q&�1D"3Q  ��8    � (�@�l>E-��$*@�7�!����E��@E<�P	�=I�<	Z3�T0 k� ��;��;	E1 4#Q&�1D"3Q  ��8    � (�?�\=E��*�<	�'�!����E��@E<�O	�=I�4	Z3�T0 k� ��:��:	E1 4#Q&�1D"3Q  ��8    � (�>�T<E���*�8����{�E��?E<�O	�<I�,	Z3�T0 k� ��:��:	E1 4#Q&�1D"3Q  ��8    � (�=�P<E���)�8����w�E��?E,�O	�<E�(	Z3�T0 k� ��;��;	E1 4#Q&�1D"3Q  ��8    � (�<�H;E����)�4����o�E��?E,�N	�;E� 
Z3�T0 k� ��;��;	E1 4#Q&�1D"3Q  ��8    � (�;�<9E����(�4�����c�E�?E,�M	�;E�
Z3�T0 k� ��;��;	E1 4#Q&�1D"3Q  ��8    � (�:�48E����(�0�����[�E�?E,�M	�:E�Z3�T0 k� ��<��<	E1 4#Q&�1D"3Q  ��8    � (�9�,8E����(�0�����S�E��?E,|M	�:E�Z3�T0 k� ��<��<	E1 4#Q&�1D"3Q  ��8    � (�8�(7E����'�0�����K�E��?E,tM	�:E� Z3�T0 k� ��<��<	E1 4#Q&�1D"3Q  ��8    � (�8� 5E�����'�0�����C�E��?E,pL	�9E��Z3�T0 k� �x<�|<	E1 4#Q&�1D"3Q  ��8    � (�8�3E����&�0 �����7�E��?E,`L	�9E��Z3�T0 k� �l;�p;	E1 4#Q&�1D"3Q  ��8    � (�8�2E����&�3����!��/�E��>@|\L	�8E��Z3�T0 k� �l9�p9	E1 4#Q&�1D"3Q  ��8    � (�81E����%�3����!��'�E��>@|TK	�8E��Z3�T0 k� �h7�l7	E1 4#Q&�1D"3Q  ��8    � (�80E����%�3����!���E��>@|PK�7E��Z3�T0 k� �h5�l5	E1 4#Q&�1D"3Q  ��8    � (�8�-E�����$�3����!���E�x>@|HJ�7E��Z3�T0 k� �`4�d4	E1 4#Q&�1D"3Q  ��8    � (�8�,D�����#�3����",��E�x>@|@J�6E��Z3�T0 k� �\3�`3	E1 4#Q&�1D"3Q  ��8    � (�8�*D����|#�3����",��E�t=@|<J�6E�Z3�T0 k� �X3�\3	E1 4#Q&�1D"3Q  ��8    � (�8�)D����t"�3����",���E�p=@|8J�5E�Z3�T0 k� �T3�X3	E1 4#Q&�1D"3Q  ��8    � (�8�(D����p!�7����",��Fh=@|0I�5E�Z3�T0 k� �L2�P2	E1 4#Q&�1D"3Q  ��8    � (�8�%D���`�7���",��F`=@|(I|3E�Z3�T0 k� �D1�H1	E1 4#Q&�1D"3Q  ��8    � (�8�#E���X�;��w���߼F\>E,$H�|3E��Z3�T0 k� �<3�@3	E1 4#Q&�1D"3Q  ��8    � (�8�"E���P;��o��	�׼FX>E, H�x2E��Z3�T0 k� �44�84	E1 4#Q&�1D"3Q  ��8    � (�8� E���H?�	}k��	�ӽFT>E,G�x2E��Z3�T0 k� �05�45	E1 4#Q&�1D"3Q  ��8    � (�8��E���<C�	}[��	�ÿFT>E,F�t1E�|Z3�T0 k� �(5�,5	E1 4#Q&�1D"3Q  ��8    � (�8��E���4C�	}W��	���D�P>E,F�t0E�xZ3�T0 k� �$5�(5	E1 4#Q&�1D"3Q  ��8    � (�8��E��,G�	}O��	���D�L>E,E�t0E�pZ3�T0 k� � 5�$5	E1 4#Q&�1D"3Q  ��8    � (�8��E��(G�	�K��	���D�L>E,D�p/E�hZ3�T0 k� �4� 4	E1 4#Q&�1D"3Q  ��8    � (�8��E�'�O�	�?��	���D�H?EC�p/E�\ Z3�T0 k� �8�8	E1 4#Q&�1D"3Q  ��8    � (�8��B�+�O�	�;��	���D�H?EB�p.E�X!Z3�T0 k� �;�;	E1 4#Q&�1D"3Q  ��8    � (�8��B�/�S�	�3��	���D�D@E B �p.E�P"Z3�T0 k� �>�>	E1 4#Q&�1D"3Q  ��8    � (�8��B�3�W�	}/��	���D�D@E A �p.E�L$Z3�T0 k� �?�?	E1 4#Q&�1D"3Q  ��8    � (�8��B�7�[�	}+��	���D�DAE�A �p.FD%Z3�T0 k� �@�@	E1 4#Q&�1D"3Q  ��8    � (�8��I?�_�	}��	���D�DBE�@ �p.F8(Z3�T0 k� �@�@	E1 4#Q&�1D"3Q  ��8 
   � (�8��IC�c�	}��	���D�DBE�? �p.F4)Z3�T0 k� �A�A	E1 4#Q&�1D"3Q  ��8 
   � (�8��IG�g�M��	���D�DCE��>l.F0*Z3�T0 k� �E�E	E1 4#Q&�1D"3Q  ��8 
   � (�8��
IG��k�M��	���D�DDE��>p.F,,Z3�T0 k� �H�H	E1 4#Q&�1D"3Q  ��8 
   � (�8��I-O���p M��	�{�D�DEE��=p.F$/Z3�T0 k� �J�J	E1 4#Q&�1D"3Q  ��8 
   � (�8��I-S�� �tM��	�{�D�DFE��=p.F 0Z3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 
   � (�8��I-S����xM��	�w�FDGB[�=t.F2Z3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 
   � (�8��I-W����x=��	�s�FHHB[�<[t.F3Z3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 
   � (�8��I-W����x=��	�s�FHHB[�<[t.F5Z3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 
   � (�8��I[����|<���	�o�FHIB[�<[t.F6Z3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 
   � (�8��I_����|<���	�k�FLKB\ <[x.E�:Z3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 
   � (�8��I_����|<���	�g�E�LLB\ <[x.E�;Z3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 	   � (�8��I_�����<���	�g�E�PMB\ <[x.E�=Z3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 	   � (�8��I-c�����<���	�g�E�TNB\<[x.E�>Z3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 	   � (�8��I-c�����,���	�c�E�TOB\<[x.E�?Z3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 	   � (�8��I-c�����,���	�c�E�XPB\<[|.B�AZ3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 	   � (�8�I-c���̀,���	�c�B�\QBl=�|/B� BZ3�T0 k� �K�K	E1 4#Q&�1D"3Q  ��8 	   � (�8�I-g���̀,���	�_�B�`RBl=�|/B� DZ3�T0 k� �K� K	E1 4#Q&�1D"3Q  ��8 	   � (�8�Ig�� ̀
 l���	�_�B�dSBl>�|/B� FZ3�T0 k� � K�$K	E1 4#Q&�1D"3Q  ��8 	   � (�8�Ig��̀ l���L[�B�hTBl>��.B� HZ3�T0 k� �$L�(L	E1 4#Q&�1D"3Q  ��8 	   � (�8�Ig���� l���L[�B�lUBl>;�.B� IZ3�T0 k� �(L�,L	E1 4#Q&�1D"3Q  ��8 	   � (�8�Ig���� l���LW�B�tVBl?;�.B� JZ3�T0 k� �(L�,L	E1 4#Q&�1D"3Q  ��8 	   � (�8�Ig���| l���LW�B�xWBl?;�.B� LZ3�T0 k� �,M�0M	E1 4#Q&�1D"3Q  ��8 	   � (�8�@g���| l���LS�B�|WF @;�.B�MZ3�T0 k� �8M�<M	E1 4#Q&�1D"3Q  ��8 	   � (�8��@g���| l���<S�B��XF$@;�-B�NZ3�T0 k� �DN�HN	E1 4#Q&�1D"3Q  ��8 	   � (�8��@g��<| l���<O�B��ZF,A��-B�QZ3�T0 k� �PO�TO	E1 4#Q&�1D"3Q  ��8 	   � (�8��	@g��<x l���<O�B��ZF0B��,B�RZ3�T0 k� �XP�\P	E1 4#Q&�1D"3Q  ��8    � (�8��	@g��<x l���<K�B��[E�4B��,B�SZ3�T0 k� �XL�\L	E1 4#Q&�1D"3Q  ��8    � (�8��
BMg�� <x l���<K�B��\E�8C��+B�TZ3�T0 k� �XJ�\J	E1 4#Q&�1D"3Q  ��8    � (�8��BMg��$<x l���,G�B��]E�<C��+B�UZ3�T0 k� �XH�\H	E1 4#Q&�1D"3Q  ��8    � (�8��BMg��0<t ����,C�E��_E�DD��*E�XZ3�T0 k� �`G�dG	E1 4#Q&�1D"3Q  ��8    � (�8��BMg��4<t ����,C�E��`E�LE��)E�YZ3�T0 k� �dG�hG	E1 4#Q&�1D"3Q  ��8    � (�8��BMg��8<t ����,C�E��aE�PE��(E�ZZ3�T0 k� �hB�lB	E1 4#Q&�1D"3Q  ��8    � (�8��BMg��<<t ����,C�E��bE�TF��(E� [Z3�T0 k� �p?�t?	E1 4#Q&�1D"3Q  ��8    � (�8��BMg��@<t  ����,C�E��cE�\F��'E�$\Z3�T0 k� �t=�x=	E1 4#Q&�1D"3Q  ��8    � (�8��BMg��L<p# ����,?�D��fE�hF�%E�,^Z3�T0 k� ��;��;	E1 4#Q&�1D"3Q  ��8    � (�8��BMg��P<p% �����?�D��gE�lG�&E�0_Z3�T0 k� ��:��:	E1 4#Q&�1D"3Q  ��8    � (�8<�BMg��X,p& �����?�D��hE�tG�&E�4`Z3�T0 k� ��9��9	E1 4#Q&�1D"3Q  ��8    � (�8<�A�g��\,p( �����?�D��iE�xG�&E�8aZ3�T0 k� ��9��9	E1 4#Q&�1D"3Q  ��8    � (�8<�A�g��h,p+ �����C�I��kE��G��'E�@cZ3�T0 k� ��8��8	E1 4#Q&�1D"3Q  ��8    � (�8<�A�g��l,p- ����,C�I��lE��G��'E�DdZ3�T0 k� ��8��8	E1 4#Q&�1D"3Q  �8    � (�8<�A�g��t,p/L���,C�I��lE��G��'E�LeZ3�T0 k� ��8��8	E1 4#Q&�1D"3Q  �8    � (�8= D�g��x,p0L���,C�I��mE��G��'E�PfZ3�T0 k� ��7��7	E1 4#Q&�1D"3Q  ��8    � (�8= D�g���,t4L���,G�JoE��F��(E�XgZ3�T0 k� ��7��7	E1 4#Q&�1D"3Q  ��8    � (�8="D�g���,t6L���,G�JpE��F �(E�\hZ3�T0 k� ��7��7	E1 4#Q&�1D"3Q  ��8    � (�8M#D�g����x9L��� lG�JqE��F �(E�`iZ3�T0 k� ��6��6	E1 4#Q&�1D"3Q  ��8    � (�8M%D�g����<L��� lG�JqE��E �)E�hjZ3�T0 k� ��6��6	E1 4#Q&�1D"3Q  ��8    � (�8M'D�g����<L��� lG�JrE��E �)E�ljZ3�T0 k� ��4��4	E1 4#Q&�1D"3Q  ��8    � (�8M*D�g����AL��� lK�BM$tE��E �)@ntlZ3�T0 k� ��2��2	E1 4#Q&�1D"3Q  ��8    � (�8M,D�g���,�CL��� lK�BM(uE��D �)@nxmZ3�T0 k� ��1��1	E1 4#Q&�1D"3Q  ��8    � (�8M.D�g���,�EL��� lK�BM,uE��D �*@n|mZ3�T0 k� ��0��0	E1 4#Q&�1D"3Q  ��8    � (�8�0D�g���,�G\��� lK�BM0vE��D �*@n�nZ3�T0 k� ��.��.	E1 4#Q&�1D"3Q  ��8    � (�8�2D�g���,�I\� � lK�BM4wE��C �*@n�oZ3�T0 k� ��-��-	E1 4#Q&�1D"3Q  ��8    � (�8�4D�g���,�K\�� lK�BM8wE��C �*@n�oZ3�T0 k� ��*��*	E1 4#Q&�1D"3Q  �8    � (�8�4D�g���,�L\�� lO�BM<xG C �*@n�pZ3�T0 k� ��'��'	E1 4#Q&�1D"3Q  ��?    � (�8�4D�g���,�N\�� lO�BM@yGD �+@n�qZ3�T0 k� ��$��$	E1 4#Q&�1D"3Q  ��?    � (�8�$6D�g���!,�R\�� lO�BMHxGD �+@n�rZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��?    � (�8�,7D�g���",�T\�� lO�BMLxGE �+@n�sZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��D    � (�8�07D�g���#,�V<���O�BMPxGE �+@n�sZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��D    � (�8�48D�g���%,�W<���S�BMTxGF �,@n�tZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��D    � (�8�89D�g���&,�Y<���S�BMXwGG �,@n�uZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��D    � (�8�@;D�g���),�]<�
� �S�BM`wGG �,@n�vZ3� T0 k� ����	E1 4#Q&�1D"3Q  ��D    � (�8�D<D�g���*,�^,��  lS�BMdwGH �,@n�vZ3� T0 k� ����	E1 4#Q&�1D"3Q  ��D    � (�8�H<D�g���,,�`,��  lS�BMhvG-I �-@n�wZ3� T0 k� ����	E1 4#Q&�1D"3Q  ��D    � (�8�L=D�g�� -,�a,��  lS�BMhvG- I �-@n�xbs� T0 k� ��� 	E1 4#Q&�1D"3Q  ��D    � (�8�P>D�g��/,�c,��  lW�BMlvG-$J �-@n�xbs��T0 k� � �	E1 4#Q&�1D"3Q  ��D    � (�8�X@D�g��2,�f- �$ lW�BMtvG-$J �-@n�ybs��T0 k� ��	E1 4#Q&�1D"3Q  ��D    � (�8�X@D�g��3,�h- �$ lW�BMxuG-(K �-@n�zbs��T0 k� �!�!	E1 4#Q&�1D"3Q  ��D    � (�8�\AD�g��5,�i �$ lW�BM|uG-,L �.@n�zbs��T0 k� ��	E1 4#Q&�1D"3Q  ��D    � (�8�`BD�g��6,�k�$ lW�BM|uG-,M �.@n�{bs��T0 k� ��	E1 4#Q&�1D"3Q  ��D    � (�8�dCD�g��8,�l�$ lW�BM�uG-0N �.@n�|bs��T0 k� ��	E1 4#Q&�1D"3Q  ��D    � (�8�dDD�g��9,�n�( lW�BM�uG-4O �.@n�|bs��T0 k� ��	E1 4#Q&�1D"3Q  ��D    � (�8�dDD�g��<,�q�( l[�BM�tG-8P �.@n�}bs� T0 k� ��	E1 4#Q&�1D"3Q  ��D    � (�8�hDD�g��>,�r�( l[�BM�tG-8Q �.@n�~Z3� T0 k� ��	E1 4#Q&�1D"3Q  ��D    � (�8�hED�g��?,�t�( l[�BM�tG-<R �/@n�~Z4 T0 k� �� 	E1 4#Q&�1D"3Q  ��D   � (�8�lFD�g��A�u�( l[�BM�tG-<S �/@n�Z4T0 k� � �$	E1 4#Q&�1D"3Q  ��D    � (�8�lGD�g��B�w�, l[�BM�sG-@T �/@n�Z4T0 k� �$�(	E1 4#Q&�1D"3Q  ��D    � (�8�lHD�g��E�y  �, l[�BM�sG-DV �/@n�Z4T0 k� �(�,	E1 4#Q&�1D"3Q  ��D    � (�8�lIL]g��G�{$"�, l[�BM�sG-DV �/@n�Z4T0 k� �,�0	E1 4#Q&�1D"3Q  ��D    � (�8�pJL]g��H�|(#�, l_�BM�sG-DW �/@n�Z4T0 k� �0�4	E1 4#Q&�1D"3Q  ��D    � (�8�pJL]g��I },$�, l_�BM�sG-DX �0@n�Z4T0 k� �4�8	E1 4#Q&�1D"3Q  ��D    � (�8�pKL]g��K0%�, l_�BM�r@�HY �0@n�Z4T0 k� �8�<	E1 4#Q&�1D"3Q  ��D    � (�8�pKL]g��L�4&�0 l\ BM�r@�HZ �0@n�Z4T0 k� �<�@	E1 4#Q&�1D"3Q   �D    � (�8�pKL]g��M�4'�0 l\ BM�r@�L[ �0@n�b�T0 k� �@ �D 	E1 4#Q&�1D"3Q  ��D    � (�8�pLL]g��P�<)�0 l\BM�r@�L\ �0@n�~b�T0 k� �D"�H"	E1 4#Q&�1D"3Q  ��D    � (�8�pML]g��Q�  @)�0 l\BM�r@�P] �0@o ~b�T0 k� �X#�\#	E1 4#Q&�1D"3Q  ��D    � (�8�lML]g��R�$~ D*�0 l\BM�q@�P^ �1@o~b�T0 k� �h$�l$	E1 4#Q&�1D"3Q  ��D    � (�8�lNL]g��T�(~ D+�0 l\BM�q@�P_ �1@o}b�T0 k� �t%�x%	E1 4#Q&�1D"3Q  ��D    � (�8�lNL]g�� U�0} H,�0 l`BM�q@�T` �1@o}b�T0 k� �|&��&	E1 4#Q&�1D"3Q  ��D    � (�8�hOL]g���V�4} L-�4 l`BM�q@�Ta �1@o}b�T0 k� ��&��&	E1 4#Q&�1D"3Q  ��D    � (�8�dOL]g���W�<| P.�4 l`BM�q@�Ta �1@o}b�T0 k� ��'��'	E1 4#Q&�1D"3Q  ��D    � (�8�dPLmg���X�@{ P/�4 l`BM�q@�Xb �1@o|b�	T0 k� ��(��(	E1 4#Q&�1D"3Q  ��D    � (�8�`PLmg���Y�H{ T0�4 l`BM�q@�Xc �1@o|b�	T0 k� ��)��)	E1 4#Q&�1D"3Q  ��D   � (�8�\QLmg���\�Pz X1�4 l`BM�p@�\d �1@o|Z4
T0 k� ��+��+	E1 4#Q&�1D"3Q  ��D    � (�8m\RLmg���]�Xy \2�4 l`BM�p@�\e �2@o|Z4
T0 k� ��,��,	E1 4#Q&�1D"3Q  ��D    � (�8mXSLmg���^}\x `3�4 l`BM�p@�\f �2@o{Z4
T0 k� ��,��,	E1 4#Q&�1D"3Q  ��D    � (�8mXSLmg���_}dw `4�4 l`BM�p@�`g �2@o{Z4T0 k� ��-��-	E1 4#Q&�1D"3Q  ��D    � (�8mXTLmg���`}hw d5�8 l`	BM�p@�`g �2@o{Z4T0 k� ��.��.	E1 4#Q&�1D"3Q  ��D    � (�8mTULmg���`}hw h5�8 ld	BM�p@�`g �2@o {Z4T0 k� ��/��/	E1 4#Q&�1D"3Q  ��D    � (�8}TVLmd ��`}lw h6�8 ld
BM�p@�`g �2@o {Z4T0 k� ��0��0	E1 4#Q&�1D"3Q  ��D    � (�8}TWLmd�a}xw p8�8 ld
BM�qE=dg �2@o$zZ4T0 k� ��1��1	E1 4#Q&�1D"3Q  ��D    � (�8}TWLmd�b}�w p8�8 ldBM�rE=dg �2@o(zZ4T0 k� ��2��2	E1 4#Q&�1D"3Q  ��D    � (�8}TWLmd�b}�w t9�8 ldBM�rE=hg �3@o(zZ4T0 k� ��3��3	E1 4#Q&�1D"3Q  ��D    � (�8}TWLmd�b}�w t:�8 ldBM�rE=lh �3@o,zZ4T0 k� ��3��3	E1 4#Q&�1D"3Q  ��D    � (�8}PWLmd	�c}�v x;�8 ldBM�sE=lh �3@o,zZ4T0 k� ��4��4	E1 4#Q&�1D"3Q  ��D    � (�8�PXLmd
�c}�v |;�8 ldBM�s@mph �3@o,zZ4T0 k� ��5��5	E1 4#Q&�1D"3Q  ��D    � (�8�PXLmd�c}�v |<�8 ldBM�s@mph �3@o0yZ4T0 k� ��6��6	E1 4#Q&�1D"3Q  ��D    � (�8�LZLmd�c}�v �=�8 lhBM�t@mli �3@o4yZ4T0 k� ��7��7	E1 4#Q&�1D"3Q  ��D    � (�8�H[Lmd�c��v �>�8 lhBM�t@mli �3@o4yZ4T0 k� ��8��8	E1 4#Q&�1D"3Q  ��D    � (�8�H[Lmd�c��v �?�8 lhBM�t@mhj �3@o8yZ4T0 k� ��8��8	E1 4#Q&�1D"3Q  ��D    � (�8�D\Lmd�d��v �?�8 lhBM�uB�hj �3@o8yZ4T0 k� ��9��9	E1 4#Q&�1D"3Q  ��D    � (�8�D\Lmd�d��v �@�8 lhBM�uB�hj �3@o8xZ4T0 k� ��:��:	E1 4#Q&�1D"3Q  ��D    � (�8@]Lmd�d��v �A�8 llBM�uB�hk �4@o<xZ4T0 k� ��:��:	E1 4#Q&�1D"3Q  ��D    � (�8<^Lmd�d��w �A�8 llBM�uB�hk �4@o<xZ4T0 k� ��;��;	E1 4#Q&�1D"3Q  ��D    � (�88^Lmd�d��w �B�8 llBN vB�hk �4@o@xZ4T0 k� ��;��;	E1 4#Q&�1D"3Q  ��D    � (�84_Lmd�c��w �B�8 llBNvE-dl �4@o@xZ4T0 k� ��<��<	E1 4#Q&�1D"3Q  ��D    � (�80`Lmd�c��w �C�8 llBNvE-dl �4@o@xZ4T0 k� ��=��=	E1 4#Q&�1D"3Q  ��D    � (�8,`Lmd�c��w �D�8 llBNvE-dl �4@oDxZ4T0 k� ��=��=	E1 4#Q&�1D"3Q  ��D    � (�8(aLmd�c��w �D�8 llBNwE-dm �4@oDwZ4T0 k� ��>��>	E1 4#Q&�1D"3Q  ��D    � (�8$bLmd�c��w �E�8 lpBNwE-`m �4@oDwZ4T0 k� ��>��>	E1 4#Q&�1D"3Q  ��D    � (�8 bLmd�c��w �E�8 lpBNwE-`m �4@oHwZ4T0 k� ��?��?	E1 4#Q&�1D"3Q  ��D    � (�8cLmd =�c��w �F�8 lpBNwE-`n �4@oHwZ4T0 k� ��?��?	E1 4#Q&�1D"3Q  ��D    � (�8-dLmd!=�c��w �F�8 lpBNx@m`n �4@oLwZ4T0 k� ��@��@	E1 4#Q&�1D"3Q  ��D    � (�8-dLmd"=�c��w �G�8 lpBNx@m\n �4@oLwZ4T0 k� ��A��A	E1 4#Q&�1D"3Q  ��D    � (�8-eLmd#=�c��w �G�8 lpBNx@m\o �4@oLwZ4T0 k� ��A��A	E1 4#Q&�1D"3Q  ��D    � (�8-eLmd$=�c��w �H�8 lpBN x@m\o �5@oPwZ4T0 k� ��B��B	E1 4#Q&�1D"3Q  ��D    � (�8-fLmd%=�d��w �H�8 ltBN x@m\o �5@oPvZ4T0 k� ��B��B	E1 4#Q&�1D"3Q  ��D    � (�8 fLmd&=�d��w �I�8 ltBN$y@mXp �5@oPvZ4T0 k� ��C��C	E1 4#Q&�1D"3Q  ��D    � (�8�fLmd'=�d��w �I�8 ltBN$x@mXp �5@oPvZ4T0 k� ��C��C	E1 4#Q&�1D"3Q  ��D    � (�8�gL]d(=�d��w �J�8 ltBN(x@mXp �5@oTvZ4T0 k� ��D��D	E1 4#Q&�1D"3Q  ��D    � (�8�gL]d)=�d��w �J�8 ltBN,x@mXq �5@oTvZ4T0 k� ��D��D	E1 4#Q&�1D"3Q  ��D    � (�8�hL]d*=�d��w �K�8 ltBN,x@mTq �5@oTvZ4T0 k� ��E��E	E1 4#Q&�1D"3Q  ��D   � (�8�hL]d+=�d��w �K�8 ltBN0w@mTq �5@oXvZ4T0 k� ��E��E	E1 4#Q&�1D"3Q  ��D    � (�8�hL]d,=�d��w �L�8 ltBN0w@mTq �5@oXvZ4T0 k� ��E��E	E1 4#Q&�1D"3Q  ��D    � (�8��iL]d,M�d��w��L�8 ltBN4w@mTr �5@oXvZ4T0 k� ��G��G	E1 4#Q&�1D"3Q  ��D    � (�8��iD�d-M�d��w��M�8 lxBN4w@mTr �5@o\uZ4T0 k� ��H��H	E1 4#Q&�1D"3Q  ��D   � (�8��iD�d.M�d��w��M�8 lxBN8v@mPr �5@o\uZ4T0 k� ��J��J	E1 4#Q&�1D"3Q  ��D    � (�8��iD�d0M�d��x��N�8 lxBN<v@mPs �5@o\uZ4T0 k� ��K��K	E1 4#Q&�1D"3Q  ��D    � (�8��jD�d1M�d��x��N�8 lxBN<v@mPs �5@o\uZ4 T0 k� ��L��L	E1 4#Q&�1D"3Q  ��D    � (�8��jD�d2M�d��x��N�8 lxBN@v@mPs �5@o`uZ4 T0 k� ��L��L	E1 4#Q&�1D"3Q  ��D    � (�8��jEmd3M�d��x��O�8 lxBN@u@mPs �5@o`uZ4 T0 k� ��M��M	E1 4#Q&�1D"3Q  ��D    � (�8L�jEmd4M�d��x��O�8 lxBNDu@mLt �6@o`uZ4 T0 k� ��M��M	E1 4#Q&�1D"3Q  ��D    � (�8L�jEmd5M|d��x��P�8 lxBNDu@mLt �6@o`uZ4 T0 k� ��M��M	E1 4#Q&�1D"3Q  ��D    � (�8L�jEm`7M|d��x��P�8 lxBNHu@mLt �6@oduZ4 T0 k� ��N��N	E1 4#Q&�1D"3Q  ��D    � (�8L�iEm`8M|d��x��P�8 l|BNHu@mLt �6@oduZ4 T0 k� ��N��N	E1 4#Q&�1D"3Q  ��D    � (�8L�iEm`9M|d��x��Q�8 l|BNLt@mLu �6@oduZ4 T0 k� ��N��N	E1 4#Q&�1D"3Q  ��D    � (�8\�iEm`;Mxd��x��Q�8 l|BNLt@mLu �6@odtZ4 T0 k� ��O��O	E1 4#Q&�1D"3Q  ��D    � (�8\�iEm\<Mxd��x��Q�8 l|BNLt@mHu �6@ohtZ4 T0 k� ��O��O	E1 4#Q&�1D"3Q  ��D    � (�8\�iEm\=Mxd��x��R�8 l|BNPt@mHu �6@ohtZ4 T0 k� ��P��P	E1 4#Q&�1D"3Q  ��D    � (�8\�hEmX?Mxd}�x��R�8 l|BNPt@mHu �6@ohtZ4 T0 k� ��P��P	E1 4#Q&�1D"3Q  ��D    � (�8\�hD=X@Mtd~ x��R�8 l|BNTt@mHv �6@ohtZ4 T0 k� ��P��P	E1 4#Q&�1D"3Q  ��D    � (�8\�hD=TBMtd~ x��S�8 l|BNTs@mHv �6@oltZ4 T0 k� ��Q��Q	E1 4#Q&�1D"3Q  ��D    � (�8\�hD=TCMtd~x��S�8 l|BNXs@mHv �6@oltZ4 T0 k� ��Q��Q	E1 4#Q&�1D"3Q  ��D    � (�8\�hD=PEMtd~x��S�8 l|BNXs@mDv �6@oltZ4 T0 k� ��Q��Q	E1 4#Q&�1D"3Q  ��D    � (�8\�hD=PFMpd~x��T�8 l|BN\s@mDw �6@oltZ4 T0 k� ��R��R	E1 4#Q&�1D"3Q  ��D    � (�8\�gEmLHMpd~x��T�8 l|BN\s@mDw �6@oltZ4 T0 k� ��R��R	E1 4#Q&�1D"3Q  ��D    � (�8\�gEmHJMpd~x��T�8 l�BN\s@mDw �6@optZ4 T0 k� ��R��R	E1 4#Q&�1D"3Q  ��D    � (�8\�gEmHKMpd~x��U�8 l�BN`r@mDw �6@optZ4 T0 k� ��S��S	E1 4#Q&�1D"3Q  ��D    � (�8\�gEmDMMpd~x��U�8 l�BN`r@mDw �6@optZ4 T0 k� ��S��S	E1 4#Q&�1D"3Q  ��D    � (�8l�gEm@OMld~w��U�8 l�BN`r@m@x �6@opsZ4 T0 k� ��S��S	E1 4#Q&�1D"3Q  ��D    � (�8l�gEm<PMldnw��V�8 l�BNdr@m@x �6@opsZ4 T0 k� ��T��T	E1 4#Q&�1D"3Q  ��D    � (�8l�gEm8RMldnw��V�8 l�BNdr@m@x �7@otsZ4 T0 k� ��T��T	E1 4#Q&�1D"3Q  ��D    � (�8l�fEm8SMldnv��V�8 l�BNhr@m@x �7@otsZ4 T0 k� ��T��T	E1 4#Q&�1D"3Q  ��D    � (�8l�fEm4UMldnv��W�8 l�BNhr@m@x �7@otsZ4 T0 k� ��T��T	E1 4#Q&�1D"3Q  ��D    � (�8l�fEm0VMhdnv��W�8 l�BNhq@m@x �7@otsZ4 T0 k� ��U��U	E1 4#Q&�1D"3Q  ��D    � (�8l�fEm0XMhdnu��W�8 l�BNlq@m@y  7@otsZ4 T0 k� ��U��U	E1 4#Q&�1D"3Q  ��D    � (�8l�fEm,YMhdnu��W�8 l�BNlq@m@y  7@otsZ4 T0 k� ��U��U	E1 4#Q&�1D"3Q  ��D    � (�8l�fEm,ZMhdnt��X�8 l�BNlq@m<y  7@oxsZ4 T0 k� ��V��V	E1 4#Q&�1D"3Q  ��D    � (�8l�fEm([Mhd^t��X�8 l�BNpq@m<y  7@oxsZ4 T0 k� ��V��V	E1 4#Q&�1D"3Q  ��D    � (�8l�fEm(\Mhd^s��X�8 l�BNpq@m<y  7@oxsZ4 T0 k� ��V��V	E1 4#Q&�1D"3Q  ��D    � (�8l�eE}(]Mdd^s��X�8 l�BNpq@m<y  7@oxsZ4 T0 k� ��V��V	E1 4#Q&�1D"3Q  ��D    � (�8l�eE}$^Mdd^r��Y�8 l�BNtp@m<z  7@oxsZ4 T0 k� ��W��W	E1 4#Q&�1D"3Q  ��D    � (�8l�eE}$_Mdd^r��Y�8 l�BNtp@m<z  7@oxsZ4 T0 k� ��W��W	E1 4#Q&�1D"3Q  ��D    � (�8l�eE}$`Mdd^q��Y�8 l�BNtp@m<z  7@o|sZ4 T0 k� ��W��W	E1 4#Q&�1D"3Q  ��D    � (�8l�eE} `Mdd^q��Y�8 l�BNxp@m<z  7@o|sZ4 T0 k� ��W��W	E1 4#Q&�1D"3Q  ��D    � (�8l�eE} a=`d�p��Z�8 l�BNxp@m8z  7@o|sZ4 T0 k� ��X��X	E1 4#Q&�1D"3Q  ��D    � (�8l�eE}b=`d�p��Z�8 l�BNxp@m8{  7@o|rZ4 T0 k� ��X��X	E1 4#Q&�1D"3Q  ��D    � (�8l�eE�b=`d�o��Z�8 l�BN|p@m8{  7@o|rZ4 T0 k� ��X��X	E1 4#Q&�1D"3Q  ��D    � (�8l�dE�c=`d�o��[�8 l�BN|p@m8{  7@o�rZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8l�dE�c=`d� n��[�8 l�BN|o@m8{  7@o�rZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8l�dE�c`d� n��[�8 l�BN�o@m8{  7@o�rZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8l�dE�c`e��n��[�8 l�BN�o@m8{  7@o�rZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8l�dKmc`e��m��[�8 l�BN�o@m8{ 7@o�rZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8l�dKmc\e��m��\�8 l�BN�o@m8| 7@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D    � (�8l�dKmc\e��m��\�8 l�BN�o@m8| 7@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D    � (�8l�dKmc=\e��l��\�8 l�BN�o@m4| 7@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D    � (�8l�dKmc=\e��l��\�8 l�BN�o@m4| 8@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D    � (�8l�dKmc=\e�l��\�8 l�BN�o@m4| 8@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D    � (�8l�cKmc=\e�l��\�8 l�BN�n@m4| 8@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D   � (�8l�cKmc=\e�l��\�8 l�BN�n@m4| 8@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D   � (�8l�cKmcm\e�l��\�8 l�BN�n@m4| 8@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D    � (�8l�cKmcm\e�l��\�8 l�BN�n@m4} 8@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D    � (�8l�cKmcm\e�l��\�8 l�BN�n@m4} 8@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D    � (�8l�cK}cm\e�l��\�8 l�BN�n@m4} 8@o�rZ4 T0 k� ��Z��Z	E1 4#Q&�1D"3Q  ��D    � (�8l�cK}cmXe�l �\�8 l�BN�n@m4} 8@o�rZ4 T0 k� ��Y� Y	E1 4#Q&�1D"3Q  ��D    � (�8l�cK}c
Xe�l �\�8 l�BN�n@m4} 8@o�rZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8l�cK}c
Xe�l �\�8 l�BN�n@m4} 8@o�rZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8l�cK}c
Xe�l �\�8 l�BN�n@m0} 8@o�rZ4 T0 k� � X�$X	E1 4#Q&�1D"3Q  ��D    � (�8l�cKmc
Te�l �\�8 l�BN�n@m0} 8@o�rZ4 T0 k� �$X�(X	E1 4#Q&�1D"3Q  ��D    � (�8\�cKmc
Te�l �\�8 l�BN�n@m0} 8@o�rZ4 T0 k� �(X�,X	E1 4#Q&�1D"3Q  ��D    � (�8\�bKmc
Te�l �\�8 l�BN�m@m0~ 8@o�rZ4 T0 k� �,X�0X	E1 4#Q&�1D"3Q  ��D    � (�8\�bKmc
Pe-�l �\�8 l�BN�m@m0~ 8@o�qZ4 T0 k� �0X�4X	E1 4#Q&�1D"3Q  ��D    � (�8\�bKmc
Le-�l �\�8 l�BN�m@m0~ 8@o�qZ4 T0 k� �0X�4X	E1 4#Q&�1D"3Q  ��D    � (�8\�bJc
Le-�l��\�8 l�BN�m@m0~ 8@o�qZ4 T0 k� �Y� Y	E1 4#Q&�1D"3Q  ��D    � (�8\�bJc
He-�l��\�8 l�BN�m@m0~ 8@o�qZ4 T0 k� �Y�Y	E1 4#Q&�1D"3Q  ��D    � (�8��bJc
Df-�l��\�8 l�BN�m@m0~ 8@o�qZ4 T0 k� �Y�Y	E1 4#Q&�1D"3Q  ��D    � (�8��bJc
-Df-�l��\�8 l�BN�m@m0~ 8@o�qZ4 T0 k� � Y�Y	E1 4#Q&�1D"3Q  ��D    � (�8��bJc
-Df-�l��\"8 l�BN�m@m0~ 8@o�qZ4 T0 k� ��Y� Y	E1 4#Q&�1D"3Q  ��D    � (�8��aJ c
-Df-�l��\"8 l�BN�m@m0~ 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��aJ c
-@f-�l��\"8 l�BN�m@m0~ 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8�aJ c
-@f-�l��\"8 l�BN�m@m0 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8�`J�c<f-�l��\"8 l�BN�m@m0 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8�`J�c<f-�l��\"8 l�BN�m@m0 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8�_J�c<f-�l��\"8 l�BN�m@m, 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8�^J�c8f-�l��\"8 l�BN�m@m, 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��^J�c8f-�l��\"8 l�BN�l@m, 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��]J�c-8f-�l��\"8 l�BN�l@m, 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��]J�c-8f-�l��\"8 l�BN�l@m, 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D   � (�8��\J�c-4f-�l��\�8 l�BN�l@m, 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��\J�c-4f-�l��\�8 l�BN�l@m, 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��[J�c-4f-�l��\�8 l�BN�l@m, 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��[K��c
M0f-�l��\�8 l�BN�l@m, 8@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��ZK��c
M0f-�l��[�8 l�BN�l@m,� 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��ZK��c
M0f-�l��[�8 l�BN�l@m, 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��ZK��c
M0f-�l��[�8 l�BN�l@m, 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��YK��c
M0f-�l��[�8 l�BN�l@m, 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��YK��c
M,f-�l��[�8 l�BN�l@m, 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��YK��c
M,f-�l��[�8 l�BN�l@m,~ 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��XK��c
M,f-�l��[�8 l�BN�l@m,~ 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��XK��c
M,f-�l��[!�8 l�BN�l@m,~ 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��XK��c
M,f-�l��[!�8 l�BN�l@m,~ 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��XK��c
M,f-�l��[!�8 l�BN�l@m,} 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��XK��c
],f-�l��[!�8 l�BN�l@m,} 9@o�qZ4 T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��D    � (�8��XK��c
],f-�l��[!�8 l�BN�l@m,} 9@o�qZ4 T0 k� ��Y� Y	E1 4#Q&�1D"3Q  ��D    � (�8��XK��c
],f-�l��[!�8 l�BN�l@m,} 9@o�qZ4 T0 k� ��Y� Y	E1 4#Q&�1D"3Q  ��D    � (�8��XK��d
],f-�l��[!�8 l�BN�l@m(} 9@o�qZ4 T0 k� ��Y� Y	E1 4#Q&�1D"3Q  ��D    � (�8��XK��d
],e-�l��[!�8 l�BN�k@m(| 9@o�qZ4 T0 k� ��Y� Y	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
M(e-�k��[!�8 l�BN�k@m(| 9@o�qZ4 T0 k� ��X� X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
M(e-�k��[!�8 l�BN�k@m(| 9@o�qZ4 T0 k� ��X� X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
M(e-�k��[!�8 l�BN�k@m(| 9@o�qZ4 T0 k� ��X� X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
M(e-�k��[�8 l�BN�k@m(| 9@o�qZ4 T0 k� ��X� X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
M(e-�k��[�8 l�BN�k@m({ 9@o�qZ4 T0 k� ��X� X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
M(e�k��[�8 l�BN�k@m({ 9@o�qZ4 T0 k� ��X� X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
M(e�k��[�8 l�BN�k@m({ 9@o�qZ4 T0 k� ��X� X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
M(d�k��[�8 l�BN�k@m({ 9@o�qZ4 T0 k� ��X� X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
M(d�k� [�8 l�BN�k@m({ 9@o�qZ4 T0 k� ��X� X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
](c�k� [�8 l�BN�k@m(z 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
](c|k� [�8 l�BN�k@m(z 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��d
](c|k� [�8 l�BN�k@m(z 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��e
]$b|k� [�8 l�BN�k@m(z 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��e
]$b|l� [�8 l�BN�k@m(z 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��e
]$bxl� [�8 l�BN�k@m(z 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��e
]$bxl� [�8 l�BN�k@m(y 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��e
]$b}xl� [�8 l�BN�k@m(y 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��e
]$b}tl� [�8 l�BN�k@m(y 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��e
]$b}tm� [�8 l�BN�k@m(y 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��e
]$b}tm� [�8 l�BN�k@m(y 9@o�qZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��e
M$b}pn� [�8 l�BN�k@m(y 9@o�pZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��f
M$b�pn� [�8 l�BN�k@m(y 9@o�pZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D   � (�8 �XK��f
M$b�pn� [�8 l�BN�k@m(x 9@o�pZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��f
M$b�lo�[�8 l�BN�k@m(x 9@o�pZ4 T0 k� � X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��f
M$b�lo�[�8 l�BN�k@m(x 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��f
$b�hp�[�8 l�BN�k@m(x 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��f
 bhp�[�8 l�BN�k@m(x 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��f
 bdq [�8 l�BN�k@m(x 9@o�pZ4 T0 k� �W�W	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��f
 bdq [�8 l�BN�k@m$x 9@o�pZ4 T0 k� �$W�(W	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��f
bdr [�8 l�BN�k@m$x 9@o�pZ4 T0 k� �0W�4W	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��f
bdr [�8 l�BN�k@m x 9@o�pZ4 T0 k� �8W�<W	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��g
b-`r [�8 l�BN�k@m x 9@o�pZ4 T0 k� �<W�@W	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��g
b-`r [�8 l�BN�j@m x 9@o�pZ4 T0 k� �@W�DW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��g
b-\r [�8 l�BN�j@mx 9@o�pZ4 T0 k� �DW�HW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��g
-b-\r [�8 l�BN�j@mx 9@o�pZ4 T0 k� �HW�LW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��g
-b-Xr [�8 l�BN�j@mx 9@o�pZ4 T0 k� �HW�LW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��g
-b
MXr [�8 l�BN�j@mx 9@o�pZ4 T0 k� �HW�LW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��g
-b
MTr [�8 l�BN�j@mx 9@o�pZ4 T0 k� �HW�LW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��g
-b
MTr [�8 l�BN�j@mx 9@o�pZ4 T0 k� �HW�LW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��h
-b
MTr [�8 l�BN�j@mx 9@o�pZ4 T0 k� �HW�LW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��h
-b
MTr [�8 l�BN�j@my 9@o�pZ4 T0 k� �HW�LW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��h
-b�Pr [�8 l�BN�j@my 9@o�pZ4 T0 k� �HW�LW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��h
-b�Pr [�8 l�BN�j@my 9@o�pZ4 T0 k� �HW�LW	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��h
-b�Lr�[�8 l�BN�j@my 9@o�pZ4 T0 k� �8X�<X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��h
b�Lr�[�8 l�BN�j@my 9@o�pZ4 T0 k� �,X�0X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��h
b�Lr�[�8 l�BN�j@my 9@o�pZ4 T0 k� � X�$X	E1 4#Q&�1D"3Q  ��D    � (�8 �XK��h
b�Hr�[�8 l�BN�j@my 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XJ�h
b�Hr�[�8 l�BN�j@my 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XJ�h
b�Dr�[�8 l�BN�j@my 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XJ�h
b�Dr�[�8 l�BN�j@my 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XJ�h
b�Dq�[�8 l�BN�j@my 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XJ�i�b�@q�[�8 l�BN�j@my 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XB��i�b�@q�[�8 l�BN�j@my 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XB��h�b�@q�[�8 l�BN�j@m y 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XB��h�b�<q�[�8 l�BN�j@m y 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XB��h�b�<q�[�8 l�BN�j@m z 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XB��h�b�<q�[�8 l�BN�j@l�z 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XB��h�b�8q�[�8 l�BN�j@l�z 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �XB��h�b�8q�[�8 l�BN�j@l�z 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �WB��h�b�8q�[�8 l�BN�j@l�z 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �WB��h�b�4q�[�8 l�BN�j@l�z 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8 �WB��h�b�4q�[�8 l�BN�j@l�z 9@o�pZ4 T0 k� �X�X	E1 4#Q&�1D"3Q  ��D    � (�8�1DA'��*_S����|0��E���D@{�'�EB�Z3�T0 k� ��	��		E1 4#Q&�1D"3Q  ��9 	   � ���2DA#��*OK���|0��E�{�D@w��EB�Z3�T0 k� ��	��		E1 4#Q&�1D"3Q  ��9 	   � ����2DA��*OC���|0��E�s�D@s��EB�Z3�T0 k� ��
��
	E1 4#Q&�1D"3Q  ��9 	   � ����3Ea��*O;��߳|0���E�o�D@k��EB�Z3�T0 k� ��
��
	E1 4#Q&�1D"3Q  ��9 	   � ����4Ea��*O3��׳|0��D�g�D@g��EB�Z3�T0 k� ��
��
	E1 4#Q&�1D"3Q  ��9 	   � ����5Ea���+O+��ϴ|0�D�_�DP_���EB�Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��9 	   � ����5E`����+O#��ô|0�D�[�DP[���EB�Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��9 	   � ����6E`���+O��|0ۯD�S�DPS���EB�Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��9 	   � ����7E`���+O��|0ǯD�G�DPG�/��EBtZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��9 	   � ��Ѽ8E`���+O���|0��D�C�DPC�/��EBpZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��9 	   � ��Ѵ9EP���+N����|0﷯D�;�DP;�/��EBlZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��9 	   � ��Ѭ9EP���+N����|0ﯯD�7�DP3�/��EBdZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��9 	   � ��Ѥ:EP���+>����|0燐D�/�DP/�/��EB`Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��9 
   � ���:EP���+>���|0D�+�E�'�/� EB\Z3�T0 k� �x�|	E1 4#Q&�1D"3Q  ��9 
   � ���;EP���t+>��w�|0D�#�E��/�EBXZ3�T0 k� �p�t	E1 4#Q&�1D"3Q  ��9 
   � ���;EP���l,>��o�|0D��E��/�EBTZ3�T0 k� �h�l	E1 4#Q&�1D"3Q  ��9 
   � ���<EP���d,>��g�|0D��E��/�EBPZ3�T0 k� �`�d	E1 4#Q&�1D"3Q  ��9 
   � ���x<EP���\,>��_�|0�{�D��E��/�EBHZ3�T0 k� �X�\	E1 4#Q&�1D"3Q  ��9 
   � ���h=EP���L,>��O�|0�k�D��E���?|EB@Z3�T0 k� �H�L	E1 4#Q&�1D"3Q  ��9 
   � ���`=EP���D,N��C�|0?c�D��E���?tEB<Z3�T0 k� �@�D	E1 4#Q&�1D"3Q  ��9 
   � ��1X=E@���<,N��;�|0?[�D���E���?lEB8Z3�T0 k� �8�<	E1 4#Q&�1D"3Q  ��9 
   � ��1P>E@��0,N��3�|0?S�D���E���?dEB4Z3�T0 k� �0�4	E1 4#Q&�1D"3Q  ��9 
   � ��1D>E@w��(,N��+�|0?K�D��E���?\EB0Z3�T0 k� �(�,	E1 4#Q&�1D"3Q  ��9 
   � ��1<>E@o�� ,N��#�|0?C�D��D����TEB,Z3�T0 k� �$�(	E1 4#Q&�1D"3Q  ��9 
   � ��14>E@g��,N���|0	�;�D���D����LEB(Z3�T0 k� �� 	E1 4#Q&�1D"3Q  ��9    � ��Q,>E@_��-N���|0	�3�D���D����D	EB$Z3�T0 k� ��	E1 4#Q&�1D"3Q  ��9    � ��Q>E@O� -N���|0	�'�D���D����4
EBZ3�T0 k� ��	E1 4#Q&�1D"3Q  ��9    � ��Q>E@G��-N{���|0	��D���D����,EBZ3�T0 k� ��	E1 4#Q&�1D"3Q  ��9    � ��Q?C�?��-Ns��|0	��D���D����$EBZ3�T0 k� ��� 	E1 4#Q&�1D"3Q  ��9    � ��Q ?C�7��-No���|0	��D���D����EBZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �}P�?C�/��-^g��߹|0	��D���D���oEBZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �{P�?C�'��-^c��׹|0	��D���D���oEBZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �yP�?C���-^[��˹|0	��D���D���o EBZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �v��?C���-^W��ù|0���D���D���n�EBZ3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �s��?C���-^S�ỹ|0���D���D���n�EB Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �q��?C���- �K�᳹|0��D���D���N�EA�Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �o�?C����- �C�᣹|0��D���D���N�EA�Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �m�@C����. �;�᛺|0�ߨD���D���N�EA�Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �k�@C����. �7�ᏺ|0�ۨD���D���N�EA�Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �i�@C����. �3�ᇺ|0�ӧD���D��N�EA�Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��9    � �f��@C���|. �/���|0�ϧD���D���EA�Z3�T0 k� �� �� 	E1 4#Q&�1D"3Q  ��9    � �d��@C���t. �'��w�|0�ǧD���D�|�EA�b��T0 k� ��"��"	E1 4#Q&�1D"3Q  ��9    � �b��@C���l. �#��o�|0�æD���D�x�EA�b��T0 k� �t"�x"	E1 4#Q&�1D"3Q  ��9    � �`��@C���d. ���g�|0���D��D�t
�E��b��T0 k� �h#�l#	E1 4#Q&�1D"3Q  ��9    � �^�x@C���\. ���_�|0���D�{�D�p�E��b��T0 k� �`$�d$	E1 4#Q&�1D"3Q  ��9    � �\�p@C���T. ���S�|0���D�s�D�l�E��b��T0 k� �X%�\%	E1 4#Q&�1D"3Q  ��9    � �Z�h@C����H. ���K�|0���D�o�D�h�E��
b��T0 k� �P%�T%	E1 4#Q&�1D"3Q  ��9    � �X�`@C����@. ���C�|0���D�g�D�d�E��
b��T0 k� �H&�L&	E1 4#Q&�1D"3Q  ��9    � �V�T@C����8. ���;�|0���D�c�Eo`xE��	b��T0 k� �<'�@'	E1 4#Q&�1D"3Q  ��9    � �T�LAC����0. ���3�|0���D�[�Eo\pE��	b��T0 k� �4(�8(	E1 4#Q&�1D"3Q  ��9    � �R�<AC���� .����#�|0���D�O�EoT`E��b��T0 k� �$)�()	E1 4#Q&�1D"3Q  ��9    � �P�4AC����.����|0���EoK�EoP.XE��Z3�T0 k� � *�$*	E1 4#Q&�1D"3Q  ��9    � �N�,AC����/����|0��EoC�EoL .PEѸZ3�T0 k� �+� +	E1 4#Q&�1D"3Q  ��9    � �L�$AC����/����|0�Eo?�EoH#.HC�Z3�T0 k� �,�,	E1 4#Q&�1D"3Q  ��9    � �J AC����/��� ��|0{�Eo7�EoD%.@C�Z3�T0 k� �-�-	E1 4#Q&�1D"3Q  ��9    � �H AC�w���/��� ��|0w�Eo3�Eo@'.8C�Z3�T0 k� �.�.	E1 4#Q&�1D"3Q  ��9    � �G AC�o���/��� �|0s�Eo+�Eo<).0 C�Z3�T0 k� ��/� /	E1 4#Q&�1D"3Q  ��9    � �F  AC�k���/��� �|0	�o�Eo'�E_4+.(!C�Z3�T0 k� ��/��/	E1 4#Q&�1D"3Q  ��9    � �E�AC�c���/��� ۼ|0	�k�Eo�E_0-. "C�Z3�T0 k� ��0��0	E1 4#Q&�1D"3Q  ��9    � �D�AC�S���/��� ˼|0	�c�Eo�E_(1.$C�Z3�T0 k� ��2��2	E1 4#Q&�1D"3Q  ��9    � �C�AC�K���/�� ü|0	�_�EoE_ 3.%C�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    � �B�BC�C��/����|0
[�EoE_5> &C�bs�T0 k� ��5��5	E1 4#Q&�1D"3Q  ��9    � �A�BC�;��/����|0
[�E_ E_7=�'C�|bs�T0 k� ��7��7	E1 4#Q&�1D"3Q  ��9    � �@�BC�3��/����|0
W�E^�E_9=�(C�tbs�T0 k� ��8��8	E1 4#Q&�1D"3Q  ��9    � �?�BC�+��/����|0
S�E^�E_;=�)C�pbs�T0 k� ��9��9	E1 4#Q&�1D"3Q  ��9    � �>�BC�#��/����|0	
S�E^�E_==�*C�hbs�T0 k� ��:��:	E1 4#Q&�1D"3Q  ��9    � �=�BC����/����|0		�O�E^�
E^�?=�+C�`bs�T0 k� ��;��;	E1 4#Q&�1D"3Q  ��9    � �<�BC�� |/���|0
	�K�E^�EN�C=�-C�Tbs�T0 k� ��=��=	E1 4#Q&�1D"3Q  ��9    � �;�BC�� t/��w�|0
	�K�E^�EN�D=�.C�Lbs�T0 k� ��>��>	E1 4#Q&�1D"3Q  ��9    � �:�BC��� l/��o�|0
	�G�C��EN�F=�/C�Dbs�T0 k� ��?��?	E1 4#Q&�1D"3Q  ��9    � �9�BC��� d/��g�|0

G�C��EN�G=�0C�< bs�T0 k� ��@��@	E1 4#Q&�1D"3Q  ��9    � �8xBC��� \0���[��0
G�C��EN�IM�1C�4 Z3�T0 k� �xA�|A	E1 4#Q&�1D"3Q  ��9    � �8pBC��� P0� �S��,
G�C�EN�JM�2C�, Z3�T0 k� �pB�tB	E1 4#Q&�1D"3Q  ��9    � �8hBC��� H0��K��,
C�C�C��KM�3D'�Z3�T0 k� �hC�lC	E1 4#Q&�1D"3Q  ��9    � �8�TBC��� 80x�;��, C�C�C��NM�5D�Z3�T0 k� �\E�`E	E1 4#Q&�1D"3Q  ��9    � �8�LBC��� 00t�3��, C�C�C��O݈6D�Z3�T0 k� �XA�\A	E1 4#Q&�1D"3Q  ��9    � �8�DCC���(0p�'��, ?�C�C��P݀7D�Z3�T0 k� �T>�X>	E1 4#Q&�1D"3Q  ��9    � �8�<CC��� 0l���, ?�C�C��Q�x8E��Z3�T0 k� �P<�T<	E1 4#Q&�1D"3Q  ��9    � �8�4CC���0h���, ?�C�C��R�p9E���Z3�T0 k� �H;�L;	E1 4#Q&�1D"3Q  ��9    � �8�,CC���0d���, n?�C�C��S�h:E���Z3�T0 k� �@;�D;	E1 4#Q&�1D"3Q  ��9    � �8� CC���0`���( n?�C�xC��T�`;E���Z3�T0 k� �8;�<;	E1 4#Q&�1D"3Q  ��9    � �8�CC����0\����( n?�C�pC��U�X<E���Z3�T0 k� �0;�4;	E1 4#Q&�1D"3Q  ��9    � �8�CC�{��0T	���( n?�C�d!C�tV�H>E���Z3�T0 k� � <�$<	E1 4#Q&�1D"3Q  ��9    � �8� CC�s��0T
���( �?�C�\"C�lW�D?E���Z3�T0 k� �=� =	E1 4#Q&�1D"3Q  ��9    � �8��CC�k��0P�ۿ�( �?�C�T#C�dW�<?E���Z3�T0 k� �=�=	E1 4#Q&�1D"3Q  ��9    � �8��CC�c��0�L�ӿ�( �?�C�L$C�\X�4@E��Z3�T0 k� �>�>	E1 4#Q&�1D"3Q  ��9    � �8��CC�[���0�H�˿�( �?�C�D%C�TX�,AE��Z3�T0 k� �?�?	E1 4#Q&�1D"3Q  ��9    � �8��CC�S���0�D�ÿ�$ �?�C�<&C�LY�$BE��Z3�T0 k� ��@� @	E1 4#Q&�1D"3Q  ��9    � �8��CC�C��0�<����$;�C�0(C�<Z�DE���Z3�T0 k� ��<��<	E1 4#Q&�1D"3Q  ��9    � �8��CC�;��0�8O���$;�D()C�4Z�DE���Z3�T0 k� ��9��9	E1 4#Q&�1D"3Q  ��9    � �8��CC�3��0�4O���$;�D *C�,Z�EE���Z3�T0 k� ��7��7	E1 4#Q&�1D"3Q  ��9    � �8��CC�+��0�,O���$;�D+C� Z��FE���Z3�T0 k� ��5��5	E1 4#Q&�1D"3Q  ��9    � �8��CC�#��0�(O���$;�D,C�[��FE�{�Z3�T0 k� ��4��4	E1 4#Q&�1D"3Q  ��9    � �8��CC���0�$O���$�;�D-C�[��GD0s�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    � �8��DC���t1�Ow�� �7�D�/C� [��HD0c�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    �  �8�DC���h1�Oo�� �7�D�0C��[��HD0[�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    �  �8�DC����`1�Oc�� �7�D�1C��[��HD0W�Z3�T0 k� ��2��2	E1 4#Q&�1D"3Q  ��9    �  �8xDEM��X1�O[�� �3�D�2C��Z��ID0O�Z3�T0 k� ��2��2	E1 4#Q&�1D"3Q  ��9    � !�8lDEM��P1��S���3�D�3C��Z�ID0G�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    � !�8dDEM��H1���K���/�D�3EM�Z��ID0?�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    � !�8�TDEMӺ�81���;���+�D�5EM�Z��ID0/�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    � !�8�LDEM˹�,1���3���'�D�6EM�Y��ID0'�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    � !�8�DCEMø�$1���+���'�D�7EM�Y��ID0�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    � !�8�<CEM���1���#���#�D�8EM�X��ID@�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    � !�8�4CEM���1�������D�8EM�X��ID@�Z3�T0 k� ��3��3	E1 4#Q&�1D"3Q  ��9    � !�8� CEM���1�������D�:EM�W�pIDO��Z3�T0 k� �|3��3	E1 4#Q&�1D"3Q  ��9    � !�8�BEM����1������N�D�;EM�W�lIDO��Z3�T0 k� �x2�|2	E1 4#Q&�1D"3Q  ��9    � !�8>BE=����1�����N�D�;EMtV�dHDO��Z3�T0 k� �p2�t2	E1 4#Q&�1D"3Q  ��9    � !�8>BE=����0������N�C�|<EMlV�\HDO� Z3�T0 k� �h2�l2	E1 4#Q&�1D"3Q  ��9    � !�8> BE=����0������N�C�t=E=dUTGDO� Z3�T0 k� �h3�l3	E1 4#Q&�1D"3Q  ��9    � !�8=�AE=w���0������M��C�d>E=PTHGDO�Z3�T0 k� �d3�h3	E1 4#Q&�1D"3Q  ��9    � !�8	��AE=s���0������M��C�\?E=HS@FDO�Z3�T0 k� �`4�d4	E1 4#Q&�1D"3Q  ��9    � !�8                                                                                                                                                                            � � �  �  �  d A�  �K����   �      6 \��� ]�$�$� �  �� W�          ��.��     W��.��                     	 Z�8           @     ���   (
	           h�  / /      ��4&�     h�b�4p    ��p          P	 Z�8         ��     ���   
	           b�   � �
      �D��     b��D��                   W	 Z�8�          ���     ���   8	 

          q�N   � �
	   �Mp�     q��M��    �|�B            V	 Z�8          ��    ���   0
3
          [�`   � �
     /���r     [�`���Y       �              Z�8           0�  #  ���   H


          ��  ��     C��/     ���/                           ���S              y  ���    		 5 	            �4          W�%c�     �m�%`(     W 4                 �         ]�     ��B   0
&


          j� $ $      k��b�     j����U�    �� �               6 �              ��@   (
 
           zg�         �>�     zY]�>�}     ���                   �         :@     ��H   0	
           9�           ��<�     9�N�9�      ,                     �         	  �     ��@   H	$
          p��      ���z�     p����s       s                 
   �         
 �     ��@   03 
           ؠ��     � ��     � ��     S                         ����               ��@   P		 5                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          X�w  ��        �����     X�w����       � "                 x                j  �       �                          X    ��       ���       X  ��           "                                                 �                         �.�4�D�M����%���>��� ������     	           
 
   �   �:� '��E       �� `e� �d @f� �� 0g  �� �c` �� d` � d� �$  d� �d d� �� e  �� @f� �d  g  
�� W� 
� X  <� f� <� f� <�  f� <�  _` >  n` ;� s` ;� s� 
� W  
�\ W  
�< W� 
�| W� 
�\ X  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �d �Q� � }����� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����8�� (�� �  ������  
�fD
��L���"����D"� �  " `   J jF��     �j   
��
��
���    "�j��" " �
� �  �  
�  [��  ��     ���       [��  ��     ���       z    ��     ��>          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �D      �� �  ���        � � �  ���        �        ��        �        ��        �    ��     X-7����        ��                         襩 4  ���                                      �                ����             [�����&��   (�8��               13 Teemu Selanne       3:29                                                                        3  3     �� �� �c�
 � CC �CD � CJ �CK  �cW � �	c_ � �
B�( �J�4 � J�4 �kI �k�9 �	C/ �C1 �C1 �C? � C#? � C$O �C%O � C'G � C(D �C/* �C5" qC9: � �- � �, _kk; o ksK �"�# �  "�5 �!�# �"
�2 �#"�# � $"�5 �%"�# �&*�2 �'"�F � ("�X �)�B �*
�Q � +*�  ,*Mx -*Sx  .*�@  *LX � 0*Bx � 1*Qx2*=x8 3*E`P 4*ShX 5*LpX  *LPP 7*DhX 8*HpX  *LPX :*HpX  *LPX  *LPX  *LPX >*HpX  *LP                                                                                                                                                                                                                         �� R         �    @ 
        �     ` P E d  ��                    ������������������������������������� ���������	�
���������                                                                                          ��    �HB�� ��������������������������������������������������������   �4, :   6 �� = � m�� ���@���@����z�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             N    .    �� 
İJ      �                             ������������������������������������������������������                                                                                                                                       ����  �  �                                           ���� ��������� � ������������������������� �������� ������ ��������������������������������  ��� ���� ��������������������� � ������������������ ���� ������������ � ������� ���������� ����������������������������� �����������������  �� ������                                   !    *    �� ��J      )  	                           ������������������������������������������������������                                                                                                                                             ����  ��                                             �  ������ ������� �����������  ���������  ����������� ������� �� ������������������ �������� � ����� � � �� � �������������� �������������������������� ����������������� ��������  ����� ������ ����������� ������ �������������������                                                                                                                                                                                                                                                                           	                                                 �              


             �   }�           8�  0�             O     [                                                      ���      �  �����  8���������������������������������������������������������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � �~� �\                                                                                                                                                                                                                                                                                      )n)n
  
F                        m      a                  m      f                                                                                                                                                                                                                                                                                                                                                                                                                       > �  
>�  P�  @�  $#�  EZm} �ɬ�D�̎����� `�f��&�˖� �N 7����y�����y�                       � {        $   �   & QW  �  �                  �                                                                                                                                                                                                                                                                                                                                    0 U K          
              !��                                                                                                                                                                                                                            Z   �� �� ����      �� M      ���� ��������� � ������������������������� �������� ������ ��������������������������������  ��� ���� ��������������������� � ������������������ ���� ������������ � ������� ���������� ����������������������������� �����������������  �� �������  ������ ������� �����������  ���������  ����������� ������� �� ������������������ �������� � ����� � � �� � �������������� �������������������������� ����������������� ��������  ����� ������ ����������� ������ �������������������             $����������������UUUU�����UUU�U{�����������������UUUW����x�����w�����������������UUuU������wxwwww����������������WwwU�������wwwwx����������������UUUU����w�xw�w������������������Uuww���uUw��uU���Uz��uz��Wz��wzu�wYW�wxw�uxwwuW���������wx��UUwwX�xuy����u������wwww�wwwwwwwwwwwUUwWuUuu�UWW�wwwwy��x���x���ww�uwuuwwx��x�����Y����������w��www�wwwy��wyx�wyx��x�U���U���U���uy��u���u��uu��uU���wx��wxxwuW�WuuxU�uWW�UUU�uWu��W�y���wx�ww��wxx����wwwwwWwwwwwuW��ww��wx��w��xww��WwxUW�wWW�wy����w����������x�www��xwx�w��w�Ww����w��xwx�xwwwx�xwww��ww�wwwwwww�Wy�x�xuw��UwuwWwuwWwxwX�xwW�wuW�z�u�Y�u�X�u�U��yUU�Uuw�yUX��UX�uWwuWuwWwUwwUUUwUUWUUUUuUUWWUUWwwuW�WUW�XUuwx�UXx�Uxwwwxww�xww����ww��UwuwwW��ww��ww��ww��xw��xwwwwwwwwwwwwxwwwxuwwxwwwwUwwwWwwwwywX��yWx�Xxy�W��uXYwWuZ��u��w���ux���w���U���U���U���u���UZ��UWUUwWuUUU�Uu��Uw��UWx�UUW��UU��UUwwwxUwww��wx��������x���w���Ux�wx�wwwwww���w���U��ww��ww�wwwuwwwWwwxWwwywww�wwx�ww��xx��wx��w����WU��WY��uY��Wx��Wy�Uxz�Xw��Xw�W���W���U��������������������������UUW�uUUX�U�U�W�uWW��WU���u���WUUUWUUwuuwwwwx��wwx�wwwwwwwwuwwwWuwwWwwwuwwx�ww�wwwx�w�xxw��wx��xw�Uw��W���Xx�U��uW��UxwUWwwUwww�w�W�x�W�y�wx��wx�Wwx�Wyz�wz��x�q��    >      9      X                       M     �  �����J����'    ��     ~�      �      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ��  � ��     � ��   	 ��  p � ��  � �� 5� �� �� �z 5� �p �$ ^$ �u� 5�  �       �� � ��   ��     ��   � �� �� �z   ���� �$ ��  � �� h �� �� �� ��  �� �� �  �� �� �z � ��� �$ R �  ��R  �      �  ��   5�������2���� g��� 	       f ^�         ��  (      5      ���t���2�������J������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                         E  �\       U TUTQ�T\�jA���̪������ UTDDEUU�����j������������������DUP UUTD�����v����������������    U�UPUDDE��\����������������        U   TE ��@ x�@ �lE �|U  E� \� �Q� _ǪE�L��\��\�������������������E�lTP��E ��P �����������UDL�_UL�_L�UL�L�̪�������U������D���EU��E��E���E���������z��Q�j�T_�z �_�  T\  E��U ��T ����|��E |P �E  @  \��\��\��Ez� Oʪ UǪ \� Eʪ�P ��E �|�P���D��lϪ�����������L��L��L�UUL�QDL�_���Ua��̪��w���E��EU��E���E��DU�����wz��   �  �E �ETOQ���j����������UO  �T  ��P ��O ��� �����O���E  T\  E   T                   ����Ǫ��\ʪ�E\ʪUE\� UDU  UT    ����������������z������DUUUUTD�������������������|���UUTDDUU�����������̧|�T�TUUDP U       ��TQ�TE TE  E                   wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwtwwwCwwt1wwCwt1wC�t1��C1����������""""���������������!���""!����,���ww��7����������������wwwwwwwwwwwwwwwwwwww7wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwws��w1wt1�wC�t1��s��s��s������"$��Gw�!������������L���q��"r��������!�����!ww�r�w�ww!�wwrwwwwwwqwwwrwwww�7ww�ww�ww��7w��w���G��'!wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                               s   D   O   w   w   v   u   f   T   �   �              3@  DDp ��4 ��tp��wpO�tpdfwGfeTwfeWwfUFwdUFweTfp�DDp���p���@�w�p   C   D   O   D   w   u   U   U  F  d  f   f   D   �   �   �DD ���7���uP��e`O�V ffg ffG Ufw UU� FUN dFw ffp DDp ��p ��@ w�p  C4 4D@O�C���O�Dt�GVfeVfdFfdFfdUfffUfffwFff�DDD���� ���                    0   G   W   W   U   E   E   w   �   �   @    fg D� O�� �� w�}�w��}����������M���M���M��������y�                    �   �   �   �   �   �   �   �   ~   w       ���w���w���~���~�DMw�������������y�                        w���w}��wt��wt��w}M�����������   M   M   ~�  p�  p   p   p      �   �   �   �               vd  eVp ffpw�Op���w���G���M�}�                                     v   ub  ub  f   `   P               "  f  U` wfP        p   p   p   p   p   p   p   p                               C4 �y�                              f  vU`vf`D�O������p}�w�  ?�  ?�  ?�  33  3#                                      f  Ug                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 " ""   "" !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                                   " ""   "" !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  "!  " ! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �    �   �   "  "�  �                "   "   "�  �            "   "  !�    ��                ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                                                                                                                                                                            �   �  �  �  	�  �  EH  ET DU CE DD4 DD3 DC0 �3 ɰ �  ,�  +�  "/  ������ � ̹�p�˚��̹���ː�̼�̻���ۜ��۩�ݍ���=��J�ܰT�� EJ�0 EJ� I�  ��  �"  ""  "/  "�� ���                    ̰ ̻ ̻	���̚�w�ݸ�	��  ����̲����"/����  ��  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� �   �".  .                            �   �    �   �       �   �   �                .                        "  .���"    �     �                   ���������������������  ��  ��  ��  �   �    �          �         �                                                                                                                 "  "(��ȩ�ܚ��ۊ����� ��  �   �   �   �   �� ��� ̻� ˽� ��� �w� �������������������������� �̻ ���         �   �       �   �   "" �+� Ȼ� ɫ� ɨ� ��                �� �I��3 ��D 
UD 
UD TD  T�  ˸  ��  �� ̰ �+ ��"/ �"/  ����  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� �   �".  .                            �   �    �   �       �    �   �     �     �  �  "   "   "   "�  �                       "   "   "�  �                            �   ���                            �   "                                                                                                  "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             �"  �""� "�  ���� �                                                                                                                                                                                       ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   �"   ".   .                  �   �   �   �   �   �   �   �                .                      �"  �""� "�    �     �                                               ���                          ����                  �   �� �       �  �  "�  "   "                                                            �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �      ��    �                                                                                                                                                                                                                                                                                                             	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           "� /���  �       �   �   �                                                   ��                                              �".��".  ���    �                      �   �      ��   �  ��  �  �  �         � ".��".��/����  �                                                                                                                                             �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   �   " � ��      �    �                   Ͱ  ˻  ˻  ۻ  ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                            �".��".  ���    �                    ".  ".  ���                                                                                                                                                                                                                        	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           "� /���  �       �   �   �                                                   ��                     �   �                      �".��".  ���    �   .  .  "/ �� �   �                            � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                          �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �"  "�  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �                    ".  ".  ���  �   "  "  "   �                        �  � �                       � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                                               	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           "� /���  �       �   �   �                       ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �                    ".  ".  ���   ���� �                             � "�"  �    � � �                                                                                                                                                           �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ���������""��""��""�����        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                          2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ DD D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�GwDGwqwDDwtwwww3333DDDD �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�""""����������A��I��I = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=""""�����A�DA�I��I�    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"��������I���I���I���I��� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(XxMAMAMMMM�M�M����3333DDDD w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xwwD�����MD��M����3333DDDD  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���4���4���4���4���4���43334DDDD �  + � � � � � � � � � � ��	� � � ��� � � � � � � � � � � ��	� � � ��� �� ����(+((�""""wwwwqqqqwGwGGG ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""wwwwwwqqDAwG M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M������������������333DDD � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�M��M��D��M����������3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DD��D�M��D����3333DDDD 5 6  X � �F � � � � � ����� � ����������� � ����� � � � � ��	F ��(X((6(5""""������DH�H� x �  l � �G � � � � � � � � � � ������������� � � � � � � � � � ��	G ��l((�x""""�������H�H��D w w x y ������H���������������������������������H�����yxww""""��������H��H��H��H�  � + w�������I�J�K�L�M�N�O � � � � � � � � � � � � � � � � � � � ��O�N�M�L�K�J�I������w(+�(DD������L��DL����3333DDDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A e ��A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,L�A�AAD��DL�����3333DDDD +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�] � ځ]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+���4���4���4L��4L��4���43334DDDD 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U �h�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5""""���������M�MMM =  U ,     !d�P���e�f�g�!�!�!�k�!�!�!�l�!�!�!�!�k�!�!�!�l�!�!�!�g�f�e���P)d((( ((,(U((=""""�������A��AA     =  U , N ,�-�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�-(,(N(,(U((=((( ��������������333DDD � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � �I��I����������������3333DDDD � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � ���A���I��I���I�����3333DDDD m � �!�A�A� � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""������������������������  � �!�AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M""""������D�D��� 
 � �!�AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�""""������������������������ - � �!�!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�wqwwqwwwwwqwwwDwwww3333DDDD 69�:���  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5qqwwwDDwtGwwww3333DDDD x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xwww4www4www4www4www4www43334DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwqwwwqwqwq + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""wwwwwwwDwGwA � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(��A�L�L�L��L���333DDDLDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDD� �� �c�
 � CC �CD � CJ �CK  �cW � �	c_ � �
B�( �J�4 � J�4 �kI �k�9 �	C/ �C1 �C1 �C? � C#? � C$O �C%O � C'G � C(D �C/* �C5" qC9: � �- � �, _kk; o ksK �"�# �  "�5 �!�# �"
�2 �#"�# � $"�5 �%"�# �&*�2 �'"�F � ("�X �)�B �*
�Q � +*�  ,*Mx -*Sx  .*�@  *LX � 0*Bx � 1*Qx2*=x8 3*E`P 4*ShX 5*LpX  *LPP 7*DhX 8*HpX  *LPX :*HpX  *LPX  *LPX  *LPX >*HpX  *LP3333DDDDAqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD��������������������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ��������������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ��������������������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE��������������������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD��������������������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD��������������������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD��������������������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� ��%��:�L�S�S�L��0�R�S�\�U�K���������8�>�7���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� ����7�\�J��<�V�I�P�[�H�P�S�S�L�������8�>�7���""""������A�D��I��""""�������D����� ����>�L�L�T�\��=�L�S�H�U�U�L��������>��<���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �>��<������A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �8�>�7���"��""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,�����������DDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �����<�L�Z�\�T�L��2�H�T�L����������������� ����4�U�Z�[�H�U�[��<�L�W�S�H�`��������������� ����.�O�H�U�N�L��2�V�H�S�P�L���������������� ������0�K�P�[��7�P�U�L�Z���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            