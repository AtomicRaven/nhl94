GST@�                                                            \     �                                                       ��  p�            � ���*�
 J��������������t���        �g      #    t���                                d8<n    �  ?    L�����  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"    
 �j,� B ��
                                                                                  ����������������������������������      ��      UUU 111 ...  &&&  ���  ��� ���         444 444 444 444                 �E� !"!         :::�����������������������������������������������������������������������������������������������������������������������������=3  03  11  03  *          �  �  �  �    	    	              ��  ��  ��  ��                  $  
          ;5 �����������������������������������������������������������������������������                                ((  H�    ��   @  #   �   �                                                                                '  !�"E!�  
$    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�fO  �Z�� |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E E ܮ                                                                                                            ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ܀~E�ӹ^��L�|�5Y��3��B���  R��'���D`T0 k� ������e1�t B50A%1r  ��   ����8܈~E�׷^��L�|�5Y��3��B���  R��&���D\T0 k� ������e1�t B50A%1r  ��   ����8�}E�۴^��L�|�4Y��3��B��  R��%���D\T0 k� ������e1�t B50A%1r  ��   ����8�}E;߳^��L�|�3Y��3��B��  R��%���DXT0 k� ������e1�t B50A%1r  ��   ����8�}E;�^��L�|�3Y��3��B��  R��$���DXT0 k� ������e1�t B50A%1r  ��   ����8�}E;�N�L�|�2Y��3��B��  R��$��DXT0 k� ������e1�t B50A%1r  ��   ����8�}E;�Nw���|�2Y��3��B�#�  R��#��DTT0 k� ������e1�t B50A%1r  ��   ����8�}E;�No���|�1Y��3��B�'�  R��#��DTT0 k� ������e1�t B50A%1r  ��   ����8�}E+�Ng���|�1Y��3��B�/�  R��"��DTT0 k� ������e1�t B50A%1r  ��   ����8�}E+�N[���|�0Y��3��B�3�  R��"��DPT0 k� ������e1�t B50A%1r  ��   ����8�|E+�NS���|�0Y��3��B�7�  R��"��DPT0 k� ������e1�t B50A%1r  ��   ����8�|E+��NK�����/Y��3��B�?�  R��!��DPT0 k� ������e1�t B50A%1r  ��   ����8��|E+��NC�����/Y��3��B�C�  R��!��DPT0 k� ������e1�t B50A%1r  ��   ����8��|E+��N;�����.Y��3��B�K�  R�� ��DPT0 k� ������e1�t B50A%1r  ��   ����8��|E,�N3�����-Y��3��B�O�  R�� ��DPT0 k� ������e1�t B50A%1r  ��   ����8� |E,�>'�����-Y��3��B�S�  R�� ��DPT0 k� ������e1�t B50A%1r  ��   ����8�|E,�>�����,Y��3��E,[�  R����J�PT0 k� ������e1�t B50A%1r  ��   ����8�|E,�>�����+Y��3��E,_�  R����J�PT0 k� ������e1�t B50A%1r  ��   ����8�{E,�>�����*Y��3��E,c�  R����J�PT0 k� ������e1�t B50A%1r  ��   ����8�${E,�>�����*Y��3��E,k�  R����J�PT0 k� ������e1�t B50A%1r  ��   ����8�,{E�=������)Y��3��E,o�  R����J�TT0 k� ������e1�t B50A%1r  ��   ����8�8{E�=������(Y��3��E,s�  R����J�TT0 k� ������e1�t B50A%1r  ��   ����8}@{E#�=������'Y��3��E,w�  R����J�TT0 k� ������e1�t B50A%1r  ��   ����8}H{E'�=����� &Y��3��E,{�  R����J�XT0 k� ������e1�t B50A%1r  ��   ����8}PzE/�=����� %Y��3��E,��  R����J�XT0 k� ������e1�t B50A%1r  ��   ����8}\zE3�=�����$Y��3��E��  R�����J�\T0 k� ������e1�t B50A%1r  ��   ����8}dyE7�=�����#Y��3��E��  R�����J�`T0 k� ������e1�t B50A%1r  ��   ����8}lyE?�=�����"Y��3��E��  R�����J�`T0 k� ������e1�t B50A%1r  ��   ����8}txEC�-�����!Y��3��E��  R�����J�dT0 k� ������e1�t B50A%1r  ��   ����8}|xEG�-����� Y��3��E��  R�����J�hT0 k� ������e1�t B50A%1r  ��   ����8}�wEO�-�����Y��3��E��  R�����J�hT0 k� ������e1�t B50A%1r  ��   ����8}�wE�S�-�����Y��3��E��  R�����J�lT0 k� ������e1�t B50A%1r  ��   ����8}�vE�[�-�����Y��3��E��  R�����J�pT0 k� ������e1�t B50A%1r  ��   ����8}�uE�_�-����}Y��3��E�  R�����J�tT0 k� ������e1�t B50A%1r  ��   ����8}�uE�g-����}Y��3��E�  R�����J�xT0 k� ������e1�t B50A%1r  ��   ����8m�tE�k�-����} Y��3��EÀ  R�����J�|T0 k� ������e1�t B50A%1r  ��   ����8m�sD�w�-{���} Y��3��E�ˀ  R�����J�T0 k� ������e1�t B50A%1r  ��   ����8m�sD̃�-w���}$Y��3��E�Ӂ  R�����J�T0 k� ������e1�t B50A%1r  ��   ����8m�rD̋�-o���}(Y��3��E�ہ  R�����J�T0 k� ������e1�t B50A%1r  ��   ����8m�qD̗�-g���}(Y��3��E�߂  R�����JҐT0 k� ����ãe1�t B50A%1r  ��   ����8m�pD̟�c���},Y��3��E��  R��!��JҔT0 k� ����âe1�t B50A%1r  ��   ����8m�oD̟�_���},Y��3��E��  R��!��JҘT0 k� ����áe1�t B50A%1r  ��   ����8m�nP��W���}0Y��3��E���  R��!��JҜT0 k� ����áe1�t B50A%1r  ��   ����8m�mP��S���m0Y��3��E���  R��!��JҤT0 k� �à�Ǡe1�t B50A%1r  ��   ����8m�lP��O���m4Y��3��E��  R��!��Eb�T0 k� ������e1�t B50A%1r  ��   ����8m�kPÌ�K���m4Y��3��E��  R��!��Eb�T0 k� ������e1�t B50A%1r  ��   ����9n jPˍ�G���m8
Y��3��E��  R��!��Eb�T0 k� ����Ýe1�t B50A%1r  ��  ����:^iPӏ�C���m8Y��3��E}�  R��!��Eb�T0 k� �Ý�ǝe1�t B50A%1r  ��   ����;^fP��;���m<Y��3��E}/�  R��!��Eb�T0 k� �ϟ�ӟe1�t B50A%1r  ��   ����<^eP��7���m<Y��3��E}7�  R��1��Eb�T0 k� �נ�۠e1�t B50A%1r  ��  ����=^ dP��3���m<Y��3��E}?�  R��1��K�T0 k� �ߡ��e1�t B50A%1r  ��   ����>�$cP���3���m<Y��3��E}G�  R��1��K�T0 k� ����e1�t B50A%1r  ��   ����?�(bP��/���=?�Y��3��E}O�  R��1��K�T0 k� ����e1�t B50A%1r  ��   ����@�,`P��+���=C�Y��3��E}W�  R��1��K�T0 k� ������e1�t B50A%1r  ��  ����A�4_P��+���=C�Y��3��E}_�  R��1��K�T0 k� �����e1�t B50A%1r  ��   ����B�8^P��'���=C�Y��3��E}g�  R��1��K�T0 k� ����e1�t B50A%1r  ��   ����C�<\P��'���=C�Y��3��E}k�  R��1��K�T0 k� ����e1�t B50A%1r  ��   ����D�D[P'��'���=C�Y��3��Ems�  R��1��K�T0 k� ����e1�t B50A%1r  ��   ����E�LWP3��#���=?�Y��3��Em�  R��1��KT0 k� ���#�e1�t B50A%1r  ��   ����G�TVP;��#���=?�Y��3��Em��  R��A��KT0 k� �'��+�e1�t B50A%1r  ��   ����I�XTPC��#���=?�Y��3��Em��  R��A��KT0 k� �/��3�e1�t B50A%1r  ��   ����K�\RPK�����=?�Y��3��Em��  R��A��KT0 k� �3��7�e1�t B50A%1r  ��   ����M�`PPO�����=?�Y��3��Em��  R��A��K$T0 k� �;��?�e1�t B50A%1r  ��   ����OhNPW�����M?�Y��3��Em��  R��A��K,T0 k� �C��G�e1�t B50A%1r  ��   ����QlMP[�����M;�Y��3��Em��  R��A��K0T0 k� �G��K�e1�t B50A%1r  ��   ����SpKP[�����M;�Y��3��Em��  R��AÏK8T0 k� �K��O�e1�t B50A%1r  ��   ����TtIE�_�M���M;�Y��3��Em��  R��AÍA�<T0 k� �W��[�e1�t B50A%1r  ��   ����V|GE�g�M���M7�Y��3��Em��  R��AǋA�D
T0 k� �c��g�e1�t B50A%1r  ��   ����X�EE�k�M���m7�Y��3��Em��  R��AǉA�H
T0 k� �o��s�e1�t B50A%1r  ��   ����Z�CE�o�M���m7�Y��3��E]��  R��AˇA�P	T0 k� �w��{�e1�t B50A%1r  ��   ����\�BE�w�M���m7�Y��3��E]��  R��QυA�T	T0 k� �����e1�t B50A%1r  �   ����]�@E�w�M���m7�Y��3��E]��  R� QσA�XT0 k� ������e1�t B50A%1r  ��   ����^�<E�w�M���m7�Y��3��E]��  R� Q�A�`T0 k� ������e1�t B50A%1r  ��  ����_�:E�w�M���]7�Y��3��O]��  R� Q�A�dT0 k� ������e1�t B50A%1r  ��   ����`��8E�{�M���]7�Y��3��O]��  R� Q߀EShT0 k� ������e1�t B50A%1r  ��   ����a��7E�{�]�L�]7�Y��3��O]ï  R�Q�ESlT0 k� ������e1�t B50A%1r  ��   ����b��5E��\��L�]7�Y��3��O]ñ  R�Q�ESpT0 k� ������e1�t B50A%1r  �   ����b��3E��\��L�]7�Y��3��O]ǲ  R�Q�EStT0 k� ������e1�t B50A%1r  �   ����b��1E���\��L�]3�Y��3��O]ǳ  R�
��ESxT0 k� ������e1�t B50A%1r �   ����b��/H탲\��L�]3�Y��3��O]Ǵ  R�
��ESxT0 k� ������e1�t B50A%1r ��   ����b �.H탴,��L�]3�Y��3��O]˶  R�
���ES|T0 k� ������e1�t B50A%1r ��   ����b �,H탵,��L�]3�Y�#�3��O]˷  R�
���ES�T0 k� ������e1�t B50A%1r ��   ����b �*H퇶,��L�]3�Y�#�3��O]ϸ  R�
���ES�T0 k� ������e1�t B50A%1r ��   ����b �(H퇸,��L�]/�Y�#�3��O]Ϲ  R�
��ES�T0 k� ������e1�t B50A%1r ��   ����b �&H틹,��L�]/�Y�#�3��O]ӻ  R�
��AS�T0 k� ����e1�t B50A%1r ��  ����b �%H���,��L�]/�Y�#�3��O]Ӽ  R�
��AS�T0 k� ����e1�t B50A%1r ��   ����b �#H���,��L�]/�Y�#�3��O]׽  R�
��AS�T0 k� �/��3�e1�t B50A%1r ��   ����b �!H��� l��L�]/�Y�#�3��O]׾  R�
��AS�T0 k� �?��C�e1�t B50A%1r ��   ����b �H��� l��L�]+�Y�#�3��O]ۿ  R�
��AS�T0 k� �O��S�e1�t B50A%1r ��  ����b �H��� l��L�]+�Y�#�3��O]��  R�
��AS�T0 k� �_��c�e1�t B50A%1r ��   ����b �I�� l��L�]+�Y�'�"s��O]��  R�
��AS�T0 k� �s��w�e1�t B50A%1r ��   ����b  I�� l��L�]+�Y�'�"s��O]��  R�
�#�AS�T0 k� ������e1�t B50A%1r ��  ����b I�� l��L�]+�Y�'�"s��O]��  R�

�'�AS�T0 k� ������e1�t B50A%1r ��   ����b I�� l��L�]+�Y�'�"s��O]��  R�

�+�AS�T0 k� ������e1�t B50A%1r ��   ����b I�� l��L�]'�Y�'�"s��O]��  R�

�+�AS�T0 k� ������e1�t B50A%1r ��   ����b I�� l��L�]'�Y�'�"s��O]��  R�

�/�AS�T0 k� ������e1�t B50A%1r ��   ����b I�� l��L�]'�Y�'�"s��E]��  R�

�3�AS�T0 k� ������e1�t B50A%1r  ��   ����b  I�� l��L�]'�Y�'�"s��E]��  S

�7�AS�T0 k� ������e1�t B50A%1r  ��   ����b $I�� l��L�]'�Y�'�"s��E]��  S

�;�AS�T0 k� ������e1�t B50A%1r  ��   ����b ,I�� l��L�]'�Y�'�"s��E]��  S	
�;�AS�T0 k� ����e1�t B50A%1r  ��   ����b 0
I�� l��L�]#�Y�+�"s��E]��  S	
�?�AS�T0 k� ����e1�t B50A%1r  /�   ����b 4I�� l��L�]#�Y�+�3��E���  S	
�C�AS�T0 k� �+��/�e1�t B50A%1r  ��   ����b 8I�� l��L�]#�Y�+�3��E���  S	
�G�AS�T0 k� �;��?�e1�t B50A%1r  ��   ����b @I�� l��L�]#�Y�+�3��E���  S	
�G�AS�T0 k� �K��O�e1�t B50A%1r  ��   ����b DI�� l��L�]#�Y�+�3��E���  S	
�K�AS�T0 k� �_��c�e1�t B50A%1r  ��   ����b HI�� l��L�]#�a�+�3��E���  S	
�O�AS�T0 k� �o��s�e1�t B50A%1r  ��   ����b P I�� l��L�]#�a�+�3��E���  U�	
�S�AS�T0 k� ������e1�t B50A%1r  ��    ����b�W�I�� l��L�]#�a�+�3��E���  U�	
�S�AS�T0 k� ������e1�t B50A%1r  ��    ����b�[�I�� l��L�]�a�+�3��D=��  U�
�W�AS�T0 k� ������e1�t B50A%1r  ��    ����b�c�I�� l��L�]�a�+�3��D=��  U�
�[�AS�T0 k� ������e1�t B50A%1r  ��    ����b�g�I�� l��L�]�a�+�3��D=��  U�
�[�AS�T0 k� ������e1�t B50A%1r  ��    ����b�o�BM�� l��L�]�a�+�3��D=��  U�
�_�AS�T0 k� ������e1�t B50A%1r  ��    ����b�s�BM�� l��L�]�a�/�"���D=��  U�
�c�AS�T0 k� ������e1�t B50A%1r  ��    ����b�{�BM�� l��L�]�a�/�"���E]��  U�
�c�AS�T0 k� ������e1�t B50A%1r  ��    ����b��BM�� l��L�]�a�/�"���E]��  U�
�g�AS�T0 k� ������e1�t B50A%1r  ��    ����b���BM�� l��L�]�a�/�"���E]��  BM
�k�AS�T0 k� ������e1�t B50A%1r  ��    ����b���BM�� l��L�]�Y�/�"���E]��  BM
�k�AS�T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� l��L�]�Y�/�"���E]��  BM
�o�AS�T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� l��L�]�Y�/�"���E]��  BM
�o�AS� T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� l�L�]�Y�/�"���E]��  BM
�s�AS� T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� l{�L�]�Y�/�"���E]��  BM
�s�AS� T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� lw�L�]�Y�/�"���E]��  BM
�w�AS� T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� lw�L�]�Y�/�"���A]��  BM
�{�AS� T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� ls�L�]�Y�/�3��A]��  BM
�{�AS� T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� lo�L�]�Y�/�3��A]��  BM
��AS� T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� lo�L�]�Y�/�3��A]��  BM
��AS� T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� lo�L�]�Y�/�3��A]��  BM
҃�AS� T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� lo�L�]�a�/�3��A]��  BM
҃�AS� T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� lo�L�]�a�/�3��A]��  BM
҇�AS� T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� lo�L�]�a�+�3��A]��  BM
҇�AS� T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� lo�L�]�a�+�3��A]��  BM
ҋ�AS� T0 k� ���#�e1�t B50A%1r  ��    ����b ��BM�� lo�L�]�a�+�3��A]��  BM
ҋ�AS� T0 k� �#��'�e1�t B50A%1r  ��    ����b ��BM�� lk�L�]�a�'�3��A]��  BM
ҏ�AS� T0 k� �'��+�e1�t B50A%1r  ��    ����b ��BM�� lk�L�]�a�'�3��A]��  BM 
ҏ�AS� T0 k� �+��/�e1�t B50A%1r  ��    ����b ��BM�� lk�L�]�a�'�3��A]��  BM 
ғ�AS� T0 k� �/��3�e1�t B50A%1r  ��    ����b ��BM�� lk�L�]�a�#�3��A]��  BM 
ғ�AS� T0 k� �3��7�e1�t B50A%1r  ��    ����b ��BM�� lg�L�]�a�#�3��A]��  BM 
ғ�AS� T0 k� �;��?�e1�t B50A%1r  ��    ����b ��BM�� lg�L�]�a�#�3��A]��  BM 
җ�AS��T0 k� �?��C�e1�t B50A%1r  ��    ����b ��BM�� lg�L�]�Y�#�4�A]��  BM 
җ�AS��T0 k� �C��G�e1�t B50A%1r  ��    ����b ��BM�� lc�L�]�Y��4�A]��  BM 
қ�AS��T0 k� �G��K�e1�t B50A%1r  ��    ����b �BM�� lc�L�]�Y��4�A]��  BM 
қ�AS��T0 k� �K��O�e1�t B50A%1r  ��    ����b �BM�� lc�L�]�Y��4�A]��  BM 
ҟ�AS��T0 k� �O��S�e1�t B50A%1r  ��    ����b �BM�� lc�L�]�Y��4�A]��  BM 
ҟ�AS��T0 k� �S��W�e1�t B50A%1r  ��    ����b �BM�� l_�L�]�Y��4�A]��  BM 
ҟ�AS��T0 k� �W��[�e1�t B50A%1r  ��    ����b �BM�� l_�L�]�Y��4�A]��  BM 
ң�AS��T0 k� �[��_�e1�t B50A%1r  ��    ����b �BM�� l_�L�]�Y��4�A]��  BM 
ң�AS��T0 k� �_��c�e1�t B50A%1r  ��    ����b �BM�� l_�L�]�Y��4�A]��  BM 
ҧ�AS��T0 k� �c��g�e1�t B50A%1r  ��    ����b �BM�� l[�L�]�Y��4�A]��  BM$
ҧ�AS��T0 k� �g��k�e1�t B50A%1r  ��    ����b #�BM�� l[�L�]�Y��4�A]��  BM$
ҧ�AS��T0 k� �k��o�e1�t B50A%1r  ��    ����b #�BM�� l[�L�]�Y��4�A]��  BM$
ҫ�AS��T0 k� �k��o�e1�t B50A%1r  ��    ����b '�BM�� l[�L�]�Y��4�A]��  BM$
ҫ�AS��T0 k� �o��s�e1�t B50A%1r  ��    ����b +�BM�� lW�L�]�Y��4�A]��  BM$
ҫ�AS��T0 k� �s��w�e1�t B50A%1r  ��    ����b /�BM�� lW�L�]�Y��4�A]��  BM$
ү�AS��T0 k� �w��{�e1�t B50A%1r  ��    ����b 3�BM�� lW�L�]�Y��4�A]��  BM$
ү�AS��T0 k� �{���e1�t B50A%1r  ��    ����b 7�BM�� lW�L�]�Y��4�A]��  BM$
ү�AS��T0 k� �����e1�t B50A%1r  ��    ����b ;�BM�� lS�L�]�Y��4�A]��  BM$
ҳ�AS��T0 k� ������e1�t B50A%1r  ��    ����b ;�BM�� lS�L�]�Y��4�A]��  BM$
ҳ�AS��T0 k� ������e1�t B50A%1r  ��    ����b ?�BM�� lS�L�]�Y��4�A]��  BM$
ҳ�AS��T0 k� ������e1�t B50A%1r  ��    ����b C�BM�� lS�L�]�Y��4�A]��  BM$
ҷ�AS��T0 k� ������e1�t B50A%1r  ��    ����b G�BM�� lS�L�]�Y��4�A]��  BM$
ҷ�AS��T0 k� ������e1�t B50A%1r  ��    ����b G�BM�� lS�L�]�Y��4�A]��  BM$
ҷ�AS��T0 k� ������e1�t B50A%1r  ��    ����b K�BM�� lS�L�]�Y��4�A]��  BM$
һ�AS��T0 k� ������e1�t B50A%1r  ��    ����b O�BM�� lS�L�]�Y��4�A]��  BM$
һ�AS��T0 k� ������e1�t B50A%1r  ��    ����b S�BM�� lS�L�]�Y��4�A]�   BM$
һ�AS��T0 k� ������e1�t B50A%1r  ��    ����b S�BM�� lO�L�]�Y��4�A]�  BM(
һ�AS��T0 k� ������e1�t B50A%1r  ��    ����b W�BM�� lO�L�]�Y��4�A]�  BM(
ҿ�AS��T0 k� ������e1�t B50A%1r  ��    ����b [�BM�� lO�L�]�Y��4�A]�  BM(
ҿ�AS��T0 k� ������e1�t B50A%1r  ��    ����b [�BM�� lO�L�]�Y��4�A]�  BM(
ҿ�AS��T0 k� ������e1�t B50A%1r  ��    ����b _�BM�� lO�L�]�Y��4�A]�  BM(
�ØAS��T0 k� ������e1�t B50A%1r  ��    ����b c�BM�� lK�L�]�Y��4�A]�  BM(
�ØAS��T0 k� ������e1�t B50A%1r  ��    ����b c�BM�� lK�L�]�Y��4�A]�  BM(
�ØAS��T0 k� ������e1�t B50A%1r  ��    ����b g�BM�� lK�L�]�Y��4�A]�  BM(
�ÙAS��T0 k� ������e1�t B50A%1r  ��    ����b k�BM�� lK�L�]�Y��4�A]�  BM(
�ǙAS��T0 k� ������e1�t B50A%1r  ��    ����b k�BM�� lK�L�]�Y��4�A]�  BM(
�ǙAS��T0 k� ������e1�t B50A%1r  ��    ����b o�BM�� lG�L�]�Y��4�A]�  BM(
�ǙAS��T0 k� ������e1�t B50A%1r  ��    ����b o�BM�� lG�L�]�Y��4�A]�  BM(
�ǙAS��T0 k� ������e1�t B50A%1r  ��    ����b s�BM�� lG�L�]�Y��4�A]�  BM(
�˙AS��T0 k� ������e1�t B50A%1r  ��    ����b w�BM�� lG�L�]�Y��4�A]�  BM(
�˙AS��T0 k� ����óe1�t B50A%1r  ��    ����b w�BM�� lC�L�]�Y���4�A]�  BM(
�˙AS��T0 k� ����óe1�t B50A%1r  ��    ����b {�BM�� lC�L�]�Y���4�A]�  BM(
�˙AS��T0 k� �ò�ǲe1�t B50A%1r  ��    ����b {�BM�� lC�L�]�Y���4�A]�	  BM(
�ϚAS��T0 k� �ǲ�˲e1�t B50A%1r  ��    ����b �BM�� lC�L�]�Y���4�A]�	  BM(
�ϚAS��T0 k� �Ǳ�˱e1�t B50A%1r  ��    ����b �BM�� lC�L�]�Y���4�A]�	  BM(
�ϚAS��T0 k� �˱�ϱe1�t B50A%1r  ��    ����b ��BM�� l?�L�]�Y���4�A]�
  BM(
�ϚAS��T0 k� �˰�ϰe1�t B50A%1r  ��    ����b ��BM�� l?�L�]�Y���4�A]�
  BM(
�ϚAS��T0 k� �ϰ�Ӱe1�t B50A%1r  ��    ����b ��BM�� l?�L�]�Y���4�A]�  BM(
�ӚAS��T0 k� �ϯ�ӯe1�t B50A%1r  ��    ����b ��BM�� l?�L�]�Y���4�A]�  BM(
�ӚAS��T0 k� �ӯ�ׯe1�t B50A%1r  ��    ����b ��BM�� l?�L�]�Y���4�A]�  BM,
�ӚAS��T0 k� �Ӯ�׮e1�t B50A%1r  ��    ����b ��BM�� l;�L�]�Y���4�A]�  BM,
�ӚAS��T0 k� �׮�ۮe1�t B50A%1r  ��    ����b ��BM�� l;�L�]�Y���4�A]�  BM,
�ӚAS��T0 k� �׭�ۭe1�t B50A%1r  ��    ����b ��BM�� l8 L�]�Y���4�A]�  BM,
�ךAS��T0 k� �ۭ�߭e1�t B50A%1r  ��    ����b ��BM�� l8 L�]�Y���4�A]�  BM,
�כAS��T0 k� �۬�߬e1�t B50A%1r  ��    ����b ��BM�� l8 L�]�Y���4�A]�  BM,
�כAS��T0 k� �߬��e1�t B50A%1r  ��    ����b ��BM�� l8L�]�Y���4�A]�  BM,
�כAS��T0 k� �߬��e1�t B50A%1r  ��    ����b ��BM�� l4L�]�Y���4�A]�  BM,
�כAS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� l4L�]�Y���4�A]�  BM,
�ۛAS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� l4L�]�Y���4�A]�  BM,
�ۛAS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� l4L�]�Y���4�A]�  BM,
�ۛAS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� l4L�]�Y���4�A]�  BM,
�ۛAS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� l4L�]�Y���4�A]�  BM,
�ۛAS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� l4L�]�Y���4�A]�  BM,
�ۛAS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� l4L�]�Y��3��A]�  BM,
�ߛAS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� l0L�]�Y��3��A]�  BM,
�ߛAS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� l0L�]�Y��3��A]�  BM,
�ߛAS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�� l0L�]�Y��3��A]�  BM,
�ߜAS��T0 k� �����e1�t B50A%1r  ��    ����b ��BM�� l0L�]�Y��3��A]�  BM,
�ߜAS��T0 k� �����e1�t B50A%1r  ��    ����b ��BM�� l0L�]�Y��3��A]�  BM,
�ߜAS��T0 k� �����e1�t B50A%1r  ��    ����b ��BM�� l0L�]�Y��3��A]�  BM,
�ߜAS��T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� l0L�]�Y��3��A]�  BM,
��AS��T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� l0L�]�Y��3��A]�  BM,
��AS��T0 k� ������e1�t B50A%1r  ��    ����b ��BM�� l,L�]�Y��3��A]�  BM,
��AS��T0 k� ������e1�t B50A%1r  ��    ����b ��BM�  l,L�]�Y��3��A]�  BM,
��AS��T0 k� ������e1�t B50A%1r  ��    ����b ��BM�  l,L�]�Y��3��A]�  BM,
��AS��T0 k� �����e1�t B50A%1r  ��    ����b ��BM�  l,L�]�Y��3��A]�  BM,
��AS��T0 k� �����e1�t B50A%1r  ��    ����b ��BM�  l,L�]�Y��3��A]�  BM,
��AS��T0 k� �����e1�t B50A%1r  ��    ����b ��BM�  l,L�]�Y��3��A]�  BM,
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM�  l,L�]�Y��3��A]�  BM,
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM� l,L�]�Y��3��A]�  BM,
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM� l,L�]�Y��3��A]�  BM,
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM� l(L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM� l(	L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM� l(	L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM� l(	L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ��BM� l(
L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b çBM� l(
L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b æBM� l(
L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b æBM� l(L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b æBM� l$L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ǦBM� l$L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ǥBM� l$L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ǥBM� l$L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ǥBM� l$L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ˥BM� l$L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ˤBM� l$L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ˤBM� l$L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ˤBM� l L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ϤBM� l L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ϤBM� l L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ϣBM� l L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ϣBM� l L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ӣBM� l L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ӣBM� l L�]�Y��3��A]�  BM0
��AS��T0 k� ����e1�t B50A%1r  ��    ����b ӣBM� l L�]�Y��3��A]�  BM0
��AS��T0 k� ���#�e1�t B50A%1r  ��    ����b ӢBM� l L�]�Y��3��A]�  BM0
��AS��T0 k� ���#�e1�t B50A%1r  ��    ����b ӢBM� lL�]�Y��3��A]�  BM0
��AS��T0 k� ���#�e1�t B50A%1r  ��    ����b עBM� lL�]�Y��3��A]�  BM0
��AS��T0 k� ���#�e1�t B50A%1r  ��    ����b עBM� lL�]�Y��3��A]�  BM0
��AS��T0 k� ���#�e1�t B50A%1r  ��    ����b עBM� lL�]�Y��3��A]�  BM0
��AS��T0 k� �#��'�e1�t B50A%1r  ��    ����b עBM� lL�]�Y��3��A]�  BM0
��AS��T0 k� �#��'�e1�t B50A%1r  ��    ����b סBM� lL�]�Y��3��A]�  BM0
��AS��T0 k� �#��'�e1�t B50A%1r  ��    ����b ۡBM� lL�]�Y��3��A]�  BM0
��AS��T0 k� �#��'�e1�t B50A%1r  ��    ����b ۡBM� lL�]�Y��3��A]�  BM0
��AS��T0 k� �#��'�e1�t B50A%1r  ��    ����b ۡBM� lL�]�Y��3��A]�  BM0
��AS��T0 k� �'��+�e1�t B50A%1r  ��    ����b ۡBM� lL�]�Y��3��A]�  BM0
��AS��T0 k� �'��+�e1�t B50A%1r  ��    ����b ۡBM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �'��+�e1�t B50A%1r  ��    ����b ߠBM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �'��+�e1�t B50A%1r  ��    ����b ߠBM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �'��+�e1�t B50A%1r  ��    ����b ߠBM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �+��/�e1�t B50A%1r  ��    ����b ߠBM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �+��/�e1�t B50A%1r  ��    ����b ߠBM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �+��/�e1�t B50A%1r  ��    ����b ߠBM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �+��/�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �+��/�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �+��/�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �/��3�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �/��3�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM0
���AS��T0 k� �/��3�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �/��3�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �/��3�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �/��3�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �/��3�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �3��7�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �3��7�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �3��7�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �3��7�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �3��7�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �3��7�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �3��7�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �3��7�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �7��;�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �7��;�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �7��;�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �7��;�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �7��;�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �7��;�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �7��;�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�  BM4
���AS��T0 k� �7��;�e1�t B50A%1r  ��    ����b �BM� lL�]�Y��3��A]�   BM4
���AS��T0 k� �;��?�e1�t B50A%1r  ��    ����bhuD����������Y|/�3��I��  C�d�g�FO�T0 k� ������e1�t B50A%1r  ��7   ����9`uD����������Y|/�3��I��  C�e�c�FO�T0 k� ������e1�t B50A%1r  ��7   ����8XtD���� �����Y|/�3��I���  C�f�c�FK�T0 k� ������e1�t B50A%1r  ��7   ����8LtD����� �����Y|/�3��I���  C�h�_�E�K�T0 k� ������e1�t B50A%1r  ��7   ����8DtD����� �����Y|/�3��I���  C�i�_�E�G�T0 k� ������e1�t B50A%1r  ��7   ����8<sC����� �����Y|/�3��I���  E^|j�[�E�G�T0 k� ������e1�t B50A%1r  ��7   ����84sC����� �����Y|/�3��I���  E^tk�[�E�G�T0 k� ������e1�t B50A%1r  ��7   ����8(sC����� �����Y|/�3��I���  E^pm�W�E�C�T0 k� ������e1�t B50A%1r  ��7   ����8 rC����� �����Y|/�3��I���  E^hn�S�E�C�T0 k� ������e1�t B50A%1r  ��7   ����8rC����� �����Y|/�3��I���  E^`o�O�E�C�T0 k� ������e1�t B50A%1r  ��7   ����8rC��������L��Y|/�3��I���  E^\p�K�E�C�T0 k� ������e1�t B50A%1r  ��7   ����8rC��������L��Y|/�3��I���  E^Tq�G�E�C�T0 k� ������e1�t B50A%1r  ��7   ����8�qC�w�������L��Y|/�3��I���  E^Ls�C�E�C�T0 k� ������e1�t B50A%1r  ��7   ����8�qC�o�������L��Y|/�3��I���  E^Dt�?�B�C�T0 k� ������e1�t B50A%1r  ��7   ����8��qC�g�������L��Y|/�3��I���  EN@u�;�B�C�T0 k� ������e1�t B50A%1r  ��7   ����8��pC�_�N�������Y|/�3��I���  EN8v�7�B�G�T0 k� ������e1�t B50A%1r  ��7   ����8��pC�W�N�������Y|/�3��I���  EN0w�3�B�G�T0 k� ������e1�t B50A%1r  ��7   ����8��pC�O�N{������Y|/�3��I���  EN(x�+�B�G�T0 k� ������e1�t B50A%1r  ��7   ����8��oC�G�Ns������Y|/�3��I���  EN x�'�B�K�T0 k� ������e1�t B50A%1r  ��7   ����8��oC�?�Nk������Y|/�3��I���  ENy#�B�K�T0 k� ������e1�t B50A%1r  ��7   ����8�oC�7�N_������Y|/�3��I���  ENz�B�O�T0 k� ������e1�t B50A%1r  ��7   ����8�nC�/�NW������Y|/�3��I���  EN{�B�O�T0 k� ������e1�t B50A%1r  ��7   ����8�nC�'�NO������Y|/�3��E���  EN{�B�S�T0 k� ������e1�t B50A%1r  ��7   ����8��nC��NC������Y|/�3��E���  EM�|�B�S�T0 k� ������e1�t B50A%1r  ��7   ����8��mC��N;������Y|/�3��E���  C��|�B�W�T0 k� ������e1�t B50A%1r  ��7   ����8��mC��>3������Y|/�3��E��  C��}��B�[�T0 k� ������e1�t B50A%1r  ��7   ����8��mC��>'������Y|/�3��E��  C��}��B�_�T0 k� ������e1�t B50A%1r  ��7   ����8�xmC���>������Y|/�3��E���  C��~��B�c�T0 k� ������e1�t B50A%1r  ��7   ����8�plD��>������Y|/�3��E���  C��~��B�c�T0 k� ������e1�t B50A%1r  ��7   ����8�dlD��>������Y|/�3��E���  C��~��B�g�T0 k� ������e1�t B50A%1r  ��7   ����8�\lD��>������Y|/�3��E���  C����E�k�T0 k� ������e1�t B50A%1r  ��7   ����8�TkD��=�������Y|/�3��E���  C����E�o�T0 k� ������e1�t B50A%1r  ��7   ����8�LkD��=�������Y|/�3��Em��  C����E�s�T0 k� ������e1�t B50A%1r  ��7   ����8�DkE���=�������Y|/�3��Em��  C����E�w�T0 k� ������e1�t B50A%1r  ��7   ����8�0jE��=�������Y|/�3��Em��  C����E��T0 k� ������e1�t B50A%1r  ��7   ����8�(jE��=�������Y|/�3��Em��  C����D߃�T0 k� �����e1�t B50A%1r  ��7   ����8  jE��=�������Y|/�3��Em��  C����D߇�T0 k� �w��{�e1�t B50A%1r  ��7   ����8 iE��-�������Y|/�3��Em��  C����Dߋ�T0 k� �o��s�e1�t B50A%1r  ��7   ����8 iE��-�������Y|/�3��Em��  C����Dߓ�T0 k� �g��k�e1�t B50A%1r  ��7   ����8 iE��-�������Y|/�3��Em��  C�x��Dߗ�T0 k� �\ �` e1�t B50A%1r  ��7   ����8�hE��-�������Y|/�3��Em��  C�p��Dߛ�T0 k� �X�\e1�t B50A%1r  ��7   ����8�hE��-�������Y|/�3��A��  C�d~�w�Dߟ�T0 k� �P�Te1�t B50A%1r  ��7   ����8�hD>{�-�������Y|/�3��A�{�  C�\~�o�Dߣ�T0 k� �L�Pe1�t B50A%1r  ��7   ����8�gD>s�-�������Y|/�3��A�w�  C�T~�g�D߫�T0 k� �D�He1�t B50A%1r  ��7   ����8�gD>k�-�������Y|/�3��A�o�  C�L}�[�D߯�T0 k� �@�De1�t B50A%1r  ��7   ����8��gD>c���������Y|/�3��A�k�  C�D}�S�D߳�T0 k� �8�<e1�t B50A%1r  ��7   ����8��gD>[��������Y|/�3��Emc�  C�<}�K�D߻�T0 k� �4�8e1�t B50A%1r  ��7   ����8߼fE^S��������Y|/�3��Em_�  C�4|�?�D��T0 k� �,	�0	e1�t B50A%1r  ��7   ����8ߴfE^K��������Y|/�3��Em[�  C�,|�7�D���T0 k� �(
�,
e1�t B50A%1r  ��7   ����8ߤeE^;�������Y|/�3��EmL  C�{B#�D���T0 k� �� e1�t B50A%1r  ��7   ����8ߘeE^3�-����Y|/�3��EmD  C�{B�D���T0 k� ��e1�t B50A%1r  ��7   ����8ߐeE^+�-{����Y|, 3��EmD  C�zB�E���T0 k� ��e1�t B50A%1r  ��7   ����8߈eE^#�-w���  Y|, 3��Em@  C�zB�E���T0 k� ��e1�t B50A%1r  ��7   ����8߀dE^�-s��#��Y|, 3��Em<  C��yA��E���T0 k� ��e1�t B50A%1r  ��7   ����8�tdE^�-o��+��Y|,3��Em8  C��yA��E���T0 k� � �e1�t B50A%1r  ��7   ����8�ldEN�-k��+��Y|,3��E]4	  C��xA��E���T0 k� ��e1�t B50A%1r  ��7   ����8�dcEN�-k��+��Y|,3��E]0  C��xA��E���T0 k� ��e1�t B50A%1r  ��7   ����8�\cEM��-k��/��Y|,3��E](  C��wA��E��T0 k� � �e1�t B50A%1r  ��7   ����8�TcEM��-k��/��Y|,3��E]$  C��wA��E��T0 k� � �e1�t B50A%1r  ��7   ����8�@bEM��o��/��Y|,3��E]  C��uA��J@�T0 k� ����e1�t B50A%1r  ��7   ����8�8bEM��o��/��Y|,3��E]  C̼u1��J@�T0 k� ����e1�t B50A%1r  ��G   ����8�0bEM��o��3�L�Y|,3��E]  C̴t1��J@'�T0 k� ����e1�t B50A%1r  ��G   ����8�$aEM��s��3�L�Y|,3��G�  C̬t1��J@/�T0 k� ����e1�t B50A%1r  ��G   ����8?aEM��s��3�L�Y|,3��G�   C̤s1��J@7�T0 k� ����e1�t B50A%1r  ��G   ����8?aEM���w��3�L�Y|,"���G��  C̜r1��E;�T0 k� ����e1�t B50A%1r  ��G   ����8?aE=���t�3�L�	Y|,"���G��  C̔r1��EC�T0 k� ����e1�t B50A%1r  ��G   ����8? `E=���x�3�L�	Y|,	"���G��  C��q1��EK�T0 k� ����e1�t B50A%1r  �G   ����8>�`E=�����7�L�Y|,
"���G��  C�|o1s�E[�T0 k� ����e1�t B50A%1r ��O   ����8>�_E=�����7�L�Y|,"���G��!  C�to1k�Ec�T0 k� ����e1�t B50A%1r ��O   ����8>�_E=����	�7�L�Y|,"���G��"  C�ln1c�Ek�T0 k� ��
��
e1�t B50A%1r ��O   ����8>�_E=����;�L�Y|0"���G��$  ELdm�_�Es�T0 k� ����e1�t B50A%1r ��O   ����8>�^CMw���;�L�Y|0"���G��%  EL\l�W�E�w�T0 k� �x�|e1�t B50A%1r ��O   ����8>�^CMo���;�<�Y|0"���G��&  ELXl�O�E��T0 k� �l�pe1�t B50A%1r ��O   ����8>�^CMg���?�<�Y|0"���G��(  ELPk�G�E���T0 k� �`�de1�t B50A%1r ��O   ����8N�]CM[���C�<�Y|03��G�*  EL@i�7�E���T0 k� �O��S�e1�t B50A%1r ��O   ����8N�]CMS���C�<�Y�03��G�,  EL8h�3�E���T0 k� �C��G�e1�t B50A%1r ��?   ����8N�\E�K���C�\�Y�03��G�-  EL0h�+�E���T0 k� �7��;�e1�t B50A%1r ��?   ����8N�\E�G��MG�\�Y�03��G�.  E<(g�#�E���T0 k� �+��/�e1�t B50A%1r	 ��?   ����8N�[E�?��MG�\�Y�03��G�/  E< f��Dг�T0 k� ���#�e1�t B50A%1r	 ��?   ����8^|[E�7��MG�\|Y�03��G�1  E<e��Dл�T0 k� ����e1�t B50A%1r
 ��?   ����8^t[E�/��MK�\xY�03��G�2  E<d��D���T0 k� ����e1�t B50A%1r
 ��?   ����8^lZE�'���MK�ltY�03��G�3  E<c��D���T0 k� �����e1�t B50A%1r
 ��?   ����8^`ZE���� �K�llY�03��G�4  E<b��D���T0 k� ������e1�t B50A%1r ��?   ����8^XZE����"�O�lhY�03��G�5  E< a��F ��T0 k� ������e1�t B50A%1r �?   ����8^PYE����#�O�ldY�0"s��G�6  E;�_1�F ��T0 k� ������e1�t B50A%1r
 ��?   ����8^HYE����$�O�l`Y�0"s��G�8  E;�^1�F ��T0 k� ������e1�t B50A%1r
 ��?   ����8^@YE����&�L l\Y�0"s��G�9  E;�]1�F ��T0 k� ������e1�t B50A%1r	 ��?   ����8�4XE���� '�L\XY�0
"s��G�:  E;�\0��F ��T0 k� �����e1�t B50A%1r ��?   ����8�$XE����)�P\PY�0
"s��E\t<  E+�Y0��F ��T0 k� ����e1�t B50A%1r ��?   ����8�WE����*�P\PY�0
"s��E\p=  E+�X ��F ��T0 k� ����e1�t B50A%1r ��?   ����8�WE���� ,�L\LY�0
"s��E\l>  E+�W ��F ��T0 k� ����e1�t B50A%1r ��?   ����8^WE����,-�L<HY�0
"s��E\h?  E+�U ��E���T0 k� ����e1�t B50A%1r ��?   ����8^ VE���~4.�L	<D Y�0
"s��E\`@  E+�T ��E���T0 k� ����e1�t B50A%1r ��?   ����8]�UEܿ�~D/�L<<!Y�0	"s��ELXA  E+�Q ��E���T0 k� ����e1�t B50A%1r ��?   ����8]�UEܷ�~P0�L<8"Y�0	3��ELPB  E+�P!�E�� T0 k� ����e1�t B50A%1r  ��?   ����8]�UEܯ�~X1�H<4#Y�4	3��ELLC  E+�N!�E�� T0 k� ���#�e1�t B50A%1r  ,�?   ����8]�TEܫ�~`1�H<0$Y�4	3��ELHD  E+�M!�E��T0 k� �#��'�e1�t B50A%1r  ��?   ����8]�TEܣ�~h2�D<0%Y�4	3��EL@D  E+�K�E��T0 k� �'��+�e1�t B50A%1r  ��?   ����8]�TE��~t2�D<,&Y�4	3��EL<E  E+�J�E��T0 k� �'��+�e1�t B50A%1r ��?   ����8M�SE��~�3�<,$(Y�4	3��EL0F  E�G�E��T0 k� �/��3�e1�t B50A%1r ��?   ����8M�SE��~�4�<,$)Y�43��EL(F  E�F�E��T0 k� �3��7�e1�t B50A%1r ��?   ����8M�SE�{�~�4�8, *Y�43��EL$F  E�D
A�E��T0 k� �7��;�e1�t B50A%1r ��?   ����8M�RE�s�n�4�4,+Y�43��E<G  E�C
A�E��T0 k� 7��;�e1�t B50A%1r ��?   ����8M�RE�k�n�4�0,,Y�43��E<G  E�A
A�E��T0 k� ;��?�e1�t B50A%1r ��?   ����8M�RE�c�n�4�0,-Y�43��E<G  B��@
A�E��T0 k� ?��C�e1�t B50A%1r ��?   ����8MpQE�S�n�4�(,0Y�43��E<G  B��=1�E��T0 k� G��K�e1�t B50A%1r ��?  ����8MhQE�K�>�4�$,1Y|43��CL G  B��<1�E��T0 k� �G��K�e1�t B50A%1r $�?   ����8M`QE�C�>�4� ,2Y|43��CK�G  B��;1�E��T0 k� �K��O�e1�t B50A%1r ��?   ����8MXPE�7�>�4�,3Y|43��CK�G  E�91#�J� T0 k� �K��O�e1�t B50A%1r ��?   ����8MDPE�'�>�3� 5Y|43��CK�F  E�7A'�J�T0 k� �K��O�e1�t B50A%1r ��?   ����8=<PE��>�3� 7Y|43��CK�F  E�5A+�J�T0 k� ,O��S�e1�t B50A%1r ��?   ����8=4PE��>�3�!8Y|43��CK�E  E�4A/�J�T0 k� ,O��S�e1�t B50A%1r ��?  ����8=(PE��>�2�!9Y|43��CK�E  E�3A/�J�	T0 k� ,O��S�e1�t B50A%1r ��?   ����8= PE��? 2� ":Y|43��CK�D  E�2A3�J�	T0 k� ,O��S�e1�t B50A%1r ��?   ����8=PE���?1��"<Y|43��CK�C  E��0A;�J�
T0 k� �S��W�e1�t B50A%1r ��?   ����8=QE���?0��#=Y�43��CK�B  E��/A?�J� 
T0 k� �S��W�e1�t B50A%1r ��?   ����8<�QE���O0��#>Y�43��E;�A  E��.QC�J�(
T0 k� �W��[�e1�t B50A%1r ��?   ����8<�QE���O/��#?Y�43��E;�A  E��-QG�J�,T0 k� �W��[�e1�t B50A%1r ��?   ����8<�RE���O .��#�@Y�4 3��E;�@  E��,QK�J�0T0 k� �W��[�e1�t B50A%1r ��?   ����8<�SF��O(-��#�BY�3�3��E;�>  E��*QW�J�<T0 k� <[��_�e1�t B50A%1r  ��?   ����8,�SF��O,,��#�CY�3�3��E;�=  E��)
�[�J�@T0 k� <[��_�e1�t B50A%1r  ��?   ����8,�TF��O0+��#�DY�3�3��E;�<  E��)
�_�J�HT0 k� <[��_�e1�t B50A%1r  .�?   ����8,�UF��O4*��#�EY�3�3��E;�;  E��(
�g�J�LT0 k� <[��_�e1�t B50A%1r  ��?  ����8,�VF��o8)��"�EY�3�3��E;�9  D۬(
�k�J�TT0 k� <_��c�e1�t B50A%1r  ��?   ����8,�VF��o<(��"�FY�3�3��E;�8  D۰'
�o�J�XT0 k� �_��c�e1�t B50A%1r  ��?   ����8,�WF��o@'��"�GY�3�3��E;�7  D۰'
�w�J�`T0 k� �_��c�e1�t B50A%1r  ��?   ����8,�YF��oD%�!�HY�3�3��E+�4  D۸&
у�J�lT0 k� �c��g�e1�t B50A%1r  ��?   ����8,�ZF��oH$� � IY�3�3��E+�3  Dۼ%
ы�J�tT0 k� �c��g�e1�t B50A%1r  ��?   ����8,�[F��oL"� � IY�/�3��E+�1  D��%
я�J�|T0 k� �c��g�e1�t B50A%1r  ��?   ����8,�\F��oL!��$IY�/�3��E+|0  D��%
ї�JрT0 k� �g��k�e1�t B50A%1r  ��?   ����8,�]E���oP ��(JY�/�3��E+|/  D��%
��JшT0 k� �g��k�e1�t B50A%1r  ��?   ����8|^E���oPܰ�(JY�/�3��E+x-  D��$
��JѐT0 k� �g��k�e1�t B50A%1r  ��?   ����8p`E���oTܨ�,KY�/�3��E+t*  D��$
��JѠT0 k� �k��o�e1�t B50A%1r  ��?  ����8lbE���_Xܨ�0KY�/�3��B�p)  D��$
��JѨT0 k� �k��o�e1�t B50A%1r  ��?   ����8dcE���_Xܨ�4KY�/�3��B�p'  D��$���JѰT0 k� �k��o�e1�t B50A%1r  ��?   ����8�`dE���_Xܤ�8LY�/�3��B�l%  D��$���JѸT0 k� �k��o�e1�t B50A%1r  ��?   ����8�\eE���_Xܤ�8LY�/�3��B�l$  D��$���J��T0 k� �o��s�e1�t B50A%1r  ��?   ����8�XfE���_Xܤ|<LY�+�3��B�l"  D��%���J��T0 k� �o��s�e1�t B50A%1r  ��?   ����8�TgB���_Xܠ|@LY�+�3��B�h!  D��%���J��T0 k� �o��s�e1�t B50A%1r  ��?   ����8�LiB���_X�|DLY�+�3��B�l  D��%���J��T0 k� �s��w�e1�t B50A%1r  ��?   ����8�LjB���_X�|HLY�+�3��B�l  D��%���J��T0 k� �s��w�e1�t B50A%1r  ��?   ����8�HkB����X��LLY�'�3��B�p  D� &���J��T0 k� �s��w�e1�t B50A%1r  ��?   ����8�DlB����T��LKY�'�3��B�p  D�&���J��T0 k� �w��{�e1�t B50A%1r  ��?   ����8�Dn@���T��PKY�'�3��B�t  D�&���C� T0 k� �w��{�e1�t B50A%1r  ��?   ����8�@o@���P		���TKY�'�3��Ct  D�'���C�T0 k� �w��{�e1�t B50A%1r  ��   ����8�<q@���L	���XJY�'�3��Cx  D�(Q��C�T0 k� �{���e1�t B50A%1r  ��   ����8�<r@���L	���\JY�'�3��C|  D� (Q��C�T0 k� �{���e1�t B50A%1r  ��   ����8�<sE����H	���\JY�'�3��C|  D�$)Q��C�$T0 k� �{���e1�t B50A%1r  ��   ����8�<tE����D	���`IY�'�3��C�  D�()Q��C�(T0 k� �{���e1�t B50A%1r  ��   ����8�<uE����@
��dIY�'�3��C�	  D�0*Q��C�0T0 k� �����e1�t B50A%1r  ��   ����8�<vE����?�
�
�dHY�'�3��E��  D�4+Q��C�4T0 k� �����e1�t B50A%1r  ��   ����8�<wE����;�
�	�hGY�'�3��E��  D�<+Q��C�8T0 k� �����e1�t B50A%1r  ��   ����8�<yE����3�
��lFY�'�3��E��  D�H-���C�@T0 k� ������e1�t B50A%1r  ��   ����8�<zE����/�	���pDY�'�3��E���  EL.���C�DT0 k� ������e1�t B50A%1r  ��   ����8�<{E����+�	���pBY�'�3��E���  ET.���C�HT0 k� ������e1�t B50A%1r  ��   ����8�@|E����#�	���t?Y�#�3��E���  E\/���C�LT0 k� ������e1�t B50A%1r  ��   ����8�@~E�����	���t?Y�#�3��E���  E\/���C�PT0 k� ������e1�t B50A%1r  �   ����8�@E�����	��|x>Y�#�3��E+��  E`.���C�TT0 k� ������e1�t B50A%1r  ��   ����8�D�E�����
�|�>Y�#�3��E+��  R�d-���C�TT0 k� ������e1�t B50A%1r  ��   ����8�HE�����
�|�=Y�#�3��E+��  R�h-���C�XT0 k� ������e1�t B50A%1r  ��   ����8�LE�����
�|�<Y�#�3��E+��  R�l,���C�XT0 k� ������e1�t B50A%1r  ��   ����8�PE������
�|�<Y�#�3��E+��  R�p,���C�\T0 k� ������e1�t B50A%1r  ��   ����8�PE�����
�|�;Y�#�3��B��  R�t+���C�\T0 k� ������e1�t B50A%1r  ��   ����8�XE�����	��|�:Y�#�3��B��  R�x+���C�\T0 k� ������e1�t B50A%1r  ��   ����8�\E�����	��|�:Y�#�3��B���  R�x*���D`T0 k� ������e1�t B50A%1r  ��   ����8�`CK����	��|�9Y�#�3��B���  R�|*���D`T0 k� ������e1�t B50A%1r  ��   ����8�dCKǿ��	��|�8Y�#�3��B���  R�)���D`T0 k� ������e1�t B50A%1r  ��   ����8�h~CKǾ^��	��|�8Y�#�3��B���  R�)���D`T0 k� ������e1�t B50A%1r  ��  ����8�p~CK˼^��L�|�7Y�#�3��B���  R�(���D`T0 k� ������e1�t B50A%1r  ��   ����8�t~CKϻ^��L�|�7Y�#�3��B���  R�(���D`T0 k� ������e1�t B50A%1r  ��   ����8�|~E�Ϻ^��L�|�6Y��3��B���  R�'���D`T0 k� ������e1�t B50A%1r  ��   ����8                                                                                                                                                                            � � �  �  �  c A�  �J����  �     � \��m| ]��s%C �  �  "Q           � ;k�    ��9m ;P    ���            ����            ��     ���   0			            D�  $ $      ��eO�     54�eO�     �                  ��        �     ���   (
             $           �O+     �4�iw    ��t              ����          ��     ���   8�

           ǟ   $ $     �(x     ǟ�(x                       		  �$          �     ���   (	            '�           .�A	)    ��*L�A	)    ��     	             ���$          ?�     ���   P
B            o. ��     B�y�    ��u��q�    �� r                 	  �p���K        �   Z  ���    8		 1               �� ��
	      V ��
    ��8 ��	    ����                     '����        �    K  ��@    		 5              �   	   j�u�B      E�u�B    U                    7         p     ��H   0            ��        ~  �    ���  �               ��        	 � !�        ��       ��F   @
%            �� $ $      ��MD�     ���MB"       %               	 D �        	       ��@   0            ��  � S	     � �f    ��� � �     f �               �� �         
 ��
`  �  ��P   0
	 

           � ]      � �u�    ��� �q\       C                    �          �     ��@   8'                 ��      �                                                                           �                               ��        ���          ��                                                                 �                           ��  ��        � N(;    ��� N    ��� "                x                j          �                               ��        � O      ��   N           "                                                �                                                          	               
 
       � �  +��       
�< U� 
� V  
� V  
�< V� 
� V� 
� W  
�< W� 
�| W� 
�\ W� 
� W  s�  n� J$ x� D� `^@ E�  _  E�  _@ �� j� � �j� �$ l  
�< W� 
�| W� 
�\ W� �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ 
�\ U� 
�� V  
�| V ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����b����      ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"     
�j,� B �
� �  �  
�       ��     � ;            ��     � ;            ��     ��u          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �       �� � �  ��        � � �  ���        �        ��        �        ��        �    ��     �l�����        ��                         ��q <  ������                                     �                 ����          
   �� ; ���%��  ���b ����           25BUF as Steen v      1:05                                                                        2  0     �"( �� �"� � �
 �"�*� �2X �2	P �2	
l �r �bS � �"4 �  " � � !� �   *9   *9 �*P �  )�` �"�P � "�b ��L �
�[* "I �B"( �B  "O �B "R �J  " � � "A � " |" "P �" "* |:!"< �B""2 |Z "6 | �$": � � %"P � �&!� �"'"* |:("< �B)"2 |Z*"6 |Z "
 �Z "
 �"-"* |:."< �B/"2 |Z0"6 |Z "
 �B2"2 |Z "6 |4"* |#5"< �+6"2 |C7"6 |K 8" �K  "D �S )�v ;*Ge <*Eu<="}T )�uE * |                                                                                                                                                                                                                         @ �   �     �               �     X P E Y  ��                     �������������������������������������� ���������	�
��������                                                                                          �� 
 ��~��� �������������������������������������������������������� ,�\, �  
��                                                                                                                                                                                                                                                                                                                                                                    ��                                                                                                                                                                                                                                                     �             L�J                                     �����������������������������������������������������                                                                                                                                                     )    ,,             ,          ,,                 	 	 ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ���               7                      C         ��  K
�J      %%  	                           ������ A���������������������������������������������                                                                                                                                                   "   � �         
      , 7      ,,              	 	 
  	 
 
 ���������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������                                                                                                                                                                                                                                                           
                                                                       �             


             �  }�    �    �#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" A C 6                                 � P}� �\                                                                                                                                                                                                                                                                             �   !�"E!�  
$                                `      a                                                                                                                                                                                                                                                                                                                                                                                                                                       j   5  : 3 ,7 7  ?Lpj  q� �����������������������������Z�����Z�����Z                       � {           �   & AG� �  �   
              �                                                                                                                                                                                                                                                                                                                                        I F   �                     !��                                                                                                                                                                                                                            Y��   �� ��        �� 3      ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ������������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&               ��                       4     �   ���������J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  p���� ��    ��Pp  ��     �f ��     �f �$ ^$ �@       �       �     �   h 
� � v           
  �   ��  
  �   �$ ^$ x x      ���  �         9    � �� g�      ��   f ^�       ��  p    �           ���� 
�*�����������     �  �          ��Φ��� 
�*���� 1| r� �  ��  yf  y<  ��������������������������������GvdDGw6wGwcfGwsfGwv6Gww6GwwcGwwcDDDDwwwwffffffffffffffffUUUUttttDDDDwwwwffffffffffffffffUUUUtttwN���t���wN��wt��wwN�wwt�wwwNwwwtGwweGwwU�tvf�wff�Fff�Fff��df��ffwwwwUUUUffffftDDft33gt5egt6Vgt5gwwwwUUUUffffDDDD3333eeeeVVVVwwwwwwwwUUUUffffDDFF35FfefDDVVFUufGfwwwwGwwwGwwwUUUUffffDDDDUUUUffffwwwwwwwuwwwuUUUUffffDDDDUUUUffffwwwwUUUUffffddDDfd33DD6VUd5eft6WwwwwUUUUffffDDGf35GfVVGvefGv6VGvwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwN�Fft�FfwN�dwt�fwwNGwwtGwwwDwwwtwt6Wwt5gwt6Wwt5gwt6Wwt5gtt6Wwt5gDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD6VGd5fGd6VGd5fGd6VGd5fGd6VGd5fGdFt5gFt6WFt5gFt6WFt5gFt6WFt5gFt6W5fGw6VGw5fGw6VGw5fGw6VGw5fGG6VGwgwwwvwwwwgwwwvwwwwgwwwvwwwwgwwwvGt6WGt5gDt6WDt5gND6WNt5gNt6WNt5g6VGd5fGf6VGw5fDD6VGU5fGf6VGf5fGfDDDDffffwwwwDDDDUUUUffffffffffffFt5gft6Wwt5gDD6WUt5gft6Wft5gft6W5fGt6VGt5fGD6VGD5fD�6VG�5fG�6VG�GwwwDwww�Gww�Dww~�Gww�Dww�DGw~�DNt6SNt5fNt6VNteeNwFVNwteNwwFfffd3333ffffVVVVeeeeVVVVeeeeffffDDDD333DffcDVVSDeecDVVSDeecDfVSDFecDUUUUDDDDDDDDDDDDDDDDDDDDDDDDDDDDD333D6ffD6VVD5fdD6VDD5fDD6VDD5fD3333ffffVVVVDDDD33335UUU5Vff5VDD3333ffffVVVVDDDD3333UUUUffffDDDD6VGfefGfVVGwDDDD3333UUUUffffDDDDffffffffwwwwDDDD3333UUUUffffDDDDft5cft6Vwt5eDDDD3333UUUUffffDDDD3333ffffeeeeDDDD3333UUUVffeVDD5V333DffcDeecDF6SDD5cDD6SDD5cDD6SDD333D6ffD5eeD6VVD5eeD6VVD5ffD6Vd5fG�fVG�efG�VVG�edw�VGw�dww�Ffffffffwwwwwwww����DDDDNNDD��������gwwwwwwwwwww��wwDDGwDDDw��DG���Dwwwwwwwwwwwww~��wwn�wwvwwwwgwwwvFfffFfffCeeeCVVVCeeeCVVVCeeeCVVVfDDDfDDDfDDDVDDDfDDDVDDDfDDDVDDDDfSDD5cDD6SDD5cDD6SDD5cDD6SDD5cDD6VDD5fDD6VDD5fDD6VDD5fDD6VDD5fD5VDD5VDD5VDD5VDD5VDD5VDD5VDD5VDDDDDDDDDADDDADDDDDDDDDDDADDDADDDDDDDDDDDDDDwDDDDDDDDDDDDDwDDDDD5VDD5VDD5VDD5VDD5VDD5VDD5VDD5VD5cDD6SDD5cDD6SDD5cDD6SDD5cDD6SDDDDfDDDfDDD5DDD6DDD5DDD6DDD5DDD6fffdfffdeeedVVVdeeedVVVdeeedVVVdCeeeCVVVCeeeCVVVCeeeCVVVCeeeCVVVfDDDVDDDfDDDVDDDfDDDVDDDfDDDVDDDD6SDD5c3D6VfD5eeD6VVDVffDDDDDDDDDDDD3333ffffeeeeVVVVffffDDDDDDDDD6VD35fDffVDeefDVVVDfffDDDDDDDDD5VDD5VDD5V335UUU5UUU5UUUVfffDDDDDDDDDDDD3333UUUUUUUUUUUUffffDDDDDD5VDD5V335VUUUVUUUVUUUVffffDDDDD5cDD6S3D5ffD6VVD5eeD6ffDDDDDDDDD5fD36VDfefDVVVDeefDfffDDDDDDDDDDDD5DDD6DDD5DDD6DDD5DDD6DDD5DDD6eeedVVVdeeedVVVdeeedVVVdeeedVVVdwwww�twwww~ww�w�wtwwtwwww~w�wwwwDDDDDDDDDADDDDDADDDDDDDDDDDtDD4DDqt4DDDD4DDsDDDDDDDDDDDD7AtCADADDADADDDDDDDADDDADDADqDADqDDDDDADDDADDDAADAADqADDAGADDDDwwwywww�www�www�www�www�www�www�������������������������www�www�www�www�www�www�www�www����������������������!�����!�-����������!-�����������!�����wwwwwwwtwwwOwww�wwt�ww�wwOGww�D��������������-��������������������������!����������-������NNNNNNNNNNNNN���FfwfDDDDDDDDDDDDNNNDNNNDNNND����gvftDDDDDDDDDDDDwts"wwB2ww22ws#Cws#4ww2twws�www�www�www�www�www�www�www�wwwywwww��������wwww������!��������wwwwww��w��w2��w���w��t���(�wy���������y���w�����y��Gwwwwt33Dt343CeeeCVVVEeeetVVVvEee�DVVzDFf�DDDfDDDVDDDe333VfffeeeeVVVVffffDDDDDDDDDDDD3333ffffeeeeVVVVffffDDDDDDD5DDD6333efffVeeeeVVVVffffDDDDeeedVVVdeeedVVVGeedgVVDzfdD�DDD�Df��NvDGN�DNN�DND~DGD��NDNt�DDDN#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFw"GC42wsDCwt�Cwt��ws�DGt�T7DfEGt{�Gwz��w���wt�Gw��wt�Gw�wtw�{�Gww��w��w2��w���w��w���x�wy����wwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wt3Gwt4wCGGttwG4�twO�wGt�GwE��wTfNw~D�����������������DD��ww�N��D�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wfuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGy�wwy�wtw�wOw�w�w�D�w2?�wCOGww�Dwwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGww23ws""wr22w244w#tD�t3~�}�ww}O3#�w""7w##'wCC#wDG2w3G~������wwwwVtwwUvwwenwwvWwwv�wwtwwtGww�3#�w""7w##'wCC#wDG2w3G~��7���wwww}�ww}�ww}�www�www}www}wwwwwwwr��ww��ww���w4��w��ww��www}ww'r'ww"GCw2wswCwtwCwtw�wswDGtwB'tww"w#w�2w�3w�3wG4wtGDwww"wr!r'wrwuUUG4wwD4wwCtwwCtww7tww7twwGtww8�3�3�3�8�3�3�33333"2#333"33UUUUwwwtwwwtwwwtwwwtwwwtwwwtwwwt��33�?33�?33�?333333#23323#3UUUUwwwwwwwwwwwwwfgvwwwwwwwwwwwwUUUUwwwtwwwtwwwtfwfdwwwtwwwtwwwtUUUUwwwwwwwwwwwwwwwwwwuwwwWwwwwwUUUUwwwWwwwWwwwWwwuwwwuwwUuwwwUwC�38C838C�38C833C332C"33C2#3UUUUwww~www~www~www~www~www~www~UUUUwfwnwvw~wfw~wvw~www~wfw~wgw~UUUUuwwwuwwwuwwwwWwwwWwwwWuwWUwwUUUUwwwwwwwwwwwwwwwwWwwwwwwwwwwwUUUUwwwdwwwdwwwdwwwdwwwdwwwdwwwdUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwUUUVwwwvwwwvwwwvwwwvwwwvwwwvwwwvGtwwGtwwGtwwGtwwGtwwGtwwGtwwGtwwwwwtwwwtwwwtwwwtwwwtwwwtwwwtwwwtww�www�www�www�www�www�www�www�w�www�www�www�www�www�www�www�wwwwwwdwwwdwwwdwwwdwwwdwwwdwwwdwwwdwwwvwwwvwwwvwwwvwwwvwwwvwwwvwwwvGtUUGTffGTffEdffEdffFdffFdffFdffUUUUfffffffffffffffffffffffff���UUUUffffffffffffffffffffffff����UU�Uff�eff�Vff�Vff�fff�fff�fʦ�f�UUU�fff�fff�fff�fff�fff�fff�fffUUUUffffffffffffffffffffffffffffwwwdwwwdd333d333d333d333d333dwwwwwwww33333333333333333333wwwvwwwv33363336333633363336FdffFdffAC333C333C333C333C333��������33333333333333333333�f�f�fFf�33�333�333�333�333�3�fff�fff33333333333333333333ffffffff33333333333333333333333d333d333d333d333d3333����wwww333333333333333333333333����wwww333633363336333633363333����wwwwC333C333C333C333C3333333����wwww33�333�333�333�333�33333����wwww�����<��5UUU5UUSU553SS2#33"532 5�����<��5UUU5UUUU555SSSS33333��������UUUUUUUU5555SSSS3333��������UUU�UU_�55=�SS]�33;������l���eUUUUUUSU552SS2#S3"3S2 0�����<��5UUU5UUSU552SS2#33"332 0����ȩ��S�UUU��US:�U59��38��009������<��UUUUUUUU5555SSSS33333������ÓUUX�UUS�SSX�553�338�003�����3���UUUU5UUUU555SSSS33333�����̚�Ue�5UX�U5Y�5X��S9��3����������UUUUUUUSU5523S2#"302 0�����<��5UUU5UUSU552SS2#33"302 0�����<��5UUV5UUUU555SSSU33353��������UUUUUUUUU5553SSS33330����l���eUUSUUU3SSS%U3"5S2#3S" "#  %                     200            "          "                         0;�  ��  �� ��  ۰  ۰  ��  ��                          #                         P"R                         "#                       "#  "                    0"                                                    �  9                     �#�� ��� ��� ��  �       02(�" �  � ��0(�������� �����   �                    "                         205            "         R 20R                                                                                    ��  ��  �� �� �  �  �  �   �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��  �S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG      w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  "!    " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  "!    " ""  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  "!  " ! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   ��  ��  ��  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    ��   �   ��� ������ �   �      �       �                        �   ��  ���  � �    �      �  �   �   �   �                                                                                                                 �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �                  ���� ���  ��    �            �   ������  ��             �  �                              �������  ���    �                    ��  ��  ���  ��  �  �  �   �                                                                                                                                                                                                    	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                                   ��                  �                        ���� ��� ����                             ����                                                                                                                                                                                                            �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �                   Ͱ  ˻  ˻  ۻ  ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                            �������  ���    �                    ��  ��  ���                                                                                                                                                                                                  	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                � ��                    ���� �                                                                                                                                                                                                        �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �           �   �     �   �                                          �   �           �   ̰  �˰                                                                                                                                                                                                         �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��                  �          �         �   �  �  �   �               �   �               � � ����� ��                                                                                                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                                  �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                �    � �  ��                  ���                                                                                                                                                                           ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r`                            ��  ����   �       �                                   �    ���  ��                    ��  ��  ���  ��  �  �  �   �                                                                                                                                                                                   �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   �  �  �  �   �   �       �  �,� �"/�""�"/� "/  �         "  "  ""  "+� �� � ��   �  "   "�  +�  
�� ��� D�D 4ETO3    �   �   �   D   E�  U�  UO                         "  "  "                                                                                                                                                                  	�  �� �� ���ܙܽɪ�͚�����͙ͼ̨��̄DC"�D32�C33�333�33P330X̽ 
�� ˪  "   ""/"""�����vv ��p ��  ��  ̽  ˸  ɚ  ��  ؛  -�� .ܰ .��  �"  �   .   "�                   � �  ��            Z   Z   Z   Z  Z  �� �� �� "� "" "" ""/ ����   �   � ���� �� ����                    �� ��������p��}`     �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                  �� �� �� }���ݪvw� w
�  ��  �� 
�� 	�� �� ��� ���+��Ҽ˝"���2+�    H   X   H   �   
          "�"    �                        ��� ��� ��ذ�̽м������ ��� ��̀��̘���D���T؊�T4�UDH�D@�TD �D8 �3: �� � + �" �"" �!"/��"/� ��� � �  �              �   ��  ��                              �       �                  "���"   "                                ���    �   "   "   "  !�� �  ��                                 � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                               �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""������������������""""���������������������""""������II������""""������IIII""""������DI�I�""""������DI�I�""""�����IIDIIIA""""��������DD""""������IADD�A��""""��������I���I�������I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD���4���4���4���4���4���43334DDDDDN��DDN��DDN��DDDDDNDDDNDDDDDNvSV~DGefS5v~D�EfSs�~D3�fUS~NC3g�U3V�C3~S35ns31Wc3Sqe5gDvS3Uw�DD��ww���w����N���������ffEUUUA3333S3333333333333333333333333333333333333333333DDDDVfwwN��DvffUwvffwwvf�wwvwwwwffffUUUU333333333333333333333333333333333333333333333333DDDD����DDDDS5UUS3fUSffUSwvfUfffeUUUU333333333333333333333333333333333333333333333333DDDDwwvfDDDDffeSUffe5ffUfSVU3S3333333333333333333333333333333333333333333333333DDDDfUU3DDNN1U  SUPeSUfeSgve1UffU3UUf5V31533133333333313331333333333333333333333333DDDD35UDD��        P   UP  5f  fn` ge� ~G>`g�s�V~G>5g�qV~G5g�V~5n13W163U3533DDNvgwDD�NDN      �� 
��        
������� ��  �� 
�������                        �������         �����
�� 	�   ���������                          �  	�� 
�� ��� ����� ��  
�  	�   �   �                                                    �   �   �                       DD~DDDD�DDDNfnDDEV�D5TdDUdD5dDUF�DenDDDDDDDDDFNDDrDDvP530   �Nwg���eN��e��Nv�N�vGN~NFd�tFd~�F6G�v6TDc%ef#%RR521520       w�DNV~��1fwfSUQfS�eUVN���tDDD����DDDDffff23S%S!" 2# 3 0   #����uf~NQgt�3n�DV~NDf�dN�GdDD~dN~�dNNcfDeVVD%5bt25gSU % 0 3                               ~  nDDDDD DD ��! %          �w D~ w~ D~�w~�~��D�DDDDDDDDDDDDDDDDDDDDDDDDDDD0S"     ~DN~�DN�DDNDDDNDDDDDDDDDDDDDDDDDDDDDDDDDDDDNDDD�DD�b#R23       DDN�DD�DDNDDD�DNDDD�DD�eNDDUDD�d�D��fdNNbdND&D�RtDSVt %"   DDG�DDDNDDDD�f�DeTnDCUVDQ5VDQFDTUnD�V�DDDDD�DDDD�DGDDGe3%  N��vN�Nv��NvNN��N��GDt��DfNgDfG�Dfd~GeeDF!VVe%%Ue"P3"S%3"Q    w~�DUg��Sgve1UUfe1�fUUD���gDDD����DDDDffff!2RR223% # 0   ��~��Vg�ewN6��5g��fnFD��vDDG�Dw�fDD�SdfRb4RU&cRV"3Q                               0  � dD �D �D  n�           w  �G  ww G� ww����~DDD�DDDDDDDDDDDDDDDDDDD�DDDR%       w�D��DD��DD�DDD�DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDNDDN�52RR        �DD�DDNDDD�DDNDDDDDNDDNFD�DEDDNFNdNNFfD��&D�b5dNR"gDPP5g  0   DDG�DDDNDDDD�f�DeEnDSUVDA5FDQVDUEnD�V�DDDDD�DDDD�DGDDGcRR2   N��vN�Nv��NvNN��N��GDt��DfNgDfG�Dfd~GeeDFRVVe5bRPR%       w~�DUg��Sgve1UUfe1�fUUD���gDDD����DDDDffff2QRU2! %0     ��~��Vg�ewN6��5g��fnFD��vDDG�Dw�fDD�VdfUed2VgR""#Q%"                             0     �  dD0�D  �D  n�            w  �G  ww G� ww����~DDD�DDDDDDDDDDDDDDDDDDD�DDD"       w�D��DD��DD�DDD�DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDNDDN�"%Q        �DD�DDNDDD�DDNDDDDDNDDNFD�DEDDNFNdNNFfD��VD�aedNRQgD0R%g RP   �DDNDDDDDDDDD�f�NeEnFSUVEA5FFQVNUEn��V��DDDN�DDDD�DgDDGSS00    ���wNDfDNgQDD�eDFN�DDdNDD�DDeDD%DG&UDFb0DuV GbU2fP5UR    ~@  vt` Vv� U� g~� ��@ DN` 00    5S  "5  20  R5           N�DD�DDDDDDDDNfnD�EV�e5TDUU�d5��UFNNenNDDDD�DDtDNDStDD%RS    �N�wD�FaDD�uDDNv�Dd�dDFDdDFndDF �DFQDDveDDfQDGUeDv%%vaP%    w�  WgF gn QU^ fw� ��D DD� "   P   RR1 0 %  5R         N�DD�DDDDDDDDNfnD�UF�d5UDUU�e4��EVNNenNDDDD�DDtDNDStDDSSU    �N�wD�FaDD�uDDNv�Dd�dDFDdDFndDFQ�DFVDDveDDfRDGUeDvRRvbRR     w�  WgF gn QU^ fw� ��D DD�     ! QQ  %P Q U% PP                     �� ~DD 䪤 �IG j�� �i��� M��K��kK���K�w�G��{Ggw�                        	�  ��  �� �  ~� � ��� ���wDD�DDD�~DD              ~� �D J� �� �� ֚ m�`K���F���K���K�w�G��{Ggw�                @   @   p   �		  	�� 	�~ ��� ��������wDD�DDD�~DD              �  ~D  �J  �  j�  �n ��@���F���K���K�w�G��{Ggw�            �   D   �   �   �   � D  �~  �z�ݙw�ݖ��wDD�DDD�~DD              �  ~D  �D  ��  n�  �n ��@���F���K���K�w�G��{Ggw�            �   D   �   I   �   � D  G~  I|�j�|�5���wDD�DDD�~DD    `   �   `  s�  G>` �uu �GVP�Ne`~��pg�FpV�Fpg�Fp~Dg`DD~ �D@                                                                                          0                               1                            "S%3"Q                         # 0    0                  "3Q                            UU  Q  SV  UU  ff DD ��   �fNvQVN�ceD�eUdNvfdN�DDD��DD�D~�NNvffD�UU�E5tEfUnEUfvff  D   D Nu1gfffg�DDn�~�d�fgfGcVDGe6NvR"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��                                 � � �� � � � � ����l(�(a(�����������������                	 
   ��� � � � � �����y(�(�����������������   ������� ������� �� ������������   � � � � � � � �����((�l(=����������������   ��	�
��������    ��������������������   ��� � � � � �����((�(( ����������������        ����     ! " # # $! % &  ��   ' (����� � � �����(-(5(Xx���������������� ) * + , - .  �Ӥ�  / 0 �  1 2�� 3 4  ��  / 5 6+*) � � � ��� � �����(�xww����������������     7 8 9 : : : : : ; < = = = = = = > ?::::: @ A B     � � � � ��� �����ww�(���������������� C CC 7 8 DD  E F G H         DD  E F G H A B CCC �� � � ��� �� ����(+((�����������������    7 8�� ���%��                 A B   �� � � ��� � ����(W(�m(`����������������   Q 7 8                       A B(Q   � � � � ��� ���	B�(a((M���������������� V W X 7 8                       A B(XWV � � � ��� � ���	C�(-(� 
(����������������� V W \ 7 8                       A B(\WV� ���� � � ��	E	D�(( (-(����������������� V W ] ^ _ ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` a b(]WV��� � � � � ��	F ��(X((6(5���������������� V W c d e f g h i j V W  k h i d e f l V W(j m(h(g(f(e(dcWV � � � � � � � ��	G ��l((�x���������������� V W n o p q ] r s t V Wn ] r u o p q v V W(t(s(r(](q(p(onWV���������H������yxww���������������� V W w f g h i d e f V W x i d e f k h y V W(f(e(d(i(h(g(f(QWV � ��O�N�M�L�K�J�I������w(+�(���������������� V W z { ] r u o p q V W | u o p q ] r u V W(q(p(o(u(r(](q }WV�A�A�V�U�T�S�R�Q���P(�((5(U(,���������������� V W ~  � � � � � � � � � � � � � � � ���(��(��(�(�((~WV�]�]�\�[�Z�Y�X���P(N(,(U((=((+���������������� � � � � � � �  �   �  � �� �� �  � �� � � � �� � � � � � � � ��� �A��(( ���������������� �     � � � � � � � � � � � �����������    � � � � � � � � ��� �A��(Xx���������������� � � � � � � � � � � � � � � � � ����������� � � � �� � � � � � � � ��� �=�:	9ww���������������� � � � � � � � � � � � � � � � � � �� � � � � � ��� � � � �� � � � � � � � ���'�>�; 
�(���������������� � � � ��� � � � � ��� � � �� � ���� � � � � ���� � � �� � � � � � ���	3?	<(+((����������������� � � � � � � � � � � � � � � � ��� � � � � � � � � � �� � � ��� � � � � � �����(W(�m(`���������������� � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �	
	
	
	
	@���(a((M���������������� � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � � �� � � � � � �����(-(� 
(����������������� � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �� � �� � � � �� ���(( (-(����������������� � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq"( �� �"� � �
 �"�*� �2X �2	P �2	
l �r �bS � �"4 �  " � � !� �   *9   *9 �*P �  )�` �"�P � "�b ��L �
�[* "I �B"( �B  "O �B "R �J  " � � "A � " |" "P �" "* |:!"< �B""2 |Z "6 | �$": � � %"P � �&!� �"'"* |:("< �B)"2 |Z*"6 |Z "
 �Z "
 �"-"* |:."< �B/"2 |Z0"6 |Z "
 �B2"2 |Z "6 |4"* |#5"< �+6"2 |C7"6 |K 8" �K  "D �S )�v ;*Ge <*Eu<="}T )�uE * |3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������@�9�1� ���������������������������������������,�>�0�	�
�������������������� � � � � � �����������������������������������������%�� ������������������,�>�0� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K������������������������1�G�S�K��<�Z�G�Z�Y�����������������������9�R�G�_�K�X��<�Z�G�Z�Y��������������������<�I�U�X�O�T�M��<�[�S�S�G�X�_�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������/�+��2�U�I�Q�K�_��8�O�M�N�Z�������������������-�G�R�M�G�X�_� � � � � � � � � � � � � � �� � ����������+�T�G�N�K�O�S� � � � � � � � � � � � � � ��� ������������������������������������ 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                       	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 