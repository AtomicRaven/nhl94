GST@�                                                           �o�                                                          U   �     
         ��  2�������J��������     ����        ��      #    ����                                d8<n    �  ?     2����  �
fD�
�L���"����D"� j   " B   J  jF�"    B�j B����
��
�"    B�jl �   B ��
   �                                                                              ����������������������������������      ��    oo b go  4  +c  c  'c      ��       	  
    	G 7� V( 	(                 �n 1         8:8�����������������������������������������������������������������������������������������������������������������������������=  0b  4  11                                         �  �  �  �                  �  
)          = �����������������������������������������������������������������������������                                $�  �   r  K�   @  #   �   �                                                                                'w w  �1n  
)�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    @c B����$R\V�|( C<@,p#�N����4Z� T0 k� ��2��2�1	�"qe1�t B  ��*    � * @c A����%R\V�|( s<@,p#�O����4Z� T0 k� ��1��1�1	�"qe1�t B  ��*    � * @c A����&R\V�|( s<@,p#�P����3Z�  T0 k� ��1��1�1	�"qe1�t B  ��*    � * @c @����&R\V�|( s<B�,p#�Q����3Z�T0 k� ��0��0�1	�"qe1�t B  ��*    � * @c ?����'R\V�|( s<B�0p#�R����2Z�T0 k� ��0��0�1	�"qe1�t B  ��*    � * @c ?����'R\V�|( s<B�0p��S��� 2Z�T0 k� ��/� /�1	�"qe1�t B  �*    � * @c >����(R\V�|( s<B�4p��T���3Z�T0 k� ��0� 0�1	�"qe1�t B  ��*    � * @c =��#�(RXV�|( �<B�4p��T���3Z�T0 k� � 1�1�1	�"qe1�t B  ��*    � * @c$=��#�(RXU�|( �<B�8p��U���3Z�T0 k� �1�1�1	�"qe1�t B  ��*    � * @c$<��#�)RXU�|( �<B�8p��V���3Z�T0 k� �1�1�1	�"qe1�t B  ��*    � * @c$;��#�)RXU�|( �<B�<p��WC��3Z�T0 k� �1�1�1	�"qe1�t B  ��*    � * @c$;��#�*RXU�|( �<B�@p��XC��3Z�T0 k� �1�1�1	�"qe1�t B  ��*    � * @c$:��#�*RXU�|( �<B�Dp��XC��3Z� T0 k� �1�1�1	�"qe1�t B  ��*    � * @c$:��#�*RXU�|( �<B�Hp��YC��4Z�$T0 k� �1�1�1	�"qe1�t B  ��*    � * @c$9��#�+RXU�|( �<B�Lp��ZC� �4Z�$T0 k� �2�2�1	�"qe1�t B  ��*    � * @c$9��#�+RXU�|( �<B�Pp��[#�!� 4Z�(T0 k� �2�2�1	�"qe1�t B  ��*   � * @c$8��#�,RXU�|( s<E�Tp��[#�"� 4Z�(T0 k� �2� 2�1	�"qe1�t B  ��*    � * @c$7��#�,RXU�|( s<E�Xp��\#�#�$4Z�,T0 k� � 2�$2�1	�"qe1�t B  ��*    � * @c$7��#�,RXU�|( s<E�\p��]#�%�(4Z�,T0 k� �$2�(2�1	�"qe1�t B  ��*    � * @c$6��#�-RXU�|( s<E�`p��^#�&�(4Z�0T0 k� �$2�(2�1	�"qe1�t B  ��*    � * @c$6��#�-RXU�|( s<E�dp��^#�'�,4Z�0 T0 k� �(2�,2�1	�"qe1�t B  ��*    � * @c$5��#�-RXU�|( s<E�hp��_#�(�05Z�4 T0 k� �,3�03�1	�"qe1�t B  ��*    � * @c$5��#�.RTU�|( s<E�pp��`�)�05Z�4 T0 k� �,3�03�1	�"qe1�t B  ��*    � * @c$4��#�.RTU�|( s<E�to��`�+�45Z�8 T0 k� �03�43�1	�"qe1�t B  ��*    � * @c(4��#�.RTU�|( s<E�xo��a�,�85Z�8!T0 k� �43�83�1	�"qe1�t B  ��*    � * @c(3��#�/RTU�|( C<E�|o��b�-�85Z�8!T0 k� �43�83�1	�"qe1�t B  ��*    � * @c(3��#�/RTU�|( C<B�n��b�/�<5Z�<!T0 k� �83�<3�1	�"qe1�t B  ��*    � * @c(2��#�/RTU�|( C<B�n��c�0�<5_�<!T0 k� �<3�@3�1	�"qe1�t B  ��*   � * @c(2��#�0RTU�|( C<B�n��d�1�@5_�<"T0 k� �<3�@3�1	�"qe1�t B  ��*    � * @c(2��#�0RTU�|( C<B�m��d�3�D6_�<"T0 k� �@3�D3�1	�"qe1�t B  ��*    � * @c(1��#�0RTU�|(  <B�l��e�4�D6_�<"T0 k� �H4�L4�1	�"qe1�t B  ��*    � * @c(1��$ 1RTU�|(  <B�l��e��6�H6_�<"T0 k� �P4�T4�1	�"qe1�t B  ��*    � * @c(0��$ 1RTU�|(  <B�k��f��7�L6_4<"T0 k� �X4�\4�1	�"qe1�t B  ��*    � * @c(0��$1RTU�|(  <B�k��g��8�L6_4<"T0 k� �\4�`4�1	�"qe1�t B  ��*    � * @c(/��$2RTU�|(  <C�j��g��:�P6_4<"T0 k� �`4�d4�1	�"qe1�t B  ��*    � * @c(/��2RTU�|( �<C�i��h��;�T6_4<"T0 k� �h8�l8�1	�"qe1�t B  ��*    � * @c(/�� 2RTU�|( �<C�i� h��<�X6_4<"T0 k� �p;�t;�1	�"qe1�t B  ��*    � * @c(.�� 3RTU�|( �@C�i�i��=�\7_48!T0 k� �t>�x>�1	�"qe1�t B  ��*    � * @c(.�� 3RTU�|( �@C�h�i��?�t7Z8"T0 k� �x>�|>�1	�"qe1�t B  �/    � * @c(-�� 3�3RTU�|( �@I3�h�j��@��7Z8"T0 k� �|>��>�1	�"qe1�t B  ��/    � * @c(-�� 3�3RTU�|( �@I3�g�j��A.$�7Z4"T0 k� �|>��>�1	�"qe1�t B  ��/    � * @c(-�� 3�3RPU�|( �DI3�g�k��B.$�7Z4"T0 k� �>��>�1	�"qe1�t B  ��/    � * @c(,�� 3�2RPU�|( �DI3�f�k��C.$�7Z4"T0 k� �?��?�1	�"qe1�t B  ��/    � * @c(,�� 3� 2RPU�|( �HI3�f�l��E.$�7Z4"T0 k� �?��?�1	�"qe1�t B  ��/    � * @c,,���3�$3RPU�|( �HIC�f�l��F.$�7Z4"T0 k� �?��?�1	�"qe1�t B  ��/    � * @c,+���3�$3RPU�|( LIC�f� m��G.$�7Z4!T0 k� ��?��?�1	�"qe1�t B  ��/    � * @c,+���3�(3RPU�|( LIC�e�$m��H.4�7Z4"T0 k� ��@��@�1	�"qe1�t B  ��/    � * @c,+���3�(3RPU�|( PIC�e�$n��I.4�7Z4"T0 k� ��@��@�1	�"qe1�t B  ��/    � * @c,*���3�,3RPU�|( TIC�e�(n��J.4�7Z4"T0 k� ��@��@�1	�"qe1�t B  ��/    � * @c,*���3�,3RPU�|( TI3�e�,o��K.4�7Z0"T0 k� ��@��@�1	�"qe1�t B  ��/    � * @c,*���3�03RPU�|( XI3�e�0o��L.4�7Z0"T0 k� ��A��A�1	�"qe1�t B  ��/    � * @c,)���3�03RPU�|( \I3�e�4o��M.4�7Z0"T0 k� ��A��A�1	�"qe1�t B  ��/    � * @c,)���3�44RPU�|( \I3�e�4p��N.4�7Z0"T0 k� �A��A�1	�"qe1�t B  ��/    � * @c,)���3�44RPU�|( `I3�e�8p��O.D�7Z0"T0 k� �A��A�1	�"qe1�t B  ��/    � * @c,(���3�84RPU�|( dIC�e�<q��P.D�7Z0"T0 k� �A��A�1	�"qe1�t B  ��/    � * @c,(���3�84RPU�|( hIC�e�<q��Q.D�7Z0"T0 k� �B��B�1	�"qe1�t B  ��/    � * @c,(���3�<4RPU�|( lIC�e�@q��R.D�7Z,#T0 k� �B��B�1	�"qe1�t B  ��/    � * @c,'���3�84RPU�|( pIC�e�@q��S.D�7Z,#T0 k� �B��B�1	�"qe1�t B  ��/    � * @c,'���3�85RPU�|( tIC�e�@q��T.D�7Z,#T0 k� �B��B�1	�"qe1�t B  ��/    � * @c,'���3�85RPU�|( xI3�e�@p��U.D�7Z,#T0 k� �C��C�1	�"qe1�t B  ��/    � * @c,'���3�85RPU�|( |I3�e�@p��U.T�7Z,$T0 k� �C��C�1	�"qe1�t B  ��/    � * @c,&���3�85RPU�|( �I3�e�@p��U.T�7Z,$T0 k� �C��C�1	�"qe1�t B  ��/    � * @c,&���3�45RPU�|( �I3�e�@o��U.T�7Z,$T0 k� �C��C�1	�"qe1�t B  ��/    � * @c,&���3�45RPU�|( � I3�f�@o��U.T�7Z($T0 k� �C��C�1	�"qe1�t B  ��/    � * @c,&���3�46RPU�|( ��!@c�f�@o��U.T�7Z($T0 k� �D��D�1	�"qe1�t B  ��/    � * @c,%��� d46RPU�|( ��"@c�f�Dn��V.T�7Z(%T0 k� �D��D�1	�"qe1�t B  ��/    � * @c,%��� d06RPU�|( ��#@c�f$Dn��V.T�7Z(%T0 k� �tD�xD�1	�"qe1�t B  ��"    � * @c,%��� d06RPU�|( ��%@c�f$Dn��V.T�7Z(%T0 k� �hD�lD�1	�"qe1�t B  ��"    � * @c,%��� d07RPU�|( ��&@c�g$Dm��V.T�7Z(%T0 k� �`E�dE�1	�"qe1�t B  ��"    � * @c,$��� d07RPU�|( ��'@c�g$Dm��V.T�7Z(&T0 k� �\E�`E�1	�"qe1�t B  ��"    � * @c,$����07RPU�|( ��(@c�g$Dm��W.T�7Z(&T0 k� �XE�\E�1	�"qe1�t B  ��"    � * @c,$����08RPU�|( ��*@c�g Dl��W.T�7Z(&T0 k� �TF�XF�1	�"qe1�t B  ��"    � * @c0$����48RPU�|( ��+B��g Dl��W.T�7Z$&T0 k� �XF�\F�1	�"qe1�t B  ��"    � * @c0#����49RLU�|( ��,B��g Dk� W.T�7Z$&T0 k� �XG�\G�1	�"qe1�t B  ��"    � * @c0#����49RLU�|( ��.B��g Dj� X.T�7Z$'T0 k� �XG�\G�1	�"qe1�t B  ��"   � * @c0#����4:RLU�|( ��/B��g Dj�X.T�7Z$'T0 k� �LJ�PJ�1	�"qe1�t B  ��"    � * @c0#����4:RLU�|( ��1B��fDi�X.T�7Z$'T0 k� �@L�DL�1	�"qe1�t B  ��"    � * @c0#����4;RLU�|( ��2K��fHi�X.T�7Z$'T0 k� �8M�<M�1	�"qe1�t B  ��"    � * @c0"����4<RLU�|( C�4K��fHh�X.T�7Z$'T0 k� �4O�8O�1	�"qe1�t B  ��"    � * @c0"����4=RLU�|( C�6K��fHh�X.T�7Z$(T0 k� �0P�4P�1	�"qe1�t B  ��"    � * @c0"��� �4=RLU�|( C�7K��fHg�X.T�7Z$(T0 k� �,Q�0Q�1	�"qe1�t B  ��"    � * @c0"��� �8>RLU�|( C�9K��f�Hf�X.T�7Z$(T0 k� �,R�0R�1	�"qe1�t B  ��"    � * @c0"��� �8?RLU�|( C�;K��f�Le�Y.T�7Z (T0 k� �,S�0S�1	�"qe1�t B  ��"    � * @c0!��� �8@RLU�|( C�=K��f�Le�Y.T�7Z (T0 k� �,T�0T�1	�"qe1�t B  ��"    � * @c0!��� �8ARLU�|( C�>K��f�Ld�Y.T�7Z (T0 k� �,U�0U�1	�"qe1�t B  ��"    � * @c0!��� �8BRLU�|( C�@K��f�Pc�Y.T�7Z )T0 k� �,V�0V�1	�"qe1�t B  ��"    � * @c0!��� �8CRLU�|( S�BK��ftPb�Y.T�7Z )T0 k� �,W�0W�1	�"qe1�t B  ��"    � * @c0!��� �8ERLU�|( S�BK��ftPa�Y.T�7Z )T0 k� �,X�0X�1	�"qe1�t B  �"    � * @c0 ���<FRLU�|( S�DK��ftP`�Y.T�7Z )T0 k� �,X�0X�1	�"qe1�t B  ��/    � * @c0 ���<GRLU�|( S�FK��ftT_�Y.T�7Z )T0 k� �0W�4W�1	�"qe1�t B ��/    � * @c0 ���@HRLU�|( T HK��ftT^�X.T�7Z )T0 k� �0W�4W�1	�"qe1�t B ��/    � * @c0 ���@IRLU�|( � HK��ftX]�Y.T�7Z *T0 k� �0W�4W�1	�"qe1�t B ��/    � * @c0 ���DKRLU�|( � IK��fdX\�Z.T�7Z *T0 k� �4W�8W�1	�"qe1�t B ��/    � * @c0 ���DDLRLU�|( � JK��fd\[�[.T�7Z *T0 k� �4V�8V�1	�"qe1�t B ��/    � * @c0���DDLRLU�|( � JK��fd\[�\.T�7Z*T0 k� �4V�8V�1	�"qe1�t B ��/    � * @c0���DDLRLU�|( � KK��fd`[�\.T�7Z*T0 k� �8V�<V�1	�"qe1�t B ��/    � * @c0���DDLRLU�|( � LK��fdd[� ].T�7Z*T0 k� �8V�<V�1	�"qe1�t B ��/    � * @c0���DDLRLU�|( � MK��fdd[� ^.T�7Z+T0 k� �8U�<U�1	�"qe1�t B ��/    � * @c0���DDLRLU�|( � NK��fdh[�$_.T�7Z+T0 k� �<U�@U�1	�"qe1�t B ��/    � * @c0���4DLRLU�|( � OK��f.�h[�$`.TX7Z+T0 k� �<U�@U�1	�"qe1�t B �/    � * @c0���4DMRLU�|( � PK��f.�h[�(a.TX7Z+T0 k� �<U�@U�1	�"qe1�t B ��/    � * @c0���4@NRLU�|( 	t RK��f.�h[�(a.TX7Z+T0 k� �@T�DT�1	�"qe1�t B ��/    � * @c0���4@NRLU�|( 	t SK��f.�h[�,b.TX7Z+T0 k� �@T�DT�1	�"qe1�t B ��/    � * @c0���4@NRLU�|( 	s�TK��f.�h[�,b.TX7Z+T0 k� @T�DT�1	�"qe1�t B ��/    � * @c0���4@NRLU�|( 	s�UK��f.�h[,c.TX7Z+T0 k� DT�HT�1	�"qe1�t B ��/    � * @c0���4<ORLU�|( 	s�VK��f.�h[,d.TX7Z,T0 k� DS�HS�1	�"qe1�t B ��/    � * @c0���48ORLU�|( 	��VK��g.�h[0d.TX7Z,T0 k� DS�HS�1	�"qe1�t B ��/    � * @c0���48ORLU�|( 	��VK��g.�h[0d.TX7Z,T0 k� HS�LS�1	�"qe1�t B ��/    � * @c0���48ORLU�|( 	��WK��h.�h[0e.TX7Z,T0 k� HS�LS�1	�"qe1�t B ��/    � * @c0���48PRLU�|( 	��WK��h.�h[0e.TX7Z,T0 k� HR�LR�1	�"qe1�t B ��/    � * @c4���48PRLU�|( ��XK��i.�h[0f.TX7Z,T0 k� LR�PR�1	�"qe1�t B ��/    � * @c4���48QRLU�|( ��YK��i.�h[0f.TX7Z,T0 k� LR�PR�1	�"qe1�t B ��/    � * @c4���44QRLU�|( ��YK��j.�h[0f.TX7Z-T0 k� �PQ�TQ�1	�"qe1�t B ��/    � * @c4���44QRLU�|( ��ZK��j.�X[0f.TX7Z-T0 k� �PQ�TQ�1	�"qe1�t B ��/    � * @c4���40QRLU�|( ��ZK��k.�X[0g.TX7Z-T0 k� �PQ�TQ�1	�"qe1�t B $�/    � * @c4���40QRLU�|( ��[K��k.�X[0g.TX7Z-T0 k� �TQ�XQ�1	�"qe1�t B ��/    � * @c4���40RRLU�|( ��[K��k.�X[0g.TX7Z-T0 k� �TQ�XQ�1	�"qe1�t B ��/    � * @c4���4,RRLU�|( ��[K��l.�X[0g.TX7Z-T0 k� �XQ�\Q�1	�"qe1�t B ��/    � * @c4���4,RRLU�!�( �[K��l.�X[0g.TX7Z-T0 k� �\Q�`Q�1	�"qe1�t B ��/    � * @c4���4(RRLU�!�( �[K��m.�X[ �0g.TX7Z-T0 k� �\Q�`Q�1	�"qe1�t B ��/    � * @c4���4(SRLU�!�( �\K��m.�X[ �0gDX7Z-T0 k� �`Q�dQ�1	�"qe1�t B ��/    � * @c4���4$SRLU�!�( �\K��m.�X[ �0gDX7Z.T0 k� �`Q�dQ�1	�"qe1�t B ��/    � * @c4���4$SRLU�!�( �\K��n.�X[ �0gDX7Z.T0 k� �dQ�hQ�1	�"qe1�t B ��/   � * @c4���4$SRLU�!�( �]K��n.�X[ �0gDX7Z.T0 k� �hQ�lQ�1	�"qe1�t B ��/    � * @c4���4$SRLU�!�( �]K��o.�X[0gDX7Z.T0 k� �hQ�lQ�1	�"qe1�t B ��/    � * @c4����$TRLU�!�( �^K��o.�X[0gDX7Z.T0 k� �lQ�pQ�1	�"qe1�t B ��/    � * @c4���� TRLU�!�( �^K��o.�X[0gDX7Z.T0 k� �lQ�pQ�1	�"qe1�t B ��/    � * @c4���� TRLU�!�( ��^K��p.�X[0gDX7Z.T0 k� pQ�tQ�1	�"qe1�t B ��/    � * @c4���� URLU�!�( ��_K��p.�X[0gDX7Z.T0 k� pQ�tQ�1	�"qe1�t B ��/    � * @c4����URLU�|( ��_K��p.�X[T0gX7Z.T0 k� tQ�xQ�1	�"qe1�t B ��/    � * @c4����VRLU�|( ��_K��q.�X[T0gX7Z.T0 k� xQ�|Q�1	�"qe1�t B ��/    � * @c4����VRLU�|( ��`K��q.�X[T0gX7Z/T0 k� xQ�|Q�1	�"qe1�t B �/    � * @c4����WRLU�|( ��`K��q.�X[T0gX7Z/T0 k� |Q��Q�1	�"qe1�t B ��/    � * @c4����XRLU�|( ��aK��r.�X[T0gX7Z/T0 k� |Q��Q�1	�"qe1�t B  ��/    � * @c4����YRLU�|( ��bB��r.�X[�0gX7Z/T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���DYRLU�|( ��bB��r.�X[�0gX7Z/T0 k� �Q��Q�1	�"qe1�t B  -�/    � * @c4���DZRLU�|( ��cB��r.�X[�0gX7Z/T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���D[RLU�|( ��cB��s.�X[�0gX7Z/T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���D \RLU�|( ӼdB��s.�X[�0g dX7Z/T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���C�\RLU�|( �dK��s.�X[�0g dX7Z/T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���C�]RLU�!�( �eK��s.�X[�0g dX7Z/T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���C�^RLU�!�( �eK��s.�X[�0g dX7Z/T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���C�_RLU�!�( �fK��s.�X[�0g dX7Z/T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���C�_RLU�!�( �fK��t.�X[�0g dX7Z/T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���C�`RLU�!�( �gK��t.�X[40g dX7Z0T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���C�aRLU�!�( �gK��t.�X[40g dX7Z0T0 k� �Q��Q�1	�"qe1�t B  ��/    � * @c4���C�aRLU�!�( �hK��t.�X[40g dX7Z0T0 k� �P��P�1	�"qe1�t B  ��/    � * @c4���C�bRLU�!�( �gK��t.�X[40g dX7Z0T0 k� �P��P�1	�"qe1�t B  ��/    � * @c4���C�cRLU�!�( �gK��t.�X[4,g dX7Z0T0 k� �P��P�1	�"qe1�t B  ��/    � * @c4���C�cRLU�!�( �gK��t.�X[4,g dX7Z0T0 k� �P��P�1	�"qe1�t B  ��/    � * @c4���C�dRLU�!�( �gK��u.�X[4,g dX7Z0T0 k� �P��P�1	�"qe1�t B  ��/   � * @c4���C�dRLU�|( �fK��u.�X[4,f dX7Z0T0 k� �P��P�1	�"qe1�t B  ��/    � * @c4���C�eRLU�|( �fK��u.�X[4(f dX7Z0T0 k� �P��P�1	�"qe1�t B  ��/    � * @c4���C�eRLU�|( �fK��u.�X[4(f dX7Z0T0 k� �P��P�1	�"qe1�t B  ��/    � * @c4���C�eRLU�|( �fK��u.�X[4$e dX7Z0T0 k� �O��O�1	�"qe1�t B  ��/    � * @c4���C�fRLU�|( �|eK��v.�X[4$e dX7Z0T0 k� �O��O�1	�"qe1�t B  ��/    � * @c4���C�fRLU�|( �xeK��v.�X[D$d dX7Z0T0 k� �O��O�1	�"qe1�t B  ��/    � * @c4���C�fRLU�|( �teK��v.�X[D d dX7Z0T0 k� �M��M�1	�"qe1�t B  ��*   � * @c4����gRLU�|( �peK��v.�X[D d dX7Z0T0 k� �K��K�1	�"qe1�t B  ��*    � * @c4����gRLU�|( �pdK��w.�X[D c dX7Z1T0 k� �|J��J�1	�"qe1�t B  ��*    � * @c4����hRLU�|( �ldK��w.�X[Dc dX7Z1T0 k� �xI�|I�1	�"qe1�t B  ��*    � * @c4����hRLU�|( �hdK��w.�X[Dc dX7Z1T0 k� �xH�|H�1	�"qe1�t B  ��*    � * @c4����iRLU�|( �ddK��w.�X[Dc dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*   � * @c4����iRLU�|( �ddK��w.�X[Dc dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����iRLU�|( �`cK��x.�X[Dc dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����jRLU�|( �\cK��x.�X[Dc dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����jRLU�|( �XcK��x.�X[Dc dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����jRLU�|( �XcK��x.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����kRLU�|( �TcK��x.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����kRLU�|( �PcK��y.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����lRLU�|( �PbK��y.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����lRLU�|( �LbK��y.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����lRLU�|( �HbK��y.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����mRLU�|( �HbK��y.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����mRLU�|( �DbK��z.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����mRLU�|( �@bK��z.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����nRLU�|( �@aK��z.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����nRLU�|( �<aK��z.�X[�c dX7Z1T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����nRLU�|( �<aK��z.�X[�c dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����oRLU�|( �8aK��z.�X[�c dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����oRLU�|( �8aK��{.�X[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����oRLU�|( �4aK��{DX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����oRLU�|( �0aK��{DX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����pRLU�|( �0`K��{DX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����pRLU�|( �,`K��{DX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����pRLU�|( �,`K��{DX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����qRLU�|( �(`K��|DX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����qRLU�|( �(`K��|DX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����qRLU�|( �$`K��|DX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4����qRLU�|( �$`K��|DX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4���|rRLU�|( � _K��|TX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4���|rRLU�|( � _K��|TX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4���|rRLU�|( �_K��|TX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4���xrRLU�|( �_K��}TX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4���xsRLU�|( �_K��|TX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4���tsRLU�|( �_K��|TX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4���tsRLU�|( �_K��|TX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4���tsRLU�|( �_K��|TX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4���ptRLU�|( �_B��{TX[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * @c4���ptRLU�|( �^B��{�T[Dc dX7Z2T0 k� �xG�|G�1	�"qe1�t B  ��*    � * C�Hs���_p� �s������C��	_��ˍ��Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8C�@s��_h���k������C�|	_��Í��Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8C�8s��_`���c������C�t	_������Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8C�0s��_X��=[������C�l	_������Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8C�$s�ۚ_P��=S������C�`	_������Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8C�s�Ӛ_L��=G������C�X	_������Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8C�s�ǚ_D��=?�����C�P	_������Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8C�sￚ_<��=7����w�C�H	_������Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8C�s﷚_4���/���o�C�@	_������Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8C��sﯚ�,
���'���c�C�4	_������Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8C��s����$	������[�C�,	_������Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�s����������S�D $	_������Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�s����������K�D 	_�����Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�s����������C�D 	_��w���Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�s������ �����;�D 	_��o����Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�s�{�����!�����/�D  	_��k����Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�s�s�����"�����'�D�	_��c����Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�s�k�����$������D�_��[����Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�s�c���˜%������D�_��S����Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�s�[��� ˘&������D�_��K����Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�s�O����ː(������D�	_��C����Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�sG����ˌ)�������D�	_��;����Z3�T0 k� �k��o��1	�"qe1�t B  ��?    ����8D�r?����ˈ*�������D�	_��3���Z3�T0 k� �h�l�1	�"qe1�t B  ��?    ����8D|r7����ˀ,�������D�	_��+���Z3�T0 k� �h�l�1	�"qe1�t B  ��?    ����8Dtr/�����|-�������D�	_��#���Z3�T0 k� �h�l�1	�"qe1�t B  ��?    ����8Dlr'�����x.�������D�	_�����Z3�T0 k� �h�l�1	�"qe1�t B  ��?    ����8Ddr�^���p0�������D�
_�����Z3�T0 k� �h�l�1	�"qe1�t B  ��?    ����8DXr�^���t1�������D�
_�����Z3�T0 k� �h	�l	�1	�"qe1�t B  ��?    ����8DPr�^���t3�������D�
_�����Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8DHr�^���t4������D�
_|�����Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8D@r��^���x5��|���D�
_x����Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8D,r�^s��x8{�|���D�
_p����Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8C�$rߚNk��|9w�|���C�
_l�׎��Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8C�rךNc��|;o�|���C�
_h �ώ��Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8C�rϚN[��|<k�����C�_d �ǎ��Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8C�rǚNO��|=c���쏿C�_d ���Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8C� r��NG�ۀ>_���쇾C�_c����Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8C��r��N?�ۀ@W�����C�__��A��Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8C��r��N7��AS�����C�_[��A�Z3�T0 k� �h�l�1	�"qe1�t B  ��? 
   ����8C��r��N/��BO����w�C�_W�A��A{�Z3�T0 k� �h!�l!�1	�"qe1�t B  ��3 
   ����8C��r��N��DC����w�C�|_O�A��Ao�Z3�T0 k� �h%�l%�1	�"qe1�t B  �3 
   ����8A]�r^����E?���\o�A_t_K�A��Ag�Z3�T0 k� �h(�l(�1	�"qe1�t B  ��3 
   ����8A]�r^����|F7�� \k�A_l_K�A{�Ac�Z3�T0 k� �d*�h*�1	�"qe1�t B  ��3 
   ����8A]�r^{���|G3��\c�A_h_G�As�A[�Z3�T0 k� �d,�h,�1	�"qe1�t B  ��3 	   ����8A]�r^s����|H/��\[�A_`_C�Ao�AS�Z3�T0 k� �d.�h.�1	�"qe1�t B  ��3 	   ����8A]�r^k����|H'�� \W�A_\_?�g�O�Z3�T0 k� �d/�h/�1	�"qe1�t B  ��3 	   ����8A]�r^c����|I#�� \O�A_T_?�_�K�Z3�T0 k� �\2�`2�1	�"qe1�t B  ��3 	   ����8A]�r^[����|JL�� \K�A_P_;�W�C�Z3�T0 k� �X5�\5�1	�"qe1�t B  ��3 	   ����8A]�r^S����|JL�� \C�A_H_7�O�?�Z3�T0 k� �T7�X7�1	�"qe1�t B  ��3 	   ����8A]�r^K����|KL�� \?�A_D_3�G�7�Z3�T0 k� �T8�X8�1	�"qe1�t B  ��3 	   ����8A]�r^G�����KL�� \7�A_<_3�?�0 Z3�T0 k� �T:�X:�1	�"qe1�t B  ��3 	   ����8A]|r^?�����LL�� 	\3�A_8_/�;�, Z3�T0 k� �T;�X;�1	�"qe1�t B  ��3 	   � �8A]tr^7�����LL�� 
\+�A_0_+�3�$ Z3�T0 k� �T<�X<�1	�"qe1�t B  ��3 	   � �8A]lr^/�����ML�� \'�A_,_'�+�  Z3�T0 k� �T=�X=�1	�"qe1�t B  ��3 	   � �8A]hr^+�����MK��� \�A_(_'�#�Z3�T0 k� �T=�X=�1	�"qe1�t B  ��3 	   � �8A]`r^#�����MK��� \�A_ _#��Z3�T0 k� �T=�X=�1	�"qe1�t B  ��3 	   � �8A]Xr^�����MK��� \�A__��Z3�T0 k� �X>�\>�1	�"qe1�t B  ��3 	   � 	�8A]Pq^�����NK�� \�A__��Z3�T0 k� �X>�\>�1	�"qe1�t B  ��3 	   � 
�8A]Lq^���ˈNK�� \�A__��Z3�T0 k� �X>�\>�1	�"qe1�t B  ��3 	   � �8A]Dq^���ˈNK��$\�A__��Z3�T0 k� �X>�\>�1	�"qe1�t B  ��3 	   � �8A]@q^���ˈNK��$[��A__� �� Z3�T0 k� �X>�\>�1	�"qe1�t B  ��3 	   � �8A]8q]���ˈNK߻�$[��A__� �� �Z3�T0 k� �X>�\>�1	�"qe1�t B  ��3 	   � �8A]0q]��{�ˈNKۺ�$[��A_ _� � �Z3�T0 k� �X?�\?�1	�"qe1�t B  ��3 	   � �8A],q]�s�[�NK׺�$[�A^�_� � �Z3�T0 k� �TC�XC�1	�"qe1�t B  ��3 	   � �8A]$q]�o�[�NK׹�$[�A^�_� � �Z3�T0 k� �PF�TF�1	�"qe1�t B  ��3 	   � �8A] q]�g�[�NKӹ�$[�A^�_� � �Z3�T0 k� �PH�TH�1	�"qe1�t B  ��3 	   � �8A]q]ߚc�[�OKϸ�$[�A^�_� ە �Z3�T0 k� �LJ�PJ�1	�"qe1�t B  ��3 	   � �8A]q]ۚ_�[�OK˸�$[ߧA^�_� ו �Z3�T0 k� �LK�PK�1	�"qe1�t B  ��3 	   � �8A]q]ӚW�[�OKǷ�$[ۦA^�_� ӕ �Z3�T0 k� �LL�PL�1	�"qe1�t B  ��3    � �8A]q]ϚS�[�OK÷�$[ӥA^�_� ˕ �Z3�T0 k� �PM�TM�1	�"qe1�t B  ��3    � �8A]q]˚K�[�OK���$[ϥA^�^�� Ǖ �Z3�T0 k� �PN�TN�1	�"qe1�t B  ��3    � �8A\�q]ÚG�[�OK���$[ˤA^�^�� Ö �Z3�T0 k� �PN�TN�1	�"qe1�t B  ��3    � �8A\�q]��C�[�OK���$[ǤA^�^�� �� �Z3�T0 k� �TN�XN�1	�"qe1�t B  ��3    � �8A\�q]��;�[�OK���$[ãA^�^�� �� �Z3�T0 k� �TO�XO�1	�"qe1�t B  ��3    � �8A\�q]��7�[�OK���$[��A^�^�� �� �Z3�T0 k� �TO�XO�1	�"qe1�t B  ��3    � �8A\�q]��3�[�OK���$[��A^�^�� �� �Z3�T0 k� �TO�XO�1	�"qe1�t B  ��3    � �8A\�q]��/�[�OK���([��A^�^�� �� �Z3�T0 k� �XO�\O�1	�"qe1�t B  ��3    � �8A\�q]��'�[�PK���([��A^�^�� �� �Z3�T0 k� �XO�\O�1	�"qe1�t B  ��3    � �8A\�q]��#�[�PK���([��A^�^�� �� �Z3�T0 k� �XO�\O�1	�"qe1�t B  ��3    � �8A\�q]���[�PK���([��A^�^�� �� �Z3�T0 k� �XO�\O�1	�"qe1�t B  ��3    �  �8A\�q]���[�PK���([��A^�^�� �� �Z3�T0 k� �\O�`O�1	�"qe1�t B  ��3    � !�8A\�q]���[�PK���([��A^�^�� �� �Z3�T0 k� �\O�`O�1	�"qe1�t B  ��3    � "�8A\�q]���[�PK���([��A^�^�� �� �Z3�T0 k� �\O�`O�1	�"qe1�t B  ��3    � #�8A\�q]���[�PK���( [��A^�^�� �� �Z3�T0 k� �`O�dO�1	�"qe1�t B  ��3    � $�8A\�q]���[�PK���(![��A^�^�� �� �Z3�T0 k� �`O�dO�1	�"qe1�t B  ��3    � %�8A\�q]���[�PK���(![��A^�^�� �� �Z3�T0 k� �`P�dP�1	�"qe1�t B  ��3    � &�8A\�q]���[�PK���("[��A^�^�� � �Z3�T0 k� �`P�dP�1	�"qe1�t B  ��3    � '�8A\�q]{���[�PK���("[��A^�^�� {� �Z3�T0 k� �dP�hP�1	�"qe1�t B  ��3    � (�8A\�q]w���[�PK��"(#[��A^�^�� w� �bs�T0 k� �dP�hP�1	�"qe1�t B  ��3    � (�8A\�q]s���[�PK��"(#[��A^�^�� s� �bs�T0 k� �dP�hP�1	�"qe1�t B  ��3    � (�8A\�q]o���[�PK��"($[��A^�^�� o� �bs�T0 k� �dP�hP�1	�"qe1�t B  ��3    � (�8A\�q]k���[�QK��"($[��A^�^�� k� �bs�T0 k� �dP�hP�1	�"qe1�t B  ��3    � )�8A\�q]g���[�QK�"(%[��A^�^�� g� �bs�T0 k� �hP�lP�1	�"qe1�t B  ��3    � )�8A\�q]c���[�QK�"(%[��A^�^�� c� �bs�T0 k� �hP�lP�1	�"qe1�t B  ��3    � )�8A\�q]_���[�QK{�"(&[àA^�^�� _� �bs�T0 k� �hP�lP�1	�"qe1�t B  ��3    � )�8A\�q][���[�QK{�"(&[àA^�^�� [� �	bs�T0 k� �hP�lP�1	�"qe1�t B  ��3    � )�8A\�q]W���[�QKw�"(&[àA^�^�� W� �	bs�T0 k� �lP�pP�1	�"qe1�t B  ��3    � )�8A\�q]W���[�QKw�"('[àA^�^�� W� |	bs�T0 k� �lP�pP�1	�"qe1�t B  ��3    � )�8A\�q]S���[�QKs�"('[àA^|^�� S� |	bs�T0 k� �lP�pP�1	�"qe1�t B  ��3    � )�8A\�q]O���[�QKs��,([ǠA^x^�� O� x	Z3�T0 k� �lP�pP�1	�"qe1�t B  ��3    � )�8A\�q]K���[�QKw��,([ǠA^x^�� K� t	Z3�T0 k� �lQ�pQ�1	�"qe1�t B  ��3    � )�8A\|q]G���[�QKw��,)[ǟA^t^�� G� t	Z3�T0 k� �pQ�tQ�1	�"qe1�t B  ��3    � )�8A\|q]G���[�QKw��,)[ǟA^p^�� C� p
Z3�T0 k� �pQ�tQ�1	�"qe1�t B  ��3    � )�8A\xq]C���[�QKw��,)[˟A^p^�� C� p
Z3�T0 k� �pQ�tQ�1	�"qe1�t B  ��3    � )�8A\tq]?���[�QK{��,*[˟A^l^�� ?� l
Z3�T0 k� �pQ�tQ�1	�"qe1�t B  ��3    � )�8A\pq];���[�QK{��,*[˟A^h^�� ;� l
Z3�T0 k� �pQ�tQ�1	�"qe1�t B  ��3    � )�8A\lq]7���[�QK{��,+[˟A^h^�� 7� h
Z3�T0 k� �tQ�xQ�1	�"qe1�t B  ��3    � )�8A\lq]7���[�RK{��,+[˟A^d^�� 7� d
Z3�T0 k� �tQ�xQ�1	�"qe1�t B  ��3    � *�8A\hq]3���[�RK��,+[ϟA^d^�� 3� d
Z3�T0 k� �tQ�xQ�1	�"qe1�t B  ��3    � *�8A\dq]/���[�RK��,,[ϟA^`^�� /� `
Z3�T0 k� �tQ�xQ�1	�"qe1�t B  ��3    � *�8A\`q]/���[�RK�",,,[ϟA^`^�� /� `b��T0 k� �tQ�xQ�1	�"qe1�t B  ��3    � *�8A\`q]+���[�RK�",,-[ϟA^\^�� +� \b��T0 k� �tQ�xQ�1	�"qe1�t B  ��3    � *�8A\\q]'���[�RK�",,-[ϟA^\^�� '� \b��T0 k� �xQ�|Q�1	�"qe1�t B  ��3    � *�8A\Xq]'���[�RK��",,-[ӟA^X^�� '� Xb��T0 k� �xQ�|Q�1	�"qe1�t B  ��3    � *�8A\Xq]#���[�RK��",,.[ӟA^T^�� #� Xb��T0 k� �xQ�|Q�1	�"qe1�t B  ��3    � *�8A\Tq]���[�RK��",,.[ӟA^T^�� � Tb��T0 k� �xQ�|Q�1	�"qe1�t B  ��3    � *�8A\Pq]���[�RK��",,.[ӟA^P^�� � Tb��T0 k� �xQ�|Q�1	�"qe1�t B  ��3    � *�8A\Pq]���[�RK��",,/[ӟA^P^�� � Pb��T0 k� �xQ�|Q�1	�"qe1�t B  ��3    � *�8A\Lq]���[�RK��",,/[ӟA^L^�� � Pb��T0 k� �|R��R�1	�"qe1�t B  ��3    � *�8A\Hq]���[�RK��",,/[ןA^L^�� � Lb��T0 k� �|R��R�1	�"qe1�t B  ��3    � *�8A\Hq]���[�RK��",,0[ןA^H^�� � Lb��T0 k� �|R��R�1	�"qe1�t B  ��3    � *�8A\Dq]���[�RK���,0[ןA^H^�� � LZ3�T0 k� �|R��R�1	�"qe1�t B  ��3    � *�8A\@q]���[�RK���,0[ןA^H^�� � HZ3�T0 k� �|R��R�1	�"qe1�t B  ��3    � *�8A\@q]���[�RK���,0[ןA^D^�� � HZ3�T0 k� �|R��R�1	�"qe1�t B  ��3    � *�8A\<q]���[�RK���,1[ןA^D^�� � DZ3�T0 k� �|R��R�1	�"qe1�t B  ��3    � *�8A\<q]���[�RK���,1[۟A^@^�� � DZ3�T0 k� ��R��R�1	�"qe1�t B  ��3    � *�8A\8q]���[�RK���,1[۟A^@^�� � @Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � *�8A\8q]���[�RK���,2[۟A^<^�� � @Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � *�8A\4q]��[�SK���,2[۟A^<^�� � @Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\4q\��{�[�SK���02[۟A^<^���� <Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\0q\��{�[�SK���02[۟A^8^���� <Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\,q\��w�[�SK���03[۟A^8^���� <Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\,q\��w�[�SK���03[ߟA^4^���� 8Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\(q\��s�[�SK���03[ߟA^4^���� 8Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\(q\��s�[�SK���03[ߟA^4^���� 4Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\$q\�o�[�SK���04[ߟA^0^���� 4Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\$q\�o�[�SK���04[ߟA^0^��� 4Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\ q\�k�[�SK���04[ߟA^,^��� 0Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\ q\�k�[�SK���04[ߟA^,^��� 0Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\ q\�k�[�SK���05[ߟA^,^��� 0Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\q\�g�[�SK��<05[�A^(^��� ,Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\q\�g�[�SK��<05[�A^(^��� ,Z3�T0 k� ��R��R�1	�"qe1�t B  ��3    � +�8A\q\�c�[�SK��<,5[�A^(^��� ,Z3�T0 k� ��S��S�1	�"qe1�t B  ��3    � +�8A\q\�c�[�SK��<,6[�A^$^��� ,Z3�T0 k� ��S��S�1	�"qe1�t B  ��3    � +�8A\q\�_�[�SK��<,6[�A^$^��� (Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\�_�[�SK���,6[�A^$^��� (Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ߚ_�[�SK���,5[�A^ ^��� (Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ߚ[�[�SK���,5[�A^ ^��� $Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ߚ[�[�SK���(5[�A^ ^��ߝ $Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ۚW�[�SK���(5[�A^ ^��ߝ $Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ۚW�[�SK���(4[�A^^��۝  Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ۚW�[�SK���(4[�A^^��۝  Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ךS�[�SK���(3[�A^^��۝  Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ךS�[�SK���(3[�A^^��ם  Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ךS�[�SK���$2[�A^^��ם Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ӚO�[�SK���$2[�A^^��ם Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � +�8A\q\ӚO�[�TK���$1[�A^^��ӝ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � ,�8A\ q\ϚK�[�TK���$1[�A^^��ӝ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � ,�8A\ q\ϚK�[�TK���$1[�A^^��ӝ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � ,�8A\ q\ϚK�[�TK���$0[�A^^��ϝ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � ,�8A[�q\ϚG�[�TK���$0[�A^^��ϝ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 	   � ,�8A[�q\˚G�[�TK���$0[�A^^��ϝ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\˚G�[�TK��� /[�A^^��˝ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\˚G�[�TK��� /[�A^^��˝ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\ǚC�[�TK��� .[�A^^��˝ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\ǚC�[�TK��� .[�A^^��˝ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\ǚC�[�TK��� .[�A^^��Ǟ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\Ú?�[�TK��� -[�A^^��Ǟ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\Ú?�[�TK��� -[�A^^��Ǟ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\Ú?�[�TK��� -[�A^^��Ǟ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\Ú;�[�TK���,[�A^^��Þ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\��;�[�TK���,[�A^^��Þ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\��;�[�TK���,[�A^^��Þ Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\��;�[�TK���+[�A^^���� Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\��7�[�TK���+[�A^^���� Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\��7�[�TK���+[�A^^���� Z3�T0 k� ��S��S�1	�"qe1�t B  ��3 
   � ,�8A[�q\��7�[�TK���*[�A^^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3 
   � ,�8A[�q\��7�[�TK���*[�A^^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3 
   � ,�8A[�q\��3�[�TK���*[�A^^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3 
   � ,�8A[�q\��3�[�TK���*[�A^^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3 
   � ,�8A[�q\��3�[�TK���)[�A^ ^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3 
   � ,�8A[�q\��3�[�TK���)[�A^ ^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3 
   � ,�8A[�q\��3�[�TK���)[�A^ ^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��/�[�TK���([�A^ ^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��/�[�TK���([�A^ ^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��/�[�TK���([�A]�^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��/�[�TK���([�A]�^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��+�[�TK���'[�A]�^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��+�[�TK���'[�A]�^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��+�[�TK���'[�A]�^���� Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��+�[�TK���'[�A]�^����  Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��+�[�TK���&[�A]�^����  Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��'�[�TK���&[�A]�^����  Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��'�[�TK���&[�A]�^����  Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8A[�q\��'�[�TK���&[�A]�^����  Z3�T0 k� ��T��T�1	�"qe1�t B  ��3    � ,�8@�x � �F pX b|  �`@�`x�tF ��T XZc� T0 k� �8F�<F�1	�"qe1�t B  ��/    �  @�x � �F pX b|  �`@�`x�tF ��T XZc� T0 k� �8F�<F�1	�"qe1�t B  /�/    �  @�x � �F pX b|  �`@�`x�tF ��T XZc� T0 k� �XF�\F�1	�"qe1�t B  ��/ 	   �  @�x ��F pX b|  �`@�`x�tF ��T XZc� T0 k� �dF�hF�1	�"qe1�t B  ��/ 	   �  @�x ��F pX b|  �`@�`x�tF ��T XZc� T0 k� �lF�pF�1	�"qe1�t B  ��/ 	   �  @�x ��F pX b|  �`@�`x�tF ��T XZc�T0 k� �tF�xF�1	�"qe1�t B  ��/ 	   �  @�x ��F pX b|   �`@�`x�tF ��T XZc�T0 k� �|F��F�1	�"qe1�t B  ��/ 	   �  @�w ��F pX b|   �`@�`x�tF ��S�XZc�T0 k� �F��F�1	�"qe1�t B  ��/ 	   �  CCw�FBpX b|$ S`A`x�tF�3�XZc�T0 k� �F��F�1	�"qe1�t B  ��/ 	   �  CCw"�FBpX |$ S`A`w�tF�3�XZc�T0 k� �F��F�1	�"qe1�t B  ��/ 	   �  CCv"�FBpX |$ S`A`w�tF�3�W_��T0 k� �F��F�1	�"qe1�t B  ��/ 	   �  CCv"�FBpX |$ S`A`w�tF�3�W_��T0 k� �F��F�1	�"qe1�t B  ��/ 	   �  CCu"�FBpX |( S`A\w�tF�3�W_��T0 k� �H��H�1	�"qe1�t B  ��* 	   �   CCuS"�FBpX |( �`C�\w�tFS���W_��T0 k� ��F��F�1	�"qe1�t B  ��* 	   � ! CCtS"�F�pXB|( �`C�\wCtFS���V_��	T0 k� ��C��C�1	�"qe1�t B  ��* 	   � " CCtS"�F�pWB|( �`C�\vCtFS���VZ��
T0 k� ��B��B�1	�"qe1�t B  ��* 	   � # E3sS"�F�pWB|( �`C�XvCtFS���VZ��T0 k� ��A��A�1	�"qe1�t B  ��* 	   � $ E3rS"�F�pWB|( �`C�XvCtFS���UZ��T0 k� ��?��?�1	�"qe1�t B  ��* 	   � % E3q��F�pWB|( �`E�XuCtF3���UZ��T0 k� ��?��?�1	�"qe1�t B  ��* 	   � & E3p��F�pWB|( 3`E�Tu�tF3���TZ��T0 k� ��>��>�1	�"qe1�t B  ��* 	   � ' E3p��F�pW�|( 3\E�Tt�tF3���TZ��T0 k� ��>��>�1	�"qe1�t B  ��* 	   � ( E#o��F�pW�|( 3\E�Pt�tF3���SZ��T0 k� ��=��=�1	�"qe1�t B  ��* 	   � ) E#m��F�pW�|( 3XE�Ls�tF3���RZ��T0 k� ��<��<�1	�"qe1�t B  ��* 	   � * E#l� �F�pW�|( 3XE�Ls�tF3��QZ��T0 k� ��=��=�1	�"qe1�t B  ��* 	   � * E#k� �F�pW�|( 3TE�Ls�tF3��PZ��T0 k� � =�=�1	�"qe1�t B  ��* 	   � * B�i� �FRpW�|( 3TE�Hr�tF3��PZ��T0 k� �>�>�1	�"qe1�t B  ��* 	   � * B�h�  DRpW�|( CPE�Hr�tF3��OZ��T0 k� �>�>�1	�"qe1�t B  ��*    � * B�gc CRpW�|( CPC�Dr�tFC��NZ��T0 k� �=�=�1	�"qe1�t B  ��*    � * B�dc�ARlW�|( CLC�@qStFC��LZ��T0 k� �;�;�1	�"qe1�t B  �*    � * E#cc�@RlW�|( CLC�<qStFC��LZ��T0 k� �;�;�1	�"qe1�t B  �*    � * E#bc�?RlW�|( CLC�8qStFC���KZ��T0 k� �?�?�1	�"qe1�t B  ��*    � * E#ac�>RlW�|( CLC�8qStFS���JZ��T0 k� �A�A�1	�"qe1�t B  ��*    � * E#`c� =RlW�|( CLC�4pStFS���IZ��T0 k� �B�B�1	�"qe1�t B  ��*    � * E#_c�$;RlW�|( CLC�4ptFS���HZ��T0 k� �C�C�1	�"qe1�t B  ��*    � * E#]c�(:RhW�|( CLC�0ptFS���GZ��T0 k� �C�C�1	�"qe1�t B  ��*    � * E#\��,9RhV�|( CLC�0ptFS���GZ��T0 k� ��C� C�1	�"qe1�t B  ��*    � * @c[��08RhV�|( SHC�0ptFC���FZ��T0 k� ��C��C�1	�"qe1�t B  ��*    � * @cY��86RhV�|( SHC�,ptFC���DZ��T0 k� ��A��A�1	�"qe1�t B  ��*    � * @cX� �<5RhV�|( SDC�,p �tFC���DZ��T0 k� ��A��A�1	�"qe1�t B  ��*    � * @cW� �@4RhV�|( SDC�,p �tFC���CZ��T0 k� ��A��A�1	�"qe1�t B  ��*    � * @cV� �D3RhV�|( SDC�,p �tFC���BZ��T0 k� ��@��@�1	�"qe1�t B  ��*    � * @cU� �H3RdV�|( S@C�(p �tF3���AZ��T0 k� ��?��?�1	�"qe1�t B  ��*   � * @cT���L2RdV�|( S@C�(p �tF3���AZ��T0 k� ��>��>�1	�"qe1�t B  ��*    � * @cS���P1RdV�|( S@C�(p �tF3���@Z��T0 k� ��>��>�1	�"qe1�t B  ��*   � * @cR���T0RdV�|( S@C�(p ctF3���?Z��T0 k� ��=��=�1	�"qe1�t B  ��*    � * @cQ���X/RdV�|( S@A�(p cxF3���?Z��T0 k� ��<��<�1	�"qe1�t B  ��*    � * @cP���X.RdV�|( c<A�(p cxG3���>Z��T0 k� ��<��<�1	�"qe1�t B  ��*    � * @cO��
�\-RdV�|( c<A�(p cxG3���=Z��T0 k� ��;��;�1	�"qe1�t B  ��*    � * @cN��
�`,RdV�|( c<A�(p cxGC���=Z��T0 k� ��:��:�1	�"qe1�t B  ��*    � * @cM��
�d,R`V�|( c<A�(p�xGC���<Z��T0 k� ��:��:�1	�"qe1�t B  ��*    � * @cL��
�h+R`V�|( c<A�(p�xGC���;Z��T0 k� ��9��9�1	�"qe1�t B  ��*    � * @cK��	�l*R`V�|( c<A�(p�|HC���;Z��T0 k� ��8��8�1	�"qe1�t B  ��*    � * @cK��	�p)R`V�|( c<A�(p�|HC���:Z��T0 k� ��8��8�1	�"qe1�t B  ��*    � * @cJ��	�t(R`V�|( c<A�(p�|H3���:Z��T0 k� ��7��7�1	�"qe1�t B  ��*    � * @cI��	�x(R`V�|( �<A�(p�I3|��9Z��T0 k� ��7��7�1	�"qe1�t B  ��*    � * @cH���|'R`V�|( �<A�(p�I3|��8Z��T0 k� ��6��6�1	�"qe1�t B  ��*    � * @cG����&R`V�|( �<BC(p�J3|��8Z��T0 k� ��5��5�1	�"qe1�t B  ��*    � * @cG����%R`V�|( �<BC(p�J3|��7Z��T0 k� ��5��5�1	�"qe1�t B  ��*    � * @c F����%R`V�|( �<BC(p�K#|��7Z��T0 k� ��4��4�1	�"qe1�t B  ��*    � * @c E����$R\V�|( C<BC(p�L#|��6Z��T0 k� ��4��4�1	�"qe1�t B  ��*    � * @c D����#R\V�|( C<BC(p�L#|��6Z� T0 k� ��3��3�1	�"qe1�t B  ��*    � * @c D����#R\V�|( C<@(p�M#|��5Z� T0 k� ��3��3�1	�"qe1�t B  ��*    � * @c C����#R\V�|( C<@(p�N#���5Z� T0 k� ��2��2�1	�"qe1�t B  ��*   � *                                                                                                                                                                             � � �  �  �  c A�  �J����   �      6 \��L. ]�)) � �� D}          � ��@     Jw ��@    ��               
    ��         7�  �  ���   8	          ��~�          � �А    ��~� �А    ��                  �         u   �  ���   0	


 
          t��          ��     toy �j    o��    y y           �         �     ���   8		          Ut�            �7P     Ut� �7P                    
 A           �p     ���   @

(          ��           . �#�     �� �#�                      
             ~�  �  ���   H

 

           ��  ��      B�
��      ���
��                              ���                �  ���    8

 '             ^�� ??   V Ŀ�     _~ �+g    �`��    v v      	 Z           \�&  .3 ��`  0

           {w / /     j �֐     {�� ��P    �� �              Z           �`�   	  ��@  (
           ["�  > >    ~��     ["��      ��    \ \     < Z           � �   
 ��A  8�          c,=  $ $      �s�     c,=s�                      	 Z          	 �     ��@   (
            7�        �-�     7�-�                       Z          
 ~      ��H   P
B          2���
      �x�     2��z�     ���                     ���C                ��@    8		 1                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          Gz�  ��        �9  � Gz�9  �                       x                j  �    
   �                          G    ��        �       G             "                                                �                          � � � � ��
 � ���          
  	     
 � 
  03� ���[       #� `o� $d p� �d 0n` �� n� �� p����< ����J ����X � �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0� ���� ����� � 
�< V� 
� W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����    *���   ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j B���
��
��"    B�j l �  B �
� �  �  
�  7    ��     �       t��  ��     � �       7    ��     �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �/B	B      ��7T ���        � �T ���        �        ��        �        ��        �    �     1�� ���        ��                         ��q < 	�� �                                    �                 ����            
 7
���%��   *   F �            21/47 (44%) rchuk y    4:40                                                                        3  3     �SC. �k C6 �HC#h C"+(B� �@ B� �cV!&cZ16	c^7. 
cbA cc0. cd)J� �J� � �CBCR �kjE � kpE � k� �
k� � � k� �c�0 � c�( �	� � �	� � �� � �� � �c~) � c�9 �c� �c� �  � � !� �""� � #"� �$� � �%
�&"�: '"�L("�:)*�I �*"� � +"� �,� � �-
� � ."M ~ �/"0 � �0"$ � � 1"? � 2*M& � 3*KN �4*6~ � 5*OvH  *&~H  *&~ � 8*OvH  *&~ � :*Kf � ;*^ � <*KV � =*Pv � >*Of � **~                                                                                                                                                                                                                         �� R              @ 
      Q �     c P E d  ��        
            �������������������������������������� ���������	�
��������                                                                                          ��    �cc�� ��������������������������������������������������������   �4, E�  ��@P���$���f������                                                                                                                                                                                                                                                                                                                                           @#�                                                                                                                                                                                                                                             	       \        ��  9<�J      J  	                           ������������������������������������������������������                                                                                                                                              �  �                  �}    ��                     ����������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� �������������������             x                       
   /     �  L�J      ,�                             ������������������������������������������������������                                                                      	                                                                   �    �              �          ��                 	 	 �������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ����                                                                                                                                                                                                                                                                        
                              	                    �             


           �   }�         wwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwww 0 I =                                 � :��{ �o�                                                                                                                                                                                                                                                                                   �1n  
)�        d      l            m      d      e      `      l                                                                                                                                                                                                                                                                                                                                                                                                         � (� �  � (��  � ��  � @��  � #��  � ��  �����������������������f�����.�����R������������                ���D : [ 
         �   & AG� �   �   
              �                                                                                                                                                                                                                                                                                                                                      p G I   �                       !��                                                                                                                                                                                                                            Y��   �� � ��      �� ]      ����������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� ��������������������������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ����             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    *      =      G                       e     �  �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ��  �� �    � �N ^$   �̞   0  ��   )   �   �   ���T     �f ��        p���� ��   p���� �$ ^h  ��     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h   ����� ��   ����� �$ ^$ /   �         ��       /   �����������J�������������� > �/ �  ��  �         ��   ���` o� #� �� o� #� �$ ^$         ��  *             ��L�����         ����J  ��  yf  y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                          �  �_ <� ���\~~����    UUU�333����~~~~����~~~~����    _�� 3�p �<� �?� �3��|��p��<�                                          �                           �   S  <  <  �  ��  S�<~~~�����~~~����~~~~����~~~~����~~~~����~~~~����~~~~����~~|����3~|3�����~|�<���<~~|;�����~~�3���    �   p  �   �   ��  �p  <�                         _  33?   S�  S�  S�  S�  S�  S�  S�  S3~~~~����~~~~����~~~~��������3333~|5 ��P ~�P ��P ~�P ��P ��P 33P <~| S�� S�~ S�� S�~ S�� S�� S33<~ �����~ �<� |?�~������<~33<�335 33? _      ~~~~����~~~~����  UU                   �        UUUU                            UUP          �                   UUU                            UUU�                            ~~~~                           wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         7v` weV "fff"O�p"��p"��p"�p3�}p-��p=��p|� }�  }�  ��  ��  ��  ��  �  �  �  �  �  "              `  eV  fff O�  ��  ��  �  �} �� �� ��  |�  }�  ��    =   }   =   =              �������}�}�}�ww~r�� ∈�������������������}�� }�� ��� ��� ����   �   �   �   �   �   �   �   C""42""#2""#2""#2""#s3342"""3333    p   p   p   p   p   p   p    ��������� ��� }�� ��  ��  ����  ��  ��  ��  ��  ��  ��  ��                          � �� ��    "               wvf wfU 7Of`w��f"�� "�p-�}p���� ��� ����x��	�� �� �� "�        f  U` f` f` �p w���� `  eV  ff  O�  ��  �� ����}�                �  �  ��  �            �  �  �   �  ��  �                     �  �  �   � `  eV  ff  O�  ��  ��  ����}���������������p	���         `  eV  ff  O�  ��  ��  ���}�     �  �  �   �  ��  �   �            ��  ��  �   ��  �   ���������������p	���                    3333UUUU                        wwww                    333333333333333333333   w  G� ws@ ws� ws$7w@wwww"                               ����������� ��� �� ��  �    `  eV  ff  O�  ��  ��  � ��}�            """"                  w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 " ""   "" "!  "" "  """ !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "!  "! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �            " ""   "" "!  "" "  """ !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                              	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                                   ��                  �                        ���� ��� ����            �   �   �   D   E�  U�  UO                         "  "  "                                                                                                                                                                 �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                   �   �                      �������  ���    ��   �  ���� �   �             �   ��  ��  ��  �  �   ��  ��                            ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                                  �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �   �                                    ��                                ��                                              �    �     �                         � ���� ��   � � �                            ����                  �   �� �       �  �  ��  �   �   �   �                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                     �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                �   ���                        � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    �   �   �                       ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ���                                                                                                                                                                                                                    �� �����ݼڜ��ک��ک��z�	��� 
�� 
�� 	�� ̘ ɪ  ��  �  �� �� ������������ ���  � � � �� �� ������ ��                      �   ��  ��  �̰ ��� ��˰�̻��̻���������ˉ�U��EP�ET �I� ٕ  �D� �L� ��� ��" ����/�"�"�""�����                         ��� �� ���"� ��   �� �        � ��� ��� ��  �                �   �     �   �               �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                                       " "  ""��",ʜ"�������  �  ��              ""  "�  ,ˠ "ʛ 򨻿��D 4U� 3D�D�EET4U�TET�EUH��UI��Y ��T   T�� H�  ������̻��̻��̻��ɻ�˚���������ɏ �����  ��  ��                �   �̰ ��� �ع���ة��ڋ̻ز���"�������"� "/  �"� ".� ��                            �   ��   ��                               �   ��   ��                  �� ������ ��      �   /   "�  "�  "�  ��                          �   O   T     ��                                 � ���� ��   � � �                                                                                                                                           �   �  �  �  	�  �  EH  ET DU CE DD4 DD3 DC0 �3 ɰ �  ,�  +�  "/  ������ � ̹�p�˚��̹���ː�̼�̻���ۜ��۩�ݍ���=��J�ܰT�� EJ�0 EJ� I�  ��  �"  ""  "/  "�� ���                    ̰ ̻ ̻	���̚�wˢ �+���"����"��"  �   �    �   �" �"� "������     �     �� �� ��
��׊��w٪�|��������            "   "   "       �         �        �   �     �       �   �   �   �   �      �                    ��� ���� �� ��  �  �  �   �                                         ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                     � 
��	�˽���w��{k��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            �  �  �  ��  �           ��  ��� �"" ""@  "D   U@  UP  U@  D   �   "   "   "/� �����               �   �   �  �  �  �  �   �   �                                       �  ���
�� ��  �   "  "  ""  ""     DH  UT@ DU@ 4ET 3ED@ D�@ ˰ �� �� 
˰  ̰  "   ""  ""  "    �   �   �   �                               �    �    ��                        �  �  �                                                                       �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �                       �   �   �               "   "   "       �         �        �   �     �       �   �   �   �   �      �                    ��� ���� ��                        ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                                          	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                           �  �   �   �   �   �  �        � �� ����   �              ���� ����                     ��     �                     �  �  �  �  �  ��  �                       �   ���                            �   �                                                                                                                    �� ̻ ��˛��  �� �˚̻���ۚ����I���䘼�^���^�٘�:�^�� ^�� D�( �) �) �) ��) ˹� ț�+��,��,����  �𫝝 ��� �ɍ ��ݨ��ډ�݊�� ��D@ �D�  J�� ݩ� ��� �ۻ �ک �ڹ�ɻ��̸���������� ����������            �   ��  ��  ��  ��  ��                                          �� ��� ��� ��  �                         �   �           �   �     �   �               �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""������������������������""""������ADAIA�A""""�������I�A�A�A""""�����DD�I""""�������DAADAI""""������IDA��""""��������DD��I�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD������������������������3333DDDD�A�AM�M�DM��M334CDDDD�A�AM�M�DDM����3333DDDDDM����DD�����3333DDDDMAM��D�DDM�����3333DDDDDD����M��DM�����3333DDDD������������DD������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��           	 
          
        ((((((( 
	(((( ����������������             ! " # $ % & '   ( $ % ) ! " # * ('(&(%($(#("(! (((���������������� + , -   . / 0 1  	 2         3       4 (((((((2	10/(.(-(,(+���������������� 5 6   7   8 9 1 :   $ % ) ! " #   ; ) ! " # $ % ) (#("(!()(%($ :198(((7(6(5����������������    <     = 8 0 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>108(=((( (<���������������� L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L����������������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7����������������  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(�����������������333333333333333333333333333333333333333333333333333333333333����  
�fD
��L���"��������������������D" � j  "  B   J jF� ����
��� �����
���� ����
��� �����
��� 0 q����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqSC. �k C6 �HC#h C"+(B� �@ B� �cV!&cZ16	c^7. 
cbA cc0. cd)J� �J� � �CBCR �kjE � kpE � k� �
k� � � k� �c�0 � c�( �	� � �	� � �� � �� � �c~) � c�9 �c� �c� �  � � !� �""� � #"� �$� � �%
�&"�: '"�L("�:)*�I �*"� � +"� �,� � �-
� � ."M ~ �/"0 � �0"$ � � 1"? � 2*M& � 3*KN �4*6~ � 5*OvH  *&~H  *&~ � 8*OvH  *&~ � :*Kf � ;*^ � <*KV � =*Pv � >*Of � **~3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0�������������������������������������������7�G�Z�Y��<�[�T�J�O�T� � � � � � � � � �:�>�/�������������������������������������������.�G�R�K��2�G�]�K�X�I�N�[�Q� � � � � � �,�>�0�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������:�>�/� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                