GST@�                                                           �j�                                                                  d     �        � 2�������J����������    ����        |�      #    ����                                d8<n    �  ?     ����  �
fD�
�L���"����D"� j   " B   J  jF�"    "�j* ,  �����
�"     �j@ �    ��
  R�                                                                              ����������������������������������       ��    ?b 0Qb 5 814  4c c   c       	 

    
   	  
      ��G 4�  ( �(                 nn 
)1         :88�����������������������������������������������������������������������������������������������������������������������������o  b  o   1  +    '           �                  	  7  V  	                  Y  !          := �����������������������������������������������������������������������������                                D              @  &   v   �                                                                                 '    
)n1n  !Y    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    	`aA�aF"�f[�|( ��Q@ ��h�:��T��T0 k� ����U8D"!S�d    ��   ��� �	`aA�aF#�d_�|( ��Q@ Рi�;��U��T0 k� �����U8D"!S�d    ��   ��� �	``A�bF%�c�c�|( ��R@ Фk�<s�U��T0 k� ��~��~U8D"!S�d    ��   ��� �	`_A�bF (� a�o�|( � S@ Шm�?s�V��
T0 k� ��|��|U8D"!S�d    ��   ��� �	$\^A�bE�$*��`�w�|( �T@ Ьn�@s�V��T0 k� ��{��{U8D"!S�d    ��   ��� �	$\^C��aE�(+��^�{�|( �T@ аo�Bs�V��T0 k� ��{��{U8D"!S�d    ��   ��� �	$\]C��bE�,-��]���|( �U@ дp�Cs�V��T0 k� ��z��zU8D"!S�d    ��   ��� �	$\]C��bE�,.�\���|( �V@ иq�Ds�U��T0 k� ��z��zU8D"!S�d    ��   ��� �	$\\C��bE�41�Y���|( �W@ ��r�Gs�T���T0 k� ��z��zU8D"!S�d    ��   ��� �	\[C��bE�83�X���|( �X@ ��s�H��T���T0 k� ��z��zU8D"!S�d    ��   ��� �	\[C��cE�<4�V���|( �X@ ��t�J��S���T0 k� �{z�zU8D"!S�d    ��   ��� �	\[C��cE�@6�U���|( �Y@ ��t�K��S���T0 k� �oz�szU8D"!S�d    ��   ��� �	`ZC��cE�D7�S���|( �Y@ ��u�L��R���T0 k� �cz�gzU8D"!S�d    ��   ��� �	`ZC��bE�H8�Rѷ�|( �Y@ ��v�M��Q���T0 k� �Wz�[zU8D"!S�d    ��   ��� �	$`ZC��bE�P:�Pѻ�|( �Z@ ��v�N��P���T0 k� �Kz�OzU8D"!S�d    ��   ��� �	$`YC��bE�X<�M���|( �\@ ��w�Q��O���T0 k� �3z�7zU8D"!S�d    ��   ��� �	$`YC��bE�\=�L���|( �]@ ��w�R��N���T0 k� �'z�+zU8D"!S�d    ��   ��� �	$\YC��bE�`?��J���|( �^@ ��x�S��M���T0 k� �z�zU8D"!S�d    ��   ��� ��\XC��aE�h@��I���|( �_@ ��x�T��L���T0 k� �z�zU8D"!S�d    ��   ��� ��\XC��aE�lA��G���|( �_@ ��x�U��K���T0 k� �z�zU8D"!S�d    ��   ��� ��\XC��`E�pB��F���|( �`@ ��x�V��J���T0 k� ��z��zU8D"!S�d    ��   ��� ��\XE3�`E�tC��D���|( �a@ � x�W��I���T0 k� ��z��zU8D"!S�d    ��   ��� ��XXE3�_E�|C��C���|( �b@ �x�X��Gc��T0 k� ��z��zU8D"!S�d    ��   ��� � �XXE3�_E��D��A���|( �c@ qx�Y��Fc��T0 k� ��z��zU8D"!S�d    ��   ��� � �XXE3�^E��E��@���|( �d@ qx�Z��Ec��T0 k� ��z��zU8D"!S�d    ��   ��� � �XXE3�]E��F��?��|( �d@ qx�[s�Dc��T0 k� ��z��zU8D"!S�d    ��O   ��� � �TXE3�]E��F��=��|( �e@ qx�\s�Bc��T0 k� ��z��zU8D"!S�d    ��O   ��� � �TXCC�\E��G��<��|( �f@ q x�]s�Ac��T0 k� ��z��zU8D"!S�d    ��O   ��� ��TXCC�[E��G��;��|( �g@ �$w�^s�@c��T0 k� ��z��zU8D"!S�d    �O    ��� ��PXCC�ZE��H �9��|( �g@ �,w�^s�>c��T0 k� ��z��zU8D"!S�d    �O    ��� ��PYCC�Y@��H �8�'�|( �h@ �0w�^c�=c��T0 k� ��z��zU8D"!S�d    ��O    ��� ��PYCC�Y@��I �7�+�|( �i@ �4v�]c�;c��T0 k� �z��zU8D"!S�d    ��O    ��� ��LY@��X@��I �6r3�|( � i@ �8v�]c�:c��T0 k� �sz�wzU8D"!S�d    ��O    ��� ��LY@��X@��I �5r7�|( �j@ �<u�]c�9c��T0 k� �g{�k{U8D"!S�d    ��O    ��� ��LY@��X@��I �3r?�|( �k@ �Du�]c�7c��T0 k� �[{�_{U8D"!S�d    ��O    ��� ��HZ@��X@��H �2rC�|( �l@ �Ht�\3�6c��T0 k� �O{�S{U8D"!S�d    ��O    ��� ��HZ@��X@��H �1rG�|( �l@ �Ls�\3�4c��T0 k� �G{�K{U8D"!S�d    ��O    ��� �HZ@��X@��H �0rO�|( �m@ �Ps�\3�3c��T0 k� �;{�?{U8D"!S�d    ��O    ��� �DZ@��X@��H �/rS�|( �m@ �Tr�\3�1c��T0 k� �/{�3{U8D"!S�d    ��O    ��� �DZ@��X@��G �.r[�|( �n@ �Xq�\3�/c��T0 k� �#{�'{U8D"!S�d    ��O    ��� �DZ@��X@��G �-r_�|( �o@ �\p�[3�.c��T0 k� �{�{U8D"!S�d    ��O    ��� �@[@��X@��G �,rc�|( �o@ �`o�[3�,c��T0 k� �{�{U8D"!S�d    ��O    ��� �@[@��X@��G �+rg�|( �p@ �dn�[3�+c��T0 k� �{�{U8D"!S�d    ��O    ��� �@[@��X@��F �*bo�|( �q@ �hm�[C�)c��T0 k� ��{��{U8D"!S�d    ��O    ��� �@[@��X@��F �)bs�|( �q@ �ll�[C�'c��T0 k� ��{��{U8D"!S�d    ��O    ��� �<[@��X@��F �(bw�|( �r@ �pk�[C�&c��T0 k� ��{��{U8D"!S�d    ��O    ��� �<[@��X@��F �'b{�|( #�r@ �tj�ZC�$c��T0 k� ��{��{U8D"!S�d    ��O   ��� �<\@��X@��E �&b�|( #�s@ �xi�ZC�"c��T0 k� ��{��{U8D"!S�d    ��O    ��� �<\@��X@��E �%b��|( #�s@ �|g�ZC�!c��T0 k� ��{��{U8D"!S�d    ��O    ��� �8\@��X@��E �$b��|( #�t@ ��f�ZC�c��T0 k� ��{��{U8D"!S�d    ��O    ��� �8\@��X@��E �#b��|( #�t@ ��e�ZC�c��T0 k� ��{��{U8D"!S�d    ��O    ��� �8\@��X@��D �"b��|( #�u@ ��d�ZC�c��T0 k� ��{��{U8D"!S�d    ��O    ��� �8\@��X@��D �!b��|( #�u@ ��b�YC�c��T0 k� ��{��{U8D"!S�d    ��O    ��� �4\@��X@��D � b��|( #�v@ ��a�YC�c��T0 k� ��{��{U8D"!S�d    ��O    ��� �4\@��X@��D � R��|( #�v@ ��`�YS�c��T0 k� ��{��{U8D"!S�d    ��O    ��� �4]@��X@��D �R��|( #�w@ Q�^�YS�c��T0 k� �w{�{{U8D"!S�d    ��O    ��� �4]@��X@��C �R��|( #�w@ Q�]�YS�c��T0 k� �k{�o{U8D"!S�d    ��O    ��� �0]@��X@��C �R��|( #�x@ Q�\�YS�c��T0 k� �c{�g{U8D"!S�d    ��O    ��� �0]@��X@��C �R��|( #�x@ Q�[�XS�c��T0 k� �W{�[{U8D"!S�d    ��O    ��� �0]@��X@��C �R��|( #�y@ Q�Y�XS�c��T0 k� �K{�O{U8D"!S�d    ��O    ��� �0]@��X@��C �R��|( #�y@ Q�X�XS�c��T0 k� �C{�G{U8D"!S�d    ��O    ��� �,]@��X@��B �⣙|( #�z@ Q�W�X3�	c��T0 k� �7{�;{U8D"!S�d    ��O    ��� �,]@��X@��B �⣗|( #�z@ Q�V�X3�c��T0 k� �+{�/{U8D"!S�d    ��O    ��� �,^@��X@��B �⣖|( #�{@ Q�U�X3�c��T0 k� �#{�'{U8D"!S�d    ��O    ��� �,^@��X@��B �⣕|( #�{@ Q�T�X3�c��T0 k� �{�{U8D"!S�d    ��O    ��� �,^@��X@� B �⣓|( #�{@ Q�S�X3�c��T0 k� �{�{U8D"!S�d    ��O    ��� �(^@��X@� B �⣒|( #�|@ a�R�W3�c��T0 k� �{�{U8D"!S�d    ��O    ��� �(^@��X@�A �⣑|( #�|@ a�Q�W3��c��T0 k� ��{��{U8D"!S�d    ��O    ��� �(^@��X@�A �⣐|( #�}@ a�P�W3��c��T0 k� ��{��{U8D"!S�d    ��O    ��� �(^@��X@�A �⟏|( #�}@ a�O�W3��c��T0 k� ��{��{U8D"!S�d    ��O    ��� �(^@��X@�A �⟍|( #�~@ a�N�W3��c��T0 k� ��{��{U8D"!S�d    ��O    ��� �$^@��X@�A �⟌|( #�~@ a�M�W3��c��T0 k� ��{��{U8D"!S�d    ��O    ��� �$_@��X@�A �⛋|( #�~@ a�L�W3��c��T0 k� ��{��{U8D"!S�d    ��O   ��� �$_@��X@�@ ��|( #�@ a�K�W3��c��T0 k� ��{��{U8D"!S�d    ��O    ��� �$_@��X@�@ ��|( #�@ a�J�W3��c��T0 k� ��{��{U8D"!S�d    ��O    ��� �$_@��X@�@ ��|( #�@ a�I�VC��c��T0 k� ��{��{U8D"!S�d    ��O    ��� �$_@��X@�@ ��|( #��@ a�H�VC��c��T0 k� ��{��{U8D"!S�d    ��O    ��� � _@��X@�@ ��|( #�@ a�G�VC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� � _@��X@�@ ��|( #�@ a�F�VC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� � _@��X@�@ ��|( #�@ a�E�VC��c��T0 k� �{|�|U8D"!S�d    ��O    ��� � _@��X@�? ��|( #�@ a�D�VC��c��T0 k� �s|�w|U8D"!S�d    ��O    ��� � _@��X@�? ��|( #�@ a�D�VC��c��T0 k� �g|�k|U8D"!S�d    ��O    ��� � _@��X@�? ��|( #�~@ a�C�VC��c��T0 k� �_|�c|U8D"!S�d    ��O    ��� � `@��X@� ? �R��|( #�~@ a�B�VC��c��T0 k� �S|�W|U8D"!S�d    ��O    ��� �`@��X@� ? �R�|( #�~@ a�A�VC��c��T0 k� �K|�O|U8D"!S�d    ��O    ��� �`@��X@�$? �R{�!�( #�~@ a�@�UC��c��T0 k� �?|�C|U8D"!S�d    ��O    ��� �`@��X@�$? �
Rw�!�( #�~@ a�@�UC��c��T0 k� �7|�;|U8D"!S�d    ��O    ��� �`@��X@�$? �
Rs�!�( �}@ a�?3UC��c��T0 k� �+|�/|U8D"!S�d    ��O    ��� �`@��X@�(> �	Ro�!�( �}@ a�>3UC��c��T0 k� �#|�'|U8D"!S�d    ��O    ��� �`@��X@�(> |	Rk�!�( �}@ a�=3UC��c��T0 k� �|�|U8D"!S�d    ��O    ��� �`@��X@�(> |Bg�!�( �}@ a�=3UC��c��T0 k� �|�|U8D"!S�d    ��O    ��� �`@��X@�,> |Bc�!�( �}@ a�<3UC��c��T0 k� �|�|U8D"!S�d    ��O    ��� �`@��X@�,> |B_�!�( �|@ a�;3UC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �`@��X@�0> |BW�!�( Ӕ|@ a�;3UC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �`@��X@�0> |BS�!�( Ӕ|@ a�:3UC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�0> |BO�!�( Ӕ|@ a�93UC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�4> |BK�|( Ӑ|@ a�9 �UC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�4> |BG�|( Ӑ{@ a�8 �TC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�4= |B?�|( �{@ a�7 �TC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�4= |2;�|( �{@ a�7 �TC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�8= |27�|( �z@ a�6 �TC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�8= |23�|( �z@ a�5 �TC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�8= |2/�|( �z@ b 5 �TC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�<= |2+�|( ��y@ b 4 �TC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�<= |2#�|( ��y@ b4 �TC��c��T0 k� ��|��|U8D"!S�d    ��O    ��� �a@��X@�<= |2�|( ��x@ b3 �TC�c��T0 k� �{|�|U8D"!S�d    ��O    ��� �a@��X@�<= |2�|( �|x@ b3 �TC�c��T0 k� �o|�s|U8D"!S�d    ��O    ��� �a@��X@�@= x2�!�( �|w@ R2 �TC{�c��T0 k� �g|�k|U8D"!S�d    ��O    ��� �a@��X@�@< x2�!�( �xv@ R1 �TC{�c��T0 k� �_|�c|U8D"!S�d    ��O    ��� �a@��X@�@< x2�!�( �xv@ R1 �TC{�c��T0 k� �S|�W|U8D"!S�d    ��O    ��� �b@��X@�D< x "�!�( �tu@ R0 �TCw�d�T0 k� �K|�O|U8D"!S�d    ��O    ��� �b@��X@�D< x "�!�( �tt@ R0 �TCw�d�T0 k� �?|�C|U8D"!S�d    ��O   ��� �b@��X@�D< x "�!�( �ts@ R/ �SCw�d�T0 k� �7|�;|U8D"!S�d    ��O    ��� �b@��X@�D< {�!��!�( �ps@ �/ �SCs�d�T0 k� �/|�3|U8D"!S�d    ��O    ��� �b@��X@�H< {�!��!�( �pr@ �. �SCs�d�T0 k� �#|�'|U8D"!S�d    ��O    ��� �b@��X@�H< {�!��!�( �lq@ �. �SCo�d�T0 k� �|�|U8D"!S�d    ��O    ��� �b@��X@�H< {�!��!�( �lp@ �- �S3o�d�T0 k� �|�|U8D"!S�d    ��O    ��� �b@��X@�H< {�!��!�( �lo@ �, �S3o�d�T0 k� �|�|U8D"!S�d    ��O    ��� �b@��X@�L< {�!�|( �hn@ �+ �S3k�d�T0 k� ��|�|U8D"!S�d    ��O    ��� �b@��X@�L< {�!�|( �hm@ �* �S3k�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �b@��X@�L< {��|( �dl@ �* �S3k�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �b@��X@�L< {��|( �dk@ �) �S3g�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �b@��X@�L; {��|( �dj@ �( �S3g�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �b@��X@�P; {��|( �`h@ �' �S3g�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �b@��X@�P; {��|( �`g@ �% �S3c�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �b@��X@�P; {���|( �`f@ �$ �S3c�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �b@��X@�P; {���|( �\e@ � # �S3_�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �b@��X@�P; {���|( �\d@ � " �S3_�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �b@��X@�T; {���|( �Xb@ � ! �S3[�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �c@��X@�T; {���|( �Xa@ �  �S3[�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �c@��X@�T; {���|( �X`@ �$ �S3W�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �c@��X@�T; {���|( �X^@ �$ �S3S�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �c@��X@�T; {���|( �T]@ �$ �S3S�d�T0 k� �{|�|U8D"!S�d    ��O    ��� �c@��X@�X; {���|( �T\@ �$ �R3O�d�T0 k� �s|�w|U8D"!S�d    ��O    ��� �c@��X@�X; w���|( �TZ@ �( �RCK�d�T0 k� �k|�o|U8D"!S�d    ��O    ��� �c@��X@�X; w���|( �TZ@ �( �RCG�d�T0 k� �_|�c|U8D"!S�d    ��O    ��� �c@��X@�X; w���|( �TY@ �( �RCG�d�T0 k� �W|�[|U8D"!S�d    ��O    ��� �c@��X@�X; w���|( �TW@ �( �RCC�d�T0 k� �O|�S|U8D"!S�d    ��O    ��� �c@��X@�X; w���|( �XV@ �, �RC?�d�T0 k� �G|�K|U8D"!S�d    ��O    ��� �c@��X@�\; w���|( �XU@ �, �QC;�d�T0 k� �;|�?|U8D"!S�d    ��O    ��� �c@��X@�\: w����|( �XT@ �, �QC7�d�T0 k� �3|�7|U8D"!S�d    ��O    ��� �c@��X@�\: w����|( �XS@ �, �QC3�d�T0 k� �+|�/|U8D"!S�d    ��O    ��� �c@��X@�\: w����|( �XR@ �0 �QC/�d�T0 k� �#|�'|U8D"!S�d    ��O    ��� �c@��X@�\: w����|( �XP@ �0
 �PC+�d�T0 k� �|�|U8D"!S�d    ��O    ��� �c@��X@�\: w���|( �XO@ �0 �PC'�d�T0 k� �|�|U8D"!S�d    ��O    ��� �c@��X@�`: w���|( �XN@ �0 �PS#�d�T0 k� �|�|U8D"!S�d    ��O    ��� �c@��X@�`: w���|( �XL@ �0 �PS�d�T0 k� ��|�|U8D"!S�d    ��O    ��� �c@��X@�`: w���|( �XK@ �4 �PS�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �c@��X@�`: w���|( �XI@ �4  �PS�d�T0 k� ��|��|U8D"!S�d    ��O   ��� �c@��X@�`: w���|( �\H@ �7� �OS�d�T0 k� ��|��|U8D"!S�d    ��O    ��� �c@��X@�`: w���|( �\G@ �7� �O	��d�T0 k� ��|��|U8D"!S�d    ��O    ��� �c@��X@�`: w���|( �\E@ �7� �O	��d�T0 k� ��|��|U8D"!S�d    ��O    ��� �c@��X@�d: w���|( �\D@ ;� �O	��d�T0 k� ��|��|U8D"!S�d    ��O    ��� �c@��X@�d: w��#�|( �\B@ ;� �O	��d�T0 k� ��|��|U8D"!S�d    ��O   ��� �c@��X@�d: w��'�|( �\A@ ;� �N	���d�T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�d: w��+�|( �\?@ ?� �N	���d�T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�d: w��3�|( �\=@ ?� � N	���d�T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�d: w��7�|( �\<@ C� � N	���d�T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�d: w��;�|( �\:@ C� � N	��d�T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�h: w��?�|( �\9@ G� � N	��d�T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�h: w��G�|( �\7@ �G� ��M	��"��T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�h: w��K�|( �\5@ �K� ��M	��"��T0 k� �{|�|U8D"!S�d    ��O    ��� �d@��X@�h: w��O�|( �\3@ �O� ��M	��"��T0 k� �s|�w|U8D"!S�d    ��O    ��� �d@��X@�h: w��W�|( �`2@ �O� ��M	��"��T0 k� �k|�o|U8D"!S�d    ��O    ��� �d@��X@�h: w��[�|( �`0@ �S� ��M	��"��T0 k� �_|�c|U8D"!S�d    ��O    ��� �d@��X@�h: w��c�|( �`.@ �W� ��M	��"��T0 k� �W|�[|U8D"!S�d    ��O    ��� �d@��X@�h9 w��g�|( �`,@ �W� ��M	��"��T0 k� �O|�S|U8D"!S�d    ��O   ��� �d@��X@�h9 w��o�|( �`+@ �[� ��L	��"��T0 k� �G|�K|U8D"!S�d    ��O    ��� �d@��X@�l9 w��w�|( �`)@ �_� ��L	��"��T0 k� �?|�C|U8D"!S�d    ��O    ��� �d@��X@�l9 w���|( �`'@ �c� ��L	��"��T0 k� �7|�;|U8D"!S�d    ��O    ��� �d@��X@�l9 w���|( �`%@ �c� ��L	��"��T0 k� �/|�3|U8D"!S�d    ��O    ��� �d@��X@�l9 w���|( �`$@ �c� ��L	��d�T0 k� �#|�'|U8D"!S�d    ��O    ��� �d@��X@�l9 w���|( �`"@ �c� ��L	��d�T0 k� �|�|U8D"!S�d    ��O    ��� �d@��X@�l9 w����|( �` @ �g� ��L	��d�T0 k� �|�|U8D"!S�d    ��O    ��� �d@��X@�l9 w����|( �`@ �k� ��K	��d�T0 k� �|�|U8D"!S�d    ��O    ��� �d@��X@�l9 w����|( �`@ �k� ��K	��d�T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�p9 w����|( �`@ �o� ��K	��d�T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�p9 w����|( �`@ �s� ��K	��d�T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�p9 w����|( �`@ �s� ��K	��d�T0 k� ��|��|U8D"!S�d    ��O    ��� �d@��X@�p9 w����|( �d@ �w� ��K	��d�T0 k� ��|��|U8D"!S�d    ��O    ��� � d@��X@�p9 w����|( �d@ �{� ��K��d�T0 k� ��|��|U8D"!S�d    ��O    ��� � d@��X@�p9 w���|( �d@ �� ��K��"��T0 k� ��|��|U8D"!S�d    ��O    ��� � d@��X@�p9 w���|( �d@ �� ��K��"��T0 k� ��|��|U8D"!S�d    ��O   ��� � d@��X@�p9 w���|( �d@ � ��J��"��T0 k� ��|��|U8D"!S�d    ��O    ��� � d@��X@�p9 w��'�|( �d@ � ��J��"��T0 k� ��|��|U8D"!S�d    ��O    ��� � d@��X@�p9 w��/�|( �d	@ � ��JR�"��T0 k� ��|��|U8D"!S�d    ��O    ��� � d@��X@�p9 w��;�|( cd@ � ��JR�"��T0 k� ��|��|U8D"!S�d    ��O    ��� � d@��X@�t9 w��C�|( cd@ 	� ��JR�"��T0 k� ��|��|U8D"!S�d    ��O    ��� � e@��X@�t9 w��K�|( cd@ 	� ��JR�"��T0 k� ��|��|U8D"!S�d    ��O    ��� � e@��X@�t9 w��S�|( cd@ 	� ��JR�"��T0 k� ��|��|U8D"!S�d    ��O    ��� � e@��X@�t9 w��[�|( cd @ 	� ��JR�"��T0 k� �|��|U8D"!S�d    ��O    ��� � e@��X@�t9 w��c�|( cg�@ 	� ��JR�"��T0 k� �w|�{|U8D"!S�d    ��O    ��� � e@��X@�t9 w��k�|( cc�@ 
�� ��JR�d�T0 k� �o|�s|U8D"!S�d    ��O    ��� � e@��X@�t9 w��s�|( cc�@ 
�� ��IR�d�T0 k� �g|�k|U8D"!S�d    ��O    ��� � e@��X@�t9 w��{�|( 3c�@ 
�� ��IR�d�T0 k� �_|�c|U8D"!S�d    ��O    ��� � e@��X@�t9 w����|( 3c�@ 
�� ��IR�d�T0 k� �W|�[|U8D"!S�d    ��O    ��� � e@��X@�t9 w����|( 3c�@ 
�� ��IR�d�T0 k� �O|�S|U8D"!S�d    ��O    ��� � e@��X@�t9 w� c��|( 3c�@ 	� ��IR�d�T0 k� �G}�K}U8D"!S�d    ��O    ��� � e@��X@�t9 s� c��|( 3_�@ 	� ��IR�d�T0 k� �?}�C}U8D"!S�d    ��O    ��� � e@��X@�t9 s� c��|( 3_�@ 	� ��IR�d�T0 k� �;}�?}U8D"!S�d    ��O    ��� � e@��X@�t9 s� c��|( 3_�@ 	� ��IR�d�T0 k� �3~�7~U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( 3_�@ 	� ��IR�d�T0 k� �+~�/~U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( 3_�@ 
�� ��IR�d�T0 k� �#�'U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( 3_�@ 
�� ��IR�d�T0 k� ��#U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( 3_�@ 
�� ��IR�d�T0 k� ����U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( 3[�@ 
�� ��IR�d�T0 k� ����U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( 3[�@ 
�� ��HR�d�T0 k� ����U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( 3[�@ r�� ��HR�d�T0 k� ����U8D"!S�d    ��O   ��� � e@��X@�x9 s� c��|( C[�@ r�� ��HR�d�T0 k� �����U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( C[�@ r�� ��HR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( C[�@ r�� ��HR�d�T0 k� �����U8D"!S�d     �O    ��� � e@��X@�x9 s� c��|( C[�@ r�� ��HR�d�T0 k� ����U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( CW�@ r����HR�d�T0 k� ����U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( CW�@ r����HR�d�T0 k� ����U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( CW�@ r����HR�d�T0 k� �߇��U8D"!S�d    ��O   ��� � e@��X@�x9 s� c��|( CW�@ r����HR�d�T0 k� �ۇ�߇U8D"!S�d    ��O    ��� � e@��X@�x9 s� c��|( CW�@ r����HR�d�T0 k� �ӈ�׈U8D"!S�d    ��O    ��� � e@��X@�|9 s� c��|( CW�@ r����HR�d�T0 k� �ω�ӉU8D"!S�d    ��O    ��� � e@��X@�|9 s� c��|( CW�@ �����HR�d�T0 k� �ˊ�ϊU8D"!S�d    ��O    ��� � e@��X@�|9 s� c��|( CW�@ �����HR�d�T0 k� �ǋ�ˋU8D"!S�d    ��O    ��� � e@��X@�|9 s� c��|( CS�@ �����HR�d�T0 k� �Ì�ǌU8D"!S�d    ��O    ��� � e@��X@�|9 s� c��|( CS�@ �����HR�d�T0 k� ����ÍU8D"!S�d    ��O    ��� � e@��X@�|9 s� c��|( CS�@ �����GR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|9 s� c� |( CS�@ �����GR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|9 s� c�|( CS�@ �����GR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|9 s� c�|( CS�@ �����GR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�|( CS�@ �����GR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�|( CS�@ �����GR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�|( CS�@ �����GR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�|( CS�@ �����GR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�|( CO�@ �����GR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�|( CO�@ �����GR�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�|( CO�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�	|( CO�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�
|( CO�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�
|( CO�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@�|8 s� c�|( CO�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CO�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CO�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CO�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CO�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CO�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CK�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CK�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CK�@ �����G�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CK�@ �����F�d�T0 k� ������U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CK�@ �����F"�d�T0 k� �����U8D"!S�d    ��O   ��� � e@��X@��8 s� c�|( CK�@ �����F"�d�T0 k� �����U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( CK�@ �����F"�d�T0 k� �����U8D"!S�d    ��O    ��� � e@��X@��8 s� c�|( 3K�@ �����F"�d�T0 k� �{���U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( 3K�@ �����F"�d�T0 k� �{���U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( 3K�@ �����F"�d�T0 k� �{���U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( 3K�@ �����F"�d�T0 k� �w��{�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( 3K�@ �����F"�d�T0 k� �w��{�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( 3K�@ �����F"�d�T0 k� �w��{�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( 3K�@ �����F"�d�T0 k� �w��{�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( 3G�@ �����F"�d�T0 k� �s��w�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( 3G�@ �����F"�d�T0 k� �s��w�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( 3G�@ �����F"�d�T0 k� �s��w�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( 3G�@ r����F"�d�T0 k� �s��w�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( cG�@ r����F"�d�T0 k� �s��w�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( cC�@ r����F"�d�T0 k� �o��s�U8D"!S�d    ��O   ��� � f@��X@��8 s� c�|( cC�@ r����F"�d�T0 k� �o��s�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( cC�@ r����F"�d�T0 k� �o��s�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( c?�@ r����F"�d�T0 k� �o��s�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( S?�@ r����F"�d�T0 k� �o��s�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( S?�@ r����F"�d�T0 k� �o��s�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( S;�@ r����F"�d�T0 k� �o��s�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( S;�@ r����F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( S7�@ r����F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( �3�@ r����F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�|( �3�@ B����F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c� |( �/�@ B����F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c� |( �+�@ B�� ��F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�!|( �+�@ B�� ��F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�!|( �'�@ B�� ��F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�"|( �#�@ B�� ��F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�"|( �#�@ B�� ��F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�"|( �#�@ B�� ��F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�#|( �#�@ B�� ��F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�#|( �#�@ B�� ��F"�d�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�$|( �#�@ B�� ��F"�d#�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�$|( �#�@ B�� ��F"�d#�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�$|( �#�@ B�� ��F"�d#�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�%|( �#�@ B�� ��F"�d#�T0 k� �k��o�U8D"!S�d    ��O    ��� � f@��X@��8 s� c�%|( S#�@ B�� ��F"�d#�T0 k� �k��o�U8D"!S�d    ��O   ��� � ��eASK�@;�X`h �\A���A��u�D@׏ ��"s� T0 k� �K��O�U8D"!�cU2d   ��O    � �N ��eASK�@;�X`h �]A���A��u�E@א ��"s� T0 k� �3��7�U8D"!�cU2d   ��O    � �L ��eASK�@;�X`h �]A���A��u�E@א ��"s� T0 k� ����U8D"!�cU2d   ��O    � �J ��eASK�@;�X`h �]A���A��u�E@א ��3� T0 k� ����U8D"!�cU2d   ��O    � �H ��fASK�@;�X`h �^A���A��u�F@א ��3� T0 k� ������U8D"!�cU2d   ��O    � 
�G ��fASK�@;�X`d �^A���A��t�F@א ��3� T0 k� ������U8D"!�cU2d   ��O    � 	�F ��fASK�@;�X`d �^A���A��t�G@א ��3� T0 k� ������U8D"!�cU2d   ��O    � �E ��fASK�@;�\ad  �^A���A��t�G@Ӑ ��3� T0 k� ������U8D"!�cU2d   ��O    � �D��A��P"��B� s�| �c�@ Sw� �c���c� T0 k� �;��?�U8D"!S�d    ��/   ��� ��A��P"��B� s�!� �c�@ Sw� �c���"�� T0 k� �;��?�U8D"!S�d    /�/   ��� ���A��P"��B� s�!� �c�@ Sw� �c���"�� T0 k� ����U8D"!S�d    ��/   ��� ���A��P��B� s�!� �c�@ �s� �c���"���T0 k� ����U8D"!S�d    $�/   ��� ���A��P�� � s�!� �c�@ �s� �c���"���T0 k� 3���U8D"!S�d    ��/   ��� ���A��P�� � s�!� �c�@ �s� �c���"���T0 k� 3���U8D"!S�d    ��/   ��� ���A��P�� � s�!�  �c�@ �k� �c���"���T0 k� 3���U8D"!S�d    ��/   ��� ���A��P�� � s�!�  �c�@ �c� �c���"���T0 k� 3���U8D"!S�d    ��/   ��� � �D��P�� � bs�!�$ Cc�@ �[�c����"���T0 k� 3���U8D"!S�d    ��/   ��� � �D��P"�� b� bs�|$ Cc�@ �S�c����c��T0 k� ����U8D"!S�d    ��/   ��� � �D��P"�� b� bs�|$ Cc�@ �K�c����c��T0 k� ����U8D"!S�d    ��/   ��� � �D��P"�� b� bs�|( Cc�@ �C�_����c��T0 k� ����U8D"!S�d    ��/   ��� � �D��P"�� b� bs�|( Cc�@ �C�_����c��T0 k� ����U8D"!S�d    ��/   ��� � c�D��P"�� b� �s�|(  c�@ �C��_���c��T0 k� ����U8D"!S�d    $�/   ���  c�D��P"�� �� �s�|(  c�@ �?��_���c��T0 k� 3���U8D"!S�d    ��/   ���  c�D��P"�� �� �s�|(  c�@ �;��_���c��T0 k� 3��#�U8D"!S�d    ��/   ���  c�D��P"� �� �s�|(  c�@ �;��_���c��T0 k� 3��#�U8D"!S�d    ��/   ���  c�D��P"� �� �s�|(  c�@ �7��[���c��T0 k� 3#��'�U8D"!S�d    ��/   ��� C�D��P� ��s�|(  �_�@ �3�C[���c��T0 k� 3#��'�U8D"!S�d    ��/   ��� C�D��P��s�|(  �_�@ �3�C[���c��T0 k� �'��+�U8D"!S�d    ��/   ��� C�D��P��s�!�(  �_�@ �/�C[���"���T0 k� �'��+�U8D"!S�d    ��/   ��� C�D��P��s�!�(  �_�@ �+�C[���"���T0 k� �+��/�U8D"!S�d    ��/   ��� �C�D��P��s�!�(  �_�@ �+�C[���"���T0 k� �/��3�U8D"!S�d    ��"   ��� �C�D��@b��Rs�!�( _�@ �'�CW���"���T0 k� �#��'�U8D"!S�d    ��"   ��� �C�D��@b߹�Rs�!�( [�@ �#�CW���"���T0 k� ����U8D"!S�d    ��"   ��� �C�D��@b۹R�Rs�!�( [�@ �#�CW���"���T0 k� ����U8D"!S�d    ��"   ��� �C�D��@b۹R�Rs�!�( [�@ ��CW���"���T0 k� ����U8D"!S�d    ��"   ��� �C�D��@�׹R�Ro�!�( �W�@ ��SW���"���T0 k� �����U8D"!S�d    ��"   ��� �S�D��@�ӹR��o�!�( �S�@ ��SS���"���T0 k� ����U8D"!S�d    ��"   ��� �S�D��@�ӹ���o�!�( �O�@ ��SS���"���T0 k� �۪�ߪU8D"!S�d    ��"   ��� �S�D��@�ӹ���k�|( �O�@ ��SS���c��T0 k� �ө�שU8D"!S�d    ��"   ��� �S�D��@�Ϲ���k�|( �O�@ C�SS���c��T0 k� �˨�ϨU8D"!S�d    ��"   ��� �S�E��@�Ϲ���g�|( SK�@ C�3S���c��T0 k� �Ǩ�˨U8D"!S�d    ��"   ��� �S�E��@�˹���g�|( SG�@ C�3S���c��T0 k� �è�ǨU8D"!S�d    ��"   ��� �S�E��@�˹���c�|( SG�@ C�3S���c��T0 k� ����èU8D"!S�d    ��"   ��� �S�E��E2˹����_�|( SC�@ C�3O���c��T0 k� ����çU8D"!S�d    ��"   ��� �S�E��E2ǹ����_�|( S?�@ C�3O���c��T0 k� ������U8D"!S�d    ��"   ��� �S�E��E2ǹ����W�|( C;�@ C�#O�%�{�c��T0 k� ������U8D"!S�d    ��"   ��� �c�E��E2ù����S�|( C7�@ C�#O�%�{�c��T0 k� ������U8D"!S�d    ��"   ��� �c�F�E"ø����S�|( C3�@ ��#S�%�w�c��T0 k� �è�ǨU8D"!S�d    �"   ��� �c F�E"ø����O�|( C/�@ ��#S�%�s�c��T0 k� �ϫ�ӫU8D"!S�d    ��/   ��� �cF�E"øA���K�|( C+�@ ��#S�%�o�c��T0 k� �׮�ۮU8D"!S�d    ��/   ��� �	SF�E"��A���C�|( 3#�@ ���#S�%�k�c��T0 k� ����U8D"!S�d    ��/   ��� �	SF�F���A���?�|( 3#�@ ���#W�%�g�c��T0 k� ������U8D"!S�d    ��/   ��� �	SF�F���A��;�|( 3�@ ���#W�%�c�c��T0 k� ����U8D"!S�d    ��/   ��� �	SF�F���A��3�|( 3�@ ���#W�%�_�c��T0 k� ����U8D"!S�d    ��/   ��� �	S	F�F���A��/�|( 3�@ ���#[�%�_�c��T0 k� ����U8D"!S�d    ��/   ��� �	c
F�F���1��+�|( 3�@ ����[�%�[�c��T0 k� ���#�U8D"!S�d    ��/   ��� �	cF�F���1��B#�|( 3�@ ����_�%�W�c��T0 k� �;��?�U8D"!S�d    ��   ��� �	cE��F���1��B�|( 3�@ ����_�%�S�c��T0 k� �7��;�U8D"!S�d    ��   ��� �	cE��F���1��B�|( �@ ����c�%�S�c��T0 k� �7��;�U8D"!S�d    ��   ��� �#E��F���A��B�|( �@ ���	3c�%�S�c��T0 k� �;��?�U8D"!S�d    ��   ��� �#E��F���A��B�|( �@ ���	3g�%�K�c��T0 k� �;��?�U8D"!S�d    ��   ��� �#Es#�F���A����|( �@ ���	3g�%�K�c��T0 k� �;��?�U8D"!S�d    ��   ��� �#Es#�F���A�����|( ��@ ���	3g�%�G�c��T0 k� �7��;�U8D"!S�d    ��   ��� �#Es'�F���A�����|( ���@ ҿ�	Cg�%�G�c��T0 k� �7��;�U8D"!S�d    ��   ��� �#Es'�F���A���|( ���@ ҷ�	Cg�%�?�c��T0 k� �7��;�U8D"!S�d    ��   ��� �#B+�F���A�A�|( ���@ ү�	Cg�%�?�c��T0 k� �3��7�U8D"!S�d    ��   ��� ��B+�F���A�A�|( B��@ ҫ�	Cg�%�;�c��T0 k� �3��7�U8D"!S�d    ��   ��� ��B+�F���Q�Aۮ|( B��@ ң�	3g�%�;�c��T0 k� �/��3�U8D"!S�d    ��   ��� ��B/�F���Q�Aׯ|( B��@ ҟ�	3g�%�7�c��T0 k� �+��/�U8D"!S�d    ��   ��� ��B/�F���Q�	A˰|( B��@ ҏ�	3g�%�3�c��T0 k� �+��/�U8D"!S�d    ��   ��� ��F3�F���Q�Añ|( B��@ ҋ�	3g�S3�c��T0 k� �;��?�U8D"!S�d    ��   ��� ��  F3�F���Q�A��|( 2��@ ��	Cg�S/�c��T0 k� �G��K�U8D"!S�d    ��   ��� ��$!F3�F���Q�1��|( 2��@ �{�	Cg�S+�c��T0 k� �O��S�U8D"!S�d    ��   ��� �$"F7�F���Q�1��|( 2��@ �s�	Cg�S'�c��T0 k� �W��[�U8D"!S�d    ��   ��� �,%F;�F���Q�1��|( 2��@ �g�	Cg�S#�c��T0 k� �_��c�U8D"!S�d    ��   ��� �0'F?�F���Q�1��|( 2��@ 2_�	3g�C�c��T0 k� �g��k�U8D"!S�d    ��   ��� 0(F?�@b��a�1��|( 2��@ 2W�	3g�C�c��T0 k� �k��o�U8D"!S�d    ��   ��� 4*FC�@b��a�1��|( 2��@ 2O�	3g�C�c��T0 k� �o��s�U8D"!S�d    ��   ��� <-FG�@b��a�1��|( 2��@ 2C�	3g�C�c��T0 k� �s��w�U8D"!S�d    ��   ��� @.BSK�@b��a�A��|( "��@ R;�	Cg�C�c��T0 k� �s��w�U8D"!S�d    ��   ��� D0BSO�E��a�A{�|( "��@ R3�	Cg�C�c��T0 k� �s��w�U8D"!S�d    ��   ��� H1BSS�E��a� Aw�|( "��@ R+�	Cg�C�c��T0 k� �s��w�U8D"!S�d    ��   ��� L3BSW�E��a�"As�|( "��@ R#�	Cg�C�c��T0 k� �s��w�U8D"!S�d    ��   ��� P5BSW�E��a�$Ak�|( "� @ R�	Cg�B��3��T0 k� �s��w�U8D"!S�d    ��   ��� X8Es_�E��a|(1c�|( "�@ R�	3g�B��3��T0 k� �p�tU8D"!S�d    ��   ��� \:Esc�E���qx*1_�|( "�@ ���	3g�B��3��T0 k� �p�tU8D"!S�d    ��   ��� `;Esg�E���qx,1W�|( �@ ���	3g�B��3��T0 k� �t
�x
U8D"!S�d    ��   ��� d=Esg�E���qt.1S�|( �@ ���	3g�B��3��T0 k� �t�xU8D"!S�d    ��   ��� l?Esk�E���qt01O�|( �@ ���	3g�B��3��T0 k� �x�|U8D"!S�d    ��   ��� p@Eso�E���qp21K�|( �@ ��� �g�B��3��T0 k� �|��U8D"!S�d    ��   ��� #tBEsp E���	Qp41G�|( �@ ��� �g�B��3� T0 k� ����U8D"!S�d    ��   ��� #�FBtEr��	Ql71;�|( ��	@ ��� �g�B��3�T0 k� �|��U8D"!S�d    ��   ��� #�HBxEr��	Ql917�|( ��
@ �� �g�2��3�T0 k� �|��U8D"!S�d    ��   ��� #�IBxEr��	Ql;!3�|( ��@ �� �g�2��3�T0 k� �|��U8D"!S�d    ��   ��� #�KB|
Er��	al<!/�|( ��@ Q��g�2��3�T0 k� �x�|U8D"!S�d    ��   ��� #�MB�Er��	ah>!+�|( ��@ Q��g�2��3�T0 k� �| �� U8D"!S�d    ��   ��� #�OEs�Er��	ah@!'�|( ��@ Q��g�2���T0 k� ��#��#U8D"!S�d    ��   ��� �REs�Er��	ahB!#�|( ��@ Q��g�2���	T0 k� ��(��(U8D"!S�d    ��   ��� �TEs�D���	QhD!�|( ��@ Q���g�B���
T0 k� ��+��+U8D"!S�d    �   ��� �VEs�D���	QhE!�|( ��@ Q{��g�B���
T0 k� ��.��.U8D"!S�d    �� 
  ��� �WH��D���	QhG!�|( ��@ Qs��c�B���T0 k� ��2��2U8D"!S�d    �� 
  ��� �YH��D���	QhH!�|( ��@ Qk��c�B���T0 k� ��5��5U8D"!S�d    �� 
  ��� C�[H��D���	QhJ!�|( ��@ Q_��c�B���T0 k� ��8��8U8D"!S�d   �� 
  ��� C�^H��!D���1hM�|( ��@ QO��_�2���T0 k� ��>��>U8D"!S�d   ��? 
  ��� C�`H��#D���1hN�|( ��@ AO��_�2����T0 k� ��A��AU8D"!S�d   ��? 
  ��� C�bH��%D�ö1hP�|( ��@ AK��[�2����T0 k� ��D��DU8D"!S�d   ��? 
  ��� C�cH��'D�÷1hR�|( ��@ AG��[�2����T0 k� ��G��GU8D"!S�d   ��? 
  ��� C�eH��)D�Ƿ1hT��|( ��@ AC��W�2����T0 k� ��J��JU8D"!S�d   ��? 
  ��� C�gH��+D�Ǹ�dU��|( ��@ A?��W�"����T0 k� ��M��MU8D"!S�d   ��? 
  ��� C�hH��,D�ǹ�dW��|( ��@ A7��S�"� ��T0 k� ��P��PU8D"!S�d   ��? 
  ��� C�lH��0D�˻�dZ��|( ��@ A7�3O�"���T0 k� ��V��VU8D"!S�d   ��?   ��� C�mH��2D�˼�d\��|( ��@ A3�3O�"���T0 k� ��Y� YU8D"!S�d    ��?   �  D oH��3D�˽�d^��|( ��@ A/�3K�����T0 k� �\�\U8D"!S�d    ��?   �  DqH��5D�Ͽ�d`��|( ��@ A+�3K�����T0 k� �_�_U8D"!S�d    ��?   �  DsH��7D����`b���|( ��@ A'�3G�����T0 k� �b�bU8D"!S�d    ��?   � 
 DtH��8D����`d���|( ��@ 1#�3G�����!T0 k� �e�eU8D"!S�d    ��?   �  DvH��:D����`e���|( ��@ 1�3C���	��"T0 k� � h�$hU8D"!S�d    /�?   �  DwH��;D����\g���|( ��@ 1�CC�����$T0 k� �$k�(kU8D"!S�d    ��?   �  D yH��=D����\i���|( �� @ 1�C?�����&T0 k� �,n�0nU8D"!S�d    ��?   �  D xH��@D����Xm���|( �"@ 1�C;�����*T0 k� �<t�@tU8D"!S�d    �?   �  D wH��BD����To���|( �#@ � C;����,T0 k� �Hp�LpU8D"!S�d   ��?   �  D wH��CD����Tq���|( �$@ � �7����.T0 k� �Xk�\kU8D"!S�d   ��?   �  D vH��DD����Pr���|( �%@ ���7����/T0 k� �hg�lgU8D"!S�d   ��?   �  4vH��FD����Lt���|( �&@ ���3����1T0 k� �tc�xcU8D"!S�d   ��?   �  4uH��GD����Lv���|( �'@ ���/����2T0 k� �|^��^U8D"!S�d   ��?   �  4uH��ID����Hw���|( � (@ 0��/����3T0 k� ��Y��YU8D"!S�d   ��?   �  4tH��JD����Dy���|( �$)@ 0�
�+����4T0 k� ��T��TU8D"!S�d   ��?   �   4tH��KD����@{���|( (*@ 0��'����5T0 k� ��O��OU8D"!S�d   ��?   � ! $sI��MD����<|���|( ,+@ 0�C'��3�7T0 k� ��J��JU8D"!S�d   ��?   � " $sI��NI����8~���|( 0,@ 0�C#��3�8T0 k� ��E��EU8D"!S�d   ��?   � " $rI��OI����8����|( 8-@ 0�C��3�9T0 k� ��@��@U8D"!S�d   ��?   � " $rI��PI����4���|( <.@ 0�C�� 3�:T0 k� ��<��<U8D"!S�d   ��?   � " $qI��QI����0���|( �@/@ 0�C��!3�:T0 k� ��7��7U8D"!S�d   ��?   � " $qI��RI����,~���|( �D1@ 0�3��#��;T0 k� ��2��2U8D"!S�d   ��?   � " $pI��SI����(~���|( �L2@ 0�3��$��<T0 k� ��-��-U8D"!S�d   ��?   � " $pI��TI���1 }���|( �P3@ @�3��&��<T0 k� ��(��(U8D"!S�d   ��?   � " $oI��VI���1|���|( �X5@ @�3�"�)��=T0 k� ����U8D"!S�d    ��?   � " $oI��WI���1|���|( �`6@ @� C�"�+��=T0 k� ����U8D"!S�d    ��?   � " $nI��WI���1{���|( �d7@ @�"C�"�,��>T0 k� ����U8D"!S�d    .�?   � " $nI��XE���Q{���|( �h9@ 0�$C�# . �>T0 k� ����U8D"!S�d    ��?   � " $mI��YE���Q{���|( �p:@ 0�&C�#0 �>T0 k� ����U8D"!S�d    �?   � " $mI��YE���Q z���|( �t;@ 0�'C�#1 �>T0 k� ����U8D"!S�d    ��?   � " $mI��ZE���P�z���|( �x<@ 0�)��3 �>T0 k� ����U8D"!S�d    ��?   � " $lI��ZE���P�y���|( �=@ 0�+��5 �=T0 k� ������U8D"!S�d    ��?   � " $lI��[O���P�y���|( �>@ 0�-�6 �=T0 k� ������U8D"!S�d    ��?   � ! $kI��[O���P�x���|( �@@  �/�8 �=T0 k� ������U8D"!S�d    ��?   �   $kI��\O�����x���|( �A@  �1�9 �<T0 k� ������U8D"!S�d    ��?   �  $kI��\O�����x���|( �B@  �3�	 ; �<T0 k� ������U8D"!S�d    ��?   �   jI��\O�����w���|( �B@  �5�
	$< �;T0 k� ������U8D"!S�d    ��?   �   jI��]O�����v���|( �D@  �9�	(? �9T0 k� ������U8D"!S�d    ��?   �   iI��]O�����v���|( ��D@  �<�	,@ �8T0 k� ������U8D"!S�d    ��?   �    iI��]O�����v���|( ��E@  �>�	#,A �7T0 k� ������U8D"!S�d    ��?   �  � iI��]O�� �u���|( ��F@  �@�	#0B �6T0 k� ������U8D"!S�d    ��?   �  � hI��]O���u���|( ��G@  �B�	#4C �5T0 k� ������U8D"!S�d    ��?   �  �$hI��]O���t���|( ��H@  �D�	#4D �4T0 k� ������U8D"!S�d    ��?   �  �$hI��]O���t���|( ��I@  �F�	#8F��3T0 k� ������U8D"!S�d    ��?   �  �(gI��]O����s��|( ��J@ �H�<G��1T0 k� ������U8D"!S�d    ��?   � 	 �(gBC�]O����s��|( ��K@ �J�@H��0T0 k� ������U8D"!S�d    ��?   �  �,gBC�]O��
��r��|( ��L@ �L� DI��/T0 k� ������U8D"!S�d    ��   �  �,fBC�]O� ��r��|( ��M@ �N�"HJ��-T0 k� ������U8D"!S�d    ��   �   �0fBC�]O� ��q��|( ��M@ �P�#LK��,T0 k� ������U8D"!S�d    ��   ��� �4fBC�^O� �xq��|( ��N@ �R�%PL��*T0 k� ������U8D"!S�d    ��   ��� �8eE��_O��lo��|( ��N@ �V�(�XN��'T0 k� �����U8D"!S�d    ��   ��� �<eE��_O��dn�'�|( ��N@ �X�*�\N��%T0 k� �w��{�U8D"!S�d    ��   ��� �@eE��`O��\n�+�|( ��O@ �Z�,�dO��#T0 k� �o��s�U8D"!S�d    ��   ��� �DdE��`F�Tm�/�|( ��O@ �\�-�hP��!T0 k� �g��k�U8D"!S�d    ��   ��� �HdE��`F�Ll�3�|( ��P@ �]�/�lQ��T0 k� �[��_�U8D"!S�d    ��   ��� �LdE��`F�Dk;�|( ��P@ ��_�1�pQ��T0 k� �S��W�U8D"!S�d    ��   ��� ��PdE��aF�@j?�|( ��Q@ ��a�2�tR��T0 k� �G��K�U8D"!S�d    ��   ��� ��TcE��aF�8jC�|( ��Q@ ��b�4�|R��T0 k� �;��?�U8D"!S�d    ��   ��� ��`cE��aF�(hO�|( ��Q@ ��e�7��S��T0 k� �#��'�U8D"!S�d    ��   ��� �	`bA�aF � gS�|( ��Q@ ��g�8��T��T0 k� ����U8D"!S�d    ��   ��� �                                                                                                                                                                            � � �  �  �  c A�  �J����  �      � \��m ]�+D+D � � f"�    �      � '     f"� '                       ~           �@     ���   (

          X]   9     � ���     X] ���           
             
 	 ] �         ��      ���   8�           8�-          !��     8�-!�       a   	            �         �      ���   	@
		          ���    5	     ���    ��_���    ��                    ��           �      ���   H	$
          %��          . �2^     %zK �*D    D z               ���          X       ���   H
	!           �5  �  	    B�
�      �5�
�                         	   �p���C         ��      ���      0            ��,�  U U      V �0�    ���p șY    ���#            C�� �         @b     ��@ 
@				         �
       j  2�    �
  2�               ��      � !�        p       ��F  0	%          ����  $ $     ~ ��@    ���� ��.      ��          A	�� ��        0       ��@   0
 
          FZ      � �O�     F# �V�    ����             0 �� �         	 p     ��H   8         ��͸  � �
	   � �U�    ���- ��>     ���            :	�� �         
 ��     ��`   P
	
         ���r ��
	      ��    ����
�    �� .                     ���c        �   �  ��@    P                   ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��d�  ��        ����    �������    |                  x        �       j  �   �   �                         ��    ��        ���      ��  ��           "                                                �                           �!�� ��
 �   � � �������  
     	          
  P   �	� ��C       = �j� >  k� �D  r� �� s  �� 0s@ �  s� �D s����X � �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā���� � �� �R� 
�\ U� 
�� V  
�| V ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���� � �����R  ������  
�fD
��L���"����D" � j  "  B   J jF�"    "�j * , ����
��"     �j @�    �
� �  �  
�      ��     � �  �    %    ��     � �       F��  ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �O�!      ��t �  ���        �t �  ��        �        ��        �        ��        �      �     [������        ��                         �7Y 	 � ���                                     �                ����               ����%��  �� � 2�� � $          �EDM 51%) derson y   0:00                                                                        2  2     � �
�b �c~ � � c� � �c� � c�� �c� � � c� � � c� � � 	c� � � 
c� � � c� � �cV � �c^ � �C.Z �C6j �
c� � c�	 | c�	 {	�$ {	�; ��" ��M eKg } K_ �"�U � "�g �"�Q �*�` �"�r � "�� ��r � 
��+!� � �"� � �#� � �$": � � %"P � �&!� � �'"* | �("< � �)"2 | *"@ |& +"P �N ,"& |^  "* |^  "  |& /"J �^  "  |N 1"& |^  "* | � 3"A � 4"P �$  " ~)  " { � 7*O~ � 8*K~  )�~ � :*K~  )�~ �<*$X �=* p � >"K x  !� p                                                                                                                                                                                                                         �� P             @ �      ( 	�     [ P E a  ��        	            	�������������������������������������� ���������	�
��������                                                                                          ��    �tM�� ��������������������������������������������������������   �4, F�  @�7������                                                                                                                                                                                                                                                                                                                                                       �R �#�                                                                                                                                                                                                                                         
     
  	  )      	  H�J     9i                             ������������������������������������������������������                                                                                                                                    
      �             �        �    �   o          
 	  
	 
 	 	 ������������ ����� ��������������������������� ������������������� �����  ������� ������������������������� �����  �������������������� �� � ����������������������� � ������������������������������������������������������� �����������             	                  �    /    � �  D�J    	  �=  	                           ������������������������������������������������������                                                                        
                                                                  �     |      �   	    |        �  �          	  
 	 
 	 	 ������ �������������� ��� ���������������� ��������������  � �������������������������� � ���� ����� ����������� � �������������������� �������� �������  ����������� ������� ������������������������������ �������   ����� �  ���             o                                                                                                                                                                                                                                                                                                     
          �             


           �   }�         wwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwww % K ?                	                 � ��o �j�                                                                                                                                                                                                                                                                                     
)n1n  !Y                    b            m                  f                                                                                                                                                                                                                                                                                                                                                                                                        P L  � ��  � ��  � (��  � #��  CfL  �ɬ������������r����������������[�����������          .   �� ����	       	  	�   & AG� �   �   
           �f�                                                                                                                                                                                                                                                                                                                                    p L L   w    p                 !�� !��                                                                                                                                                                                                                        Y   �� �~ ��      �� ?    
������������ ����� ��������������������������� ������������������� �����  ������� ������������������������� �����  �������������������� �� � ����������������������� � ������������������������������������������������������� ����������������� �������������� ��� ���������������� ��������������  � �������������������������� � ���� ����� ����������� � �������������������� �������� �������  ����������� ������� ������������������������������ �������   ����� �  ���   �� �     $���������������������������������������������������ƫ��f���f���f������˻�fff�fffffffffffffffffff��������f˻�ff�fffffffffffffffff������������ɚ��l���fʹ�fɺ�fj�����������������������������������x��������������������wy����������ff��ff��ff��ffyffl�lfh�l�e�f�efffffffff��f�uz�UUX�UUU�UUW�UU��ffffffflfff�ffl��l̼������������fl��ff���fʺzf���f��������ɻ�vʻ�����������������������x�������x��x������������������������������ffǖffg�ffǜffŋffg�ffe�ffe�ffgUUw�UUw�UUW�UUy�UW��UX�fUY��Uy������y���z��Ƽ��fʚ�lk��jf��l˅y�xvj�f�j�l�j�f�i�f�j�Ƹʫ�w˫�u̪��x��������x���x������������������������������x��wx���������w��y�ˋi��W����U�h�U�jWUyfUu�f�X�ff�UUU�UUUzUUWxUUW�UUw�UU��UU��UU�x�UX��UW��UY��XY����̹x�i�W��Uy����������������ƺ����������̪˺˻�����������˺����ɫ������z�ʗ������z����x����������������������l�ffj�fff�fff��ff���f�̼ffʻf����UUwwUUUW�UwX�UwweU�whUUUlUUUfUUUx��f�fff���̗X��x���y���x���w���l�j�k�̵�˦f�ʻ��˻��̻��l��fl�U{˼�����l����fff�˻��̘��uUUUU��w�ʪ�ʩ�X�uUUUUUUUW��fffff�ffgZf��������UUW�UUU���W�ffU�ffU�ff�zf�UWg�UWūUW�v�U�[�U�X�y�XuX�W�Ux������̚��Ɗ��f��lf�l�l����x�˅�l��f�Wff�Vffu�fiWff�VffU�ffZfff�fffffffffffffffffffffffffffffff$�I    :      >     ��                       \     �   ���������J    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$ ^h  ��     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@       �           ��  �h  �  �����2���J J  � �� U ��� �  ���  �         ��   ���� j� = �� j� = �$ ^$         �� d��           +C��m|��           ����J  �&  yf  y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �   3       �  �3 3�=������<��̼��� �3 33==ƙ�<ə�ƙ�3ƙ��ƙ���i� 3= ��3=�l�ә��<��l<��l<��l<���<    �   3=  �30 ��� ���=��������                        +   3     0  �<  3� 3� =� =� 0� 0������������������3�33033�0�3�0��;f��;��̽�������3��3��<���<�f���̳=�=�������3303<�<00�<30�3����������������=��=��3�3�=�3�0  �=  �3  �3� ��0 ̳0 �0 �0  0� =� =� 3�  3�  �<  0  33�0�3�0�3�0�3303�303�303�303303��<���0<��0<033<033003300330033030�30�<00�<0330333033303330333033�0��<���0�03303303=03=03��0 ̳0 ��0 �3� �3� �=  0  3�     �                           <�03=��3=�� 3��  �=  �        033003300330�330��303= ��33    330333033303330333<��333ݰ    0=�0<3���;�3 �=  3�             �                           wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                                    �����   �   �   �   ����                                     	�  		  	 � 	 	 	   	   	   	   	  ��                  ��   	   	   	   	   	   	 	 	 � 		  	�                 �   	    �   	    �   	    �   	   	   �  	   �  	   �  	   �                                                       �����   �   �   �   ����                                     
�  

  
 � 
 
 
   
   
   
   
  ��                  ��   
   
   
   
   
   
 
 
 � 

  
�                 �   
    �   
    �   
    �   
   
   �  
   �  
   �  
   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    "! ""! " "" """ "!   " ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """               "  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                        ""   "! " ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                          �  �  �  �  �  �w �� �� ɪ �˙ ����������ٙ�ڪ�٘���TK�UZ� ET� 4UJ EJ D� �ܻ ��� ڙ �� �"�  �" ""  �"   �   �   �   �   �   }   p   �   �   �   �   �   �   �"  ۲  ۲  ��  �   @   T   �   �   D   �   ��� �   �  /�  "/� "" ""� ���         0 2 !2 #!0 #      �  �   �   ��  �                               �   �       ����   �       �                                   �    ���  ��                    ��  ��  ���  �  �  �   �   ��  �                            �   ���                            �   �                                                                                                                            ��	����ɪ�ܙ����ݼ "-� "� J.��#��C>Z�C U�D �Z�#�U"�C"�� ���                �  �˰ ̻� �wp ׶� �vp �w� ɪ� ��� ��� �ۙ ��� �
� �" 0�" 0.�@ "�            ����˰ + �"  "" "  � �     �  �  ��  �   �           �          �  �� ��� ��   �                    �   �   �   �  �� 	  
  �  ",  ""  �"   "                      ��  ��  �          ���� ��� ����                                    � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                                 �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                 �� �̽���ݪ۽w�}�֪�vv���p���    �   �                                �   �       �    �                     �   �  �  �                    ��  ��  ���                         ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                                 �   �  �  �  ��  ��  C�  U=  UJ  DZ  D  E  �4 
�: ���+��"��""� """ ""   �   �                        ɪ��ɪw̚�p�������������˻��۽��ݸ�̲-ۻ"""�""�2"�@  �C  �D  �T  D@  �   �   �   "�  "     �� �  �                                        ܰ ˻ �ݚ��w{`  g`  w                      �  �  ��"� ��� "                                  �   �                      �������  ���    �              �  �� ��  �    � ���                                                �   ���                            �   �                                                                                                                         	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                                   ��                  �                        ���� ��� ����                            ��  ��  ���   ���� �                                                                                                                                                                                       �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���         �  �  ��  �   �                     �� �� �� �� �݉���̙�  ���                              �������  �                     �  �   �  �  ��  �  ��  �                                                                                                                    �  �  ��  �                                                                                        �  ɪ� ɪ� ̚� �ȍ ͷ  "�  "� .( 3># �4�
�T��T�"�UN"�UN(�Dɜ� ʨ����, � /�������� � ��                                ��  ��  ��  g}  �א vz� gz� ̊� �ɩ 8̜ D<� T� @��  �� ɀ ��  ��  "   .          �  ��� �������  ��                           "  "  "  "                       �  ��  ��  ww  ��  vv  w        �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                �"�!/"�  �                                                                                                                                                                                  ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r`"   "  !�    ��                              �                        ���� ��� ����                              �   �      ��   �  ��  �  �  �         � �������������  �                � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                              �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �          
 "� ""� ""� "                       �                             ���                         �  ��                    �����                         �     �                                       �   ���                            �   �                                                                                                                 �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                /���"/�  ��                    �                                                                            �               �  �  ��  �   �   �                               ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                         �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��  ��  �   ��  �                    �     �                                       �   ���                            �   �                                                                                                          �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��                   �   ��� �̰         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
�b �c~ � � c� � �c� � c�� �c� � � c� � � c� � � 	c� � � 
c� � � c� � �cV � �c^ � �C.Z �C6j �
c� � c�	 | c�	 {	�$ {	�; ��" ��M eKg } K_ �"�U � "�g �"�Q �*�` �"�r � "�� ��r � 
��+!� � �"� � �#� � �$": � � %"P � �&!� � �'"* | �("< � �)"2 | *"@ |& +"P �N ,"& |^  "* |^  "  |& /"J �^  "  |N 1"& |^  "* | � 3"A � 4"P �$  " ~)  " { � 7*O~ � 8*K~  )�~ � :*K~  )�~ �<*$X �=* p � >"K x  !� p3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.����������������������������������������� ��5�K�\�O�T��=�U�J�J� � � � � � � � � � �/�.�7�����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������2�0�.� ���������������������������������������/�.�7�	�
�������������������� � � � � � �����������������������������������������%��������������������/�.�7� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�A�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                