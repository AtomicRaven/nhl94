GST@�                                                            \     �                                               T���       �  �            ���2�������ʰ������������������        �g     #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"��   " `  J  jF��    "�j "����
��
��     �j�� 
   ��
  ��                                                                              ����������������������������������      ��    bb= QQ0 4 111 44              		 

                     ��� �   � �                 nn ))
         88�����������������������������������������������������������������������������������������������������������������������������o  b  o   4  +c  c  'c            �        	  
      	G  7�  V(  	(                  n  1          :8 �����������������������������������������������������������������������������                                ��  �   �  z�   @  #   �   �                                                                                '        )n)n
  1n    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�9O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE E �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    `(i@�pT@��P8I@`$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `(i@�pT@��P<J@`$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `(i@�pT@���<J@`$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `(i@�pT@���<J@`$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `(i@�pT@���<J@`$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,i@�pT@���<J@`$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,i@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,i@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,i@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,i@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,i@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,i@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,i@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YC�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,j@�pT@���<J@`$YA tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pT@���<J@`$YA tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pT@���<J@`$YA tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pT@���<J@`$YA tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pT@���<J@`$YA tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pT@���<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pT@���<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pT@���<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,jK�pTL����<J@`$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,jK�pTL����<JK�$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,jK�pTL����<JK�$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,jK�pTL����<JK�$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,jK�pTL����<JK�$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,jK�pTL����<JK�$Y@�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,jK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,jK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,jK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,jK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pTL����<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pT@��@<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pT@��@<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,iK�pT@��@<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,iK�pT@��@<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,iK�pT@��@<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,iK�pT@��@<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,iK�pT@��@<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,iK�pT@��@<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,iK�pT@��@<JK�$YK�tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   F �P +���6A�#�E� `W�`8
0g� ��
�X3� T0 k� ����&�1D"3Ad 59)4#Q  ��   �   AF �P +���7A�#�E� `W�p8
0g� ��
�\3� T0 k� ����&�1D"3Ad 59)4#Q  ��    �   @F #�P +���7A�#�E�$`W�p8
0g� ��
�`3� T0 k� ����&�1D"3Ad 59)4#Q  ��    �   ?�F '�P /���8D�#�E�$`W�p8
0g� ��
�h3� T0 k� ����&�1D"3Ad 59)4#Q  ��    �   >�F /�P /���9D�#�E�$`[�p8
0k� ��
�t3� T0 k� ����&�1D"3Ad 59)4#Q  ��    �   =�F 3�P 3���9D�#�E�$`W�p8
0k� ��
�x3� T0 k� ����&�1D"3Ad 59)4#Q  ��    �   <�E�7�P 3���:D�#�E�(`W�p8
0k� ��
р3� T0 k� ����&�1D"3Ad 59)4#Q  ��    �   ;�E�;�P 3���:D�'�E�(PW�p8	0o� ��
ф3� T0 k� ����&�1D"3Ad 59)4#Q  ��    �   :�E�C�P7���:D�'�E�(PW�p<	0o� ��
ь3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �   9�E�G�P7���:D�'�E�(PW�p<	0o� ��
ѐ3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �   7�E�K�P7���;D�'�@o(PW�p<0o� ��
ј3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �   5�E�W�P;���;D�'�@o(PS�p<0s� ��
Ѥ3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �   3�E�[�P;���;D�'�@o(PS�p@0s� ��
Ѭ3� T0 k� ���&�1D"3Ad 59)4#Q  ��)    �   1�E�c�B�;���;D�'�@o(PO�p@0s� ��
Ѵ3� T0 k� ���&�1D"3Ad 59)4#Q  ��)    �   /�E�g�B�;���;D�+�@o(�O�p@0w� ��
Ѽ3� T0 k� ���&�1D"3Ad 59)4#Q  ��)    �   -�E�o�B�?���;D�+�@o(�K�p@0w� ��
��3� T0 k� ���&�1D"3Ad 59)4#Q  ��)    �   +�E�w�B�?���;D�/�@o(�G�pD0w� ��
��3� T0 k� �	��	&�1D"3Ad 59)4#Q  ��)    �   )� E���B�C���;D�3�@o(�C�pD0w� ��
��3� T0 k� �	��	&�1D"3Ad 59)4#Q  ��)    �   '�$E���B�G��;E3�@(P?�pD0w� ��
��3� T0 k� �	��	&�1D"3Ad 59)4#Q  ��)    �   %�$E���B�G��;E3�@(P;�pD0w� ��a�3� T0 k� �	��	&�1D"3Ad 59)4#Q  ��)    �   #�(E���B�G��;E7�@(P;�pD0{� ��a�3� T0 k� �	��	&�1D"3Ad 59)4#Q  ��	    �   !�(E���B�K��;E7�@(P7�pD0{� ��a�3� T0 k� �
��
&�1D"3Ad 59)4#Q  ��	    �   �,E���B�K��;E;�@(P3�pD0{� ��b 3� T0 k� �
��
&�1D"3Ad 59)4#Q  ��	    �   �0E���B�K�>�;E;�@(P/�pD0� ��b3� T0 k� �
��
&�1D"3Ad 59)4#Q  ��	    �   �4E���B�K�>�;Eo?�@(P'�pH0� ��b3� T0 k� �
��
&�1D"3Ad 59)4#Q  ��	    �   �8E���B�O�>�;EoC�@(P�pH0� ��b 3� T0 k� �
��
&�1D"3Ad 59)4#Q  ��	    �   �<E���B�O�>�;EoC�@(P�pH0�� ��b(3� T0 k� �
��
&�1D"3Ad 59)4#Q  ��	    �   <E���B�O�>�;EoC�@(P�pH0�� ��03� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �   @E���B�O�n�;EoC�@(@�pH0�� ��83� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �   DE���B�O�n�;EoG�@$@�pH0�� ��@3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �   DE���B�S�n�;E_G�@$@�pL0�� ��H3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �   HE���B�S�n�;E_G�@$@�pL0�� ��P3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �    LE���B�S�n�;E_G�@$O��pL0�� ��\3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �    LE���B�S�
�;E_G�@$O��pL0�� ��d3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �    PE��@`S�
�;E_G�@$O�pL0�� ��l3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �    TE��@`S�
�;E_G�@$O�pL0�� ��t3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �    TE��@`S�
�;E_G�@$O�pL0�� ��|3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �    XE��@`S�
�;KG�@$��pP0�� ���3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �    XE�#�@`S�
�;KG�@$�ۂpP0�� ���3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �    \E�'�@�S�
�;KG�@$	�ׂpP0�� ���3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �   \E�/�@�S�
�;KG�@$	�ρpP0�� ���3� T0 k� ���&�1D"3Ad 59)4#Q  ��	    �   `E�3�@�S�
�;KG�B�$	�ˁpP0�� ���3� T0 k� ���&�1D"3Ad 59)4#Q  �	    �   dE�?�@�S���;K?G�B�(	O��pP0�� ���3� T0 k� ���&�1D"3Ad 59)4#Q  �	   �   hE�C�A S���;K?G�B�(	O��pP0�� ���3� T0 k�  ���&�1D"3Ad 59)4#Q  ��    �    hE�G�A S���;K?G�B�(	O��pT 0�� ���3� T0 k�  ���&�1D"3Ad 59)4#Q  ��    �    lE�K�A S���;K?G�D�(	O��pT 0�� ���3� T0 k�  ���&�1D"3Ad 59)4#Q  ��    �    lE�S�A S���;K?G�D�(	O��pT 0�� ���3� T0 k�  ���&�1D"3Ad 59)4#Q  ��   �    pE�W�A S���;D�G�D�,	O��pT 0�� ��� 3� T0 k�  ���&�1D"3Ad 59)4#Q  ��    �    pE�[�APS���;D�K�D�,
O��pT 0�� ��� 3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �tE�[�APS���;D�K�D�,
O��pT 0�� ���!3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �xE�_�APS���;D�K�D�,
��pW�0�� � �!3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �|E�c�APS���;D�K�D�0��pW�0�� � �"3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �|E�g�APS���;D�O�D�0��p[�0�� �  "3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   ��E�g�A�S���;D�O�D�4��p[�0�� � "3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �E�k�A�S���;D�O�D�4�p[�0�� � #3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �E�k�A�S���;D�S�D�8{�p[�0�� � #3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �E�o�A�S���;D�S�D�8w�p[�0�� � $3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �E�o�A�S���;D�W�D�<o�p[�0�� �  $3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �E�o�D�S���;D�W�D�@k�p[�0�� � (%3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �E�s�D�S���;D�[�D�@g�p[�0�� � ,%3� T0 k� ���&�1D"3Ad 59)4#Q  ��    �   �E�s�D�S���;D�[�D�Dc�p[�0�� � 4%3� T0 k� ���&�1D"3Ad 59)4#Q  ��/    �   �E�s�D�S���;D�\ D�D_�p_�0�� �<&3� T0 k� ���&�1D"3Ad 59)4#Q  ��/    �   �E�s�D�S���;D�`D�H[�p_�0�� �@&3� T0 k� ���&�1D"3Ad 59)4#Q  ��/    �   �E�s�A�S���;D�`LLW�p_�0�� �D'3� T0 k� ���&�1D"3Ad 59)4#Q  ��/    �   �E�s�A�S���;D�dLPS�p_�0�� �L'3� T0 k� ���&�1D"3Ad 59)4#Q  ��/    �    �E�s�A�S���;D�hLPO�p_�0�� �P'3� T0 k� ���&�1D"3Ad 59)4#Q  ��/    �    �L1s�A�S���;D�lLTK�p_�0�� �X(3� T0 k� ���&�1D"3Ad 59)4#Q  ��/    �    �L1s�A�S���;D�pLXG�p_�0�� �\(3� T0 k� ���&�1D"3Ad 59)4#Q  ��/   �    �L1s�F S���;D�pLXC�pc�0�� �`)3� T0 k� ���&�1D"3Ad 59)4#Q  ��/    �    �L1s�F S���;D�tL\?�pc�0�� �h)3� T0 k� ���&�1D"3Ad 59)4#Q  ��/    �    �L1w�F S���;D�tL`;�p` 0�� �l)3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    �L1w�F W���;D�xL`7�p` 0�� �p*3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    �L1w�F W���;D�|Ld3�p` 0�� �x*3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    �L1w�E�W���;D�|Ld/�p`0�� �|*3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �L1w�E�[���;D��	Lh+�pd0�� ��+3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �L1w�E�[���;D��
Lh+�pd0�� ��+3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LAw�E�_���;D��Ll'�pd0�� ��+3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LAw�E�_�� ;E�L�l#�pd0�� ��,3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LAw�@_��;E�L�p�pd@�� ��,3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��LAw�@c��;E�L�p�pd@�� ��,3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��LAw�@c��;E�L�t�pd@�� ��-3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��LAw�@c��;E�L�t�ph@�� ��-3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��LAw�@g��;E�L�x�ph@�� ��-3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��LAw�@g�� ;E�L�x�ph@�� ��-3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��LAw�@k��$;E�L�|�ph@�� ��.3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��LA{�@k��(;E�L�| �ph@�� ��.3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��LA{�@k��,;E�L��!�ph@�� ��.3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   � LA{�@o��0;D��L��!�phP�� ��/3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   � LA{�@o��4;D��L��"��plP�� ��/3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LA{�@o��8;D��L��"��plP�� ��/3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LA{�@s��@;D��L��#��plP�� ��/3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LA{�@s��D;D��L��$��plP�� ��03� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LA{�@s��H;D��L��$��plP�� ��03� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LA{�@s��L;D��L��%�plP�� ��03� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LA{�@s��P;D��L��%�plP�� ��03� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LA{�@s��T;D�� L��&�plP�� ��13� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LA{�@s��X;D��!L��&�ppP�� ��13� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   � LA{�@s��\;D��#L��'��pP�� ��13� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �  LA{�@s��`;D��%L��'��pP�� ��13� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �$!LA{�@w��d;D��&L��(��pP�� ��13� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �$"LA{�@w��d;D��(L��)��pP�� ��23� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �(#LA{�@w��h;D��*L��)ߊ�pP�� ��23� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �($LA{�@w��l;D��,L��*ߊ�pP�� ��2"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,%LA{�@w��p;D��-L��*ۋ�pP�� ��2"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,&LA�@w��t;F�/L��*׋�pP�� ��3"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,'LA�@{��x;F�1L��+׋�pP�� ��3"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �0(LA�@{��|;F�3L��+Ӌ`tP�� ��3"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �0)LA�@{���;F�4L��,Ӌ`tP�� � 3"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �0*LA�@{���;F�6L��,ϋ`tP�� � 3"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �0+LA�@{���;F�8L��,ϋ`tP�� �4"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �4,LA�@{���<F�:L��,ˋ`tP�� �4"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �4,LA�@{���<D� ;L��,ˋ`t	P�� �4"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �4-LA�@���<D�=L��,ǋ`t	P�� �4"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �4.LA�@���<D�?L��,ǌ`t	P�� �43� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   �8/LA�@���=D�@L��-Ì`t	P�� �53� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �80LA�@���=D�BL��-Ì�t	P�� �53� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �81LA�@���=I�CL��-Ì�x	P�� �53� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �82L1�@���=I�EL��-���x	P�� �53� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �<3L1�@���=I�FL�-���x
P�� �53� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   <3L1�@����>I�GL�-���x
P�� � 53� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   <4L1�@����>I�IL�-���x
P�� � 63� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   <5L1�@����>J JL�-���x
P�� �$63� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   @6L1�@����>J  KL�.���x
P�� �$63� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   @7E��@����>J  LL�.���x
P�� �(63� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   @7E��@����?J $MDߴ.���x
P�� �(6"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   @8E��@����?J $NDߴ.���xP�� �,6"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   D9E��@����?I�$OD߸.���xP�� �07"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   D9E��@����?I�$PD߸.���xP�� �07"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   D:A��@����?I�(QD߼/���xP�� �47"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   D;A�{�@����@I�(QD߼/���|P�� �47"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   D<A�{�@����@I�(RD��/���|P�� �87"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   H<A�{�@����@J (SD��0���|P�� �87"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   H=A�{�@����@J (SD��0���|P�� �<7"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   H>A�{�@����@J (TD��0���|P�� �<8"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   H>A�{�@����AJ (TD��0���|P�� �@8"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   H?D�w�@����AJ (UD��0���|P�� �@83� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   H?D�w�@����AI�(UD��1���|P�� �D83� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   L@D�w�@����BI�(VD��1���|P�� �D83� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   LAD�w�@����BI�(VD��2���|P�� �H83� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   LAD�w�L�����BI�(VD��2���|P�� �H83� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   LBD�w�L�����BI�(WD��2���|P�� �H83� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   LBD�w�L�����CJ (WD��2���|P�� �L93� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   PCD�s�L�����CJ (WD��3���|P�� �L93� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   PDD�s�L�����CJ (WD��3���|P�� �P93� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   PDD�s�L�����DJ (WD��4����P�� �P93� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   PED�s�L�����DJ (WD��4����P�� �T93� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   PED�s�L�����DI�(WD��5����P�� �T93� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   PFD�s�L�����EI�(WD��6����P�� �T93� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   PFD�s�L�����EI�(WD��6����P�� �X93� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   TGD�o�L�����EI�(WD��7����P�� �X93� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   TGD�o�L�����FI�(WD��8����P�� �X:3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   THD�o�L�����F@(WD� 8����P�� �\:3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   THD�o�L�����F@(WE�9����P�� �\:3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   TID�o�L�����G@(WE�:����P�� �`:3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   TID�o�L�����G@(WE�;����P�� �`:3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   XJD�o�L�����G@(WE�<����P�� �`:3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   XJD�o�L�����G@(WE�=����P�� �d:3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   XKD�k�L�����H@(WE�>����P�� �d:3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   XKD�k�L�����H@(WE� >����P�� �d:3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   XKD�k�L�����H@(WE�$?����P�� �h:3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �XLD�k�L�����IK�(WEp,@����P�� �h;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �XLD�k�L�����IK�(WEp0A����P�� �h;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �XMD�k�L�����IK�(WEp4B����P�� �l;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\MD�k�L�����IK�(WEp8D����P�� �l;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\ND�k�L�����JK�(WEp<E����P�� �l;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\ND�k�L�����JK�(WEpDF����P�� �l;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\ND�k�L�����JK�(WEpHG����P�� �p;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\OLQg�@����JK�(WEpLH����P�� �p;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\OLQg�@����JK�(WEpPJ����P�� p;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\PLQg�@����KK�(WEpTK����P�� t;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\PLQg�@����KK�(WEpXL���P�� t;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\QLQg�@����KK�(WEp\N���P�� t;3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �XRLQg�@����KK�(WE``O���P�� t<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �XRLQg�@����LK�(WE`dP���P�� x<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �XSLQg�@����LK�(WE`hR���P�� x<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �XTLQg�@����LK�(WE`lS{���P�� x<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �TULQg�@����LK�(XE`lU{���P�� |<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �TULQg�@����LK�(XE`pV{���P�� |<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �TVLQg�@����LK�,XE`tX{���P�� |<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �PWLQc�@����LK�,XE`xY{���P�� |<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �PXLQc�@����LK�,XE`x[{���P�� |<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LYLac�@����LK�,XE`|\w���P�� �<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �LZLac�@����LK�,XE`|^w���P�� �<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �H[Lac�@����MK�,XEP�_w���P�� �<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �D[Lac�@����MK�,XEP�aw���P�� �<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �D\Lac�@����MK�,YEP�bw���P�� �<3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �<^Lac�@��� MK�0YEP�ew���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �8_Lac�@��� MK�0YL�gs���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �4`Lac�@��� MK�0YL�hs���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �0`Lac�@��� MK�0YL�js���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �0aLac�@��� MK�0YL�ks���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �(bLac�@��� MK�0YL�ls���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �$cLac�@��� MK�0YL�ns���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   � cLa_�@���MK�0YL�os���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �dLa_�@���MK�0ZL�ps���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �eLa_�@���NK�0ZL�qo���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �fLa_�@���NK�4ZL�so���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �fLa_�@���NK�4ZL�to���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �gLa_�@���NK�4ZL�uo���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �hLa_�@���NK�4ZL�vo���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��hLa_�@���NK�4ZL �wo���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��iLa_�@���NK�4ZL �yo���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��jLa_�@���NK�4ZL �zo���P�� �=3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��jLa_�@���NK�4ZL �{k���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��kLa_�@���NK�4ZL �|k���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��lLa_�@���NK�4ZL �}k���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��lLa_�@���NK�4[L �~k���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��mLa_�@���NK�8[L �k���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��mLa_�@���NK�8[L ��k���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��nLa_�@���NK�8[L ��k���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �nLa_�@���NK�8[L ��k���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �oLa_�@���NK�8[L �k���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �oLa_�L����NK�8\L �k���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �oLa[�L����NK�8\L �g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   �nLa[�L����NK�<\L �g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �nLa[�L����NK�<\L ��g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �nLa[�L����NK�<\L �g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��nLa[�L����NK�<]L �g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��mLa[�L���� NK�<]L �g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   ��mLa[�L���� NK�<]L �g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   ��mLa[�L����$NK�@]L �~g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   ��lLQ[�L����$NK�@]L �~g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �xlLQ[�L����$NK�@^L �~g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �tkLQ[�L����(NK�@^L �~g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �lkLQ[�L����,NK�@^L �}g���P���>3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �lkLQ[�L����,NK�@^L �}c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   	�hkLQ[�L����0MK�<^L �}c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   	�dlD�[�L����0MK�<^L �}c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   	�`lD�[�L����0MK�<^L �}c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   	�\lD�[�L����0MK�<^L �|c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   	�\lD�[�L����4MK�<^L �|c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   	�\lD�[�L����4MK�<^L �|c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   	�\lD�[�L��� 4MK�<^L �|c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   	�\lD�[�L��� 4MK�<^L �|c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   	�\lEq[�L��� 4MK�<^L �{c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   	�\lEqX L��� 4MK�<^L �{c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lEqXL��� 4MK�<^L �{c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lEqTL��� `4MK�<^L �{c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lEqTL��� `4MK�<^L �{c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1TL��� `4MK�<^L �{c���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1T@�� `4MK�<^L �zc���P���?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1T@�� `8MK�<^L�z_���P��|?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1P@��@8M@<^L�z_���P��|?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1P
@��@8N@<^L�z_���P��|?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1P@��@8N@<^L�z_���P��|?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1P@��@8N@<^L�z_���P��|?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1P@��@8N@<^L�y_���P��|?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1P@��@8N@<^AP�y_���P��|?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1L@��@8N@<^AP�y_���P��x?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1L@��@8N@<^AP�y_���P��x?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1L@��@8N@<^AP�y_���P��x?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1L@�� �8N@<^AP�y_���P��x?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lL1L@�� �8N@<^C��x_���P��x?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lLAL@�� �8N@<^C��x_���P��x?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lLAH@�� �8N@<^C��x_���P��x?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lLAH@�� �8N@<^C��x_���P��x?3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lLAH@�� �8N@<^C��w_���P��t@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lLAH@�� �8N@<^C��w_���P��t@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lLAH@�� `8N@<^C��v_���P��t@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lLAH@�� `8N@<^C��v_���P��t@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   �\lLAD@�� `8N@<^C��u_���P��t@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lLAD@�� `8N@<^C��u_���P��t@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �\lLAD@�� `8N@<^C��t[���P��t@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P\lLAD@�� `8N@<^C��t[���P��t@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P`lLAD@�� `8N@<^C��t[���P��p@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P\lLAD@�� `8N@<^C��t[���P��p@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P\lLAD@�� `8N@<^C��s[���P��p@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P\lLAD @�� `8N@<^C��s[���P��p@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P\lLA@!@�� `8N@<^C��s[���P��p@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P\lLA@!@�� `8N@<^C��r[���P��p@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P\lLA@"@�� 8N@<^C��r[���P��p@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P\lLA@#@�� 8N@<^C��r[���P��p@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   P\lLA@$@�� 8N@<^C��r[���P��p@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P\lLA@$@�� 8N@<^C��r[���P��p@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   `\lLA@%@�� 8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA@&@�� 8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA@&@�� 8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA<'@�� 8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA<(@�� 8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA<(@�� 8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA<)@�� 8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA<*@�� 8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA<*@��@8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA<+@��@8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA<+@��@8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA<,@��@8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA<-@��@8N@<^C��r[���P��l@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA8-@��@8N@<^C��r[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA8.@��@8N@<^C��r[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\lLA8.@��@8N@<^C��r[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `\mLA8/@��@8N@<^C��q[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `XmLA8/@��@8N@<^C��q[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `XmLA80@��@8N@<^C��p[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `TmLA80@��@8N@`<^C��p[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   `TmL181@��p8N@`<^C��o[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `TmL181@��p8N@`<^C��o[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `TmL182@��p8N@`<^C��n[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `TmL182@��p8N@`<^C��n[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `TmL183@��p8N@`<^C��n[���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `TmL183@��p8N@`<^C��nW���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `TmD144@��p8N@`<^C��nW���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `PnD144@��p8N@`<^C��mW���P��h@3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `PnD145@��p8NK�<^C��mW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `LnD146@��p8NK�<^C��lW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `LnD106@��p8NK�<^C��lW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `LnD107@��p8NK�<^C��kW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `HnD108@��p8NK�<^C��jW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   `HnEa,8@��p8NK�<^C��jW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   `DnEa,9@���8NK�<^C��iW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `DnEa(:@���8NK�<^C��iW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `@oEa(;@���8NK�<^C��hW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `@oEa$<@���8NK�<^C��hW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `<oEa$=@���8NK�<^C�|hW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `<oEQ >L����8NK�<^C�|gW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   `<oEQ>L����8NK�<^C�|gW���P��dA3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P8oEQ?L����8NK�<^C�|gW���P��dA"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P8oEQ@L����8NK�<^C�xgW���P��dA"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P4oEQAL����8NK�<^C�xfW���P��dA"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P4oC�BL����8NK�<^C�xfW���P��dA"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P4pC�CL����8NK�<^C�xfW���P��dA"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P0pC�DL����8NK�<^C�xfW���P��dA"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P0pC�DL����8NK�<^C�xfW���P��dA"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P0pC� EL����8NK�<^C�xfW���P��dA"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P0pC��FL����8NK�<^C�xfW���P��dA"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,pC��GL����8NK�<^C�xfW���P��`A"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,pC��GL����8NK�<^A xfW���P��`A"s� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,pC��HL����8NK�<^A xfW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,pC��IL����8NK�<^A xfW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,pC��JL����8NK�<^A xfW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P,pC��JL����8NK�<^A xfW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,pC��KL����8NK�<^A xfW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,pC��LL����8NK�<^C�xfW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,pC��LL����8NK�<^C�xfW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,oC��ML����8NK�<^C�xfW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,oC�NL����8NK�<^C�xfW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,oC�NL����8NK�<^C�xfW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,oC�OL����8NK�<^K�xeW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,nC�PL����8NK�<^K�xeW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,nC�PL����8NK�<^K�xeW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,nC�QL����8NK�<^K�xeW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,nD �QL����8NK�<^K�xeW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,nD �R@���8NK�<^K�xeW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,nD �R@���8NK�<^K�xeW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,nD |S@���8MK�<^K�xeW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,nD xT@���8MK�<^K�xeW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �,nI�xT@���4MK�@]K�xeW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �(nI�xT@���4MK�<]K�xeW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �(nI�tT@���0LK�<]K�xdW���P��`A"�� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   �(mI�tT@���0LK�8]K�xdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (mI�tT@��p,LK�8]L xdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (mI�tT@��p,KK�4]L xdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (mI�tT@��p,KK�4]L xdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (mI�pT@��p(KK�4]L xdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (mI�pT@��p(JK�0\L xdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (lI�pT@��p$JK�0\L xdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (lI�pT@�� $JK�0\L tdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (lI�pT@�� $IK�,\L tdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (kI�pT@��  IK�,[L tdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (kI�pT@��  IK�,[L tdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (kI�pT@��  HK�,[L tdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (kAPpT@��� HK�([L tdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (kAPpT@��� GK�(ZL tdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (kAPpT@���GK�(ZL tdW���P��`A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �    (kAPpT@��� FK�$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �    (kAPpT@��� FK�$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   @(kAPpT@��� EK�$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   @(kAPpT@��� EK�$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   @(kA pT@��� EK�$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   @(kA pT@��� EK�$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   @(kA pT@��� DK�$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �(jA pT@���$D@`$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �(jA pT@���$D@`$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �(jA pT@���$D@`$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �(jA pT@���(D@`$ZL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �(jA pT@���(D@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   �(jA pT@���(D@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(jA pT@���,D@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(jA pT@��@,D@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(jA pT@��@,E@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)   �   P(j@�pT@��@,E@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(i@�pT@��@0E@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(i@�pT@��@0F@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(i@�pT@��@0F@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(i@�pT@��@4G@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(i@�pT@��@4G@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(i@�pT@��@4H@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(i@�pT@��@4H@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(i@�pT@��P8I@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(i@�pT@��P8I@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �   P(i@�pT@��P8I@`$YL tdW���P��\A3� T0 k� ����&�1D"3Ad 59)4#Q  ��)    �                                                                                                                                                                               � � �  �  �  d A�  �K����   �      6 \��� ]�11 @ � i�@   � �	   � h�     i�@ h�                   ]	 Z           ���     ���   0	&


          T�  � �	   � ��     T ��     ��          	 Z          p�  
  ���   (	 
          ����    
	     )�    ���� )�                   ? Z           b      ���   0
           Jl   4 4    ��     JV �.    ��r            Z Z           ��     ���   H$
          Y|  � �
	   / 	x     Yz 	x                    	 Z           ��    ���   03 
           d��  � �	   C ��     d� ۿ     V               R	 Z          %��  !  ���   H	D
 
          ��p�       W��ts    ��p���ts                   \ 6         �       ��@   8	 

          ��        k $�     �� $�                    i 5         ��     ��@    		�          ��          :��    �� :��                  	    ��          `�     ��B   8
)           Ϻ       � B
k     Ϻ B
k                        �         	 ?�     ��H  0
3
          A{�  � �
    �~�     A{�~�                     A �         
  
`     ��P   H


           VD ��
     � ��      VD ��                            ���g             �  ��@    		 5 	                 ��      �                                                                           �                               ��        ���          ��                                                                 �                          �{  ��        � 9�=     �{ 9�=         "                 x                j  �    	   �                              ��        � :          :           "                                                �                            )  	 �� $ : B ��� 9 :         
       	  
  �   /D 3��K       � @[� ʄ  \` �� 0\� �$ @]  ˤ ]� �� ]� �D e  �� 0i` �  i� �D j  �D  ]` �� ]���� ����  ����. ����< ����J ����X � �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }����� � � }����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����    ����  ������  
�fD
��L���"����D"� �  " `   J jF��    "�j "���
��
���     �j��  
  �
� �  �  
�      ��     � B      ��    ��     � )           ��     � B          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �)33      ��= �  ���        � �T ���        �        ��        �        ��        �  	  }�     �� ��        ��                         T�) , � ���                                      �                 ����            	  B	���&��     ��           �    26 Robert Reichel                                                                                   4  4     �TcW �lc_ � �K/S � K7[ � K8K �K9K � K;S � K<V �	B�e �
B�e �B�M �B�E � B�] � B�L �CJ � CZ �C D � C"L �J�S �J�K � J�R �J�K �J�H �KCc �KF[ � KIb �KJ[ �KLX �ck � cs �K � �  � �!c � � "c� � � #� �$c� � �%c� �&"� � � '"� �(� � �)
� �*"� � � +"� �,"� � �-*� � �."� � � /"� �0� � � 
� �2*� � �3"� � � 4"� �5� � � 
� � 
�(  "Q u  9"B u(  "Q u  ;"C u(  "K u �  "L u �>*m �  "L u                                                                                                                                                                                                                         �� P         �     @ 
        	�     c P E e  ��        	            ������������������������������������� ���������	�
���������                                                                                          ��    ��~�0� ��������������������������������������������������������   �4, >   B h�� }  �@M��@��� �"���������'�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 
  	  .    �� �D�J ��    �                             ������������������������������������������������������                                                                    
                                                                    J��� <��                                             ���������������������������� � ��������������������� ������ ����� ��� ��������������������� ������� �������������������������������� ����������������� ����� ������� ���������������� � ������������ � ������������ ������ ����������� ������� ���� � ��                                  f    %     � �\�J      e�                             ������������������������������������������������������                                                                                                                   
                   ���Y-�  �                                           ����� �������������� �������� �� �� �������������� ��� ��� �� ���������������������� ��������� ����������������������������������� �  �� ����������� ������������� ��������������������� � ��� �������� ��� ����������� ��� � ����                                                                                                                                                                                                                                                                           	                     
                             �              


            �   }�           �      8�            oW                                                         ���  S�      I  J5  =��������������������������������������������������������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � ��I �\                                                                                                                                                                                                                                                                                        )n)n
  1n        e            m                  k            `                                                                                                                                                                                                                                                                                                                                                                                                         > �  
>�  @�  2�  J�  Bm] ���������]�̞�n���������� �V W������������                      �� o        $   �   & QW  �   �                  �                                                                                                                                                                                                                                                                                                                                        K K   �   	                  !��                                                                                                                                                                                                                            Z��   �� �� ��      �� 4      ���������������������������� � ��������������������� ������ ����� ��� ��������������������� ������� �������������������������������� ����������������� ����� ������� ���������������� � ������������ � ������������ ������ ����������� ������� ���� � ������� �������������� �������� �� �� �������������� ��� ��� �� ���������������������� ��������� ����������������������������������� �  �� ����������� ������������� ��������������������� � ��� �������� ��� ����������� ��� � ����             $����������������˪�������������������������������������f��ff��ff�������̺�ff�fffffffffffffffffff����ƹ��ffʻfff�fffjffffffffffff��������������������ʺ��l���f˪������������������������������������������������������������������fff�fff�fff�ffk�ffi�ff��ff��ff�ffffffff�fff�x�����w��xx�������wfffffff�ffff�fffww��ww�x����wx��fk��ff��ff��ffʹffj��fʪ�f�ˊ�k������������ʚ��������������������������������������������˫��ʫ��ff��fl��fl��ff̫fff�ffʬ�f���f�����������wu���w��l������f����W��������xww��Wy�l����x������k���W�fi���j���j���f����˘�����y�y�y����������������������������������������������������ʻ����ʫɚ�����l���ƨ�lƘ�j���k���̜i���j���kxx���wx������wx������������ƈx����������������wW����w�������������������������z����������˫��̺������������������������������������������������������������ʺ������k������������������������������������������x�j���˙�x�˘��̩�x������x���xx�x������x������wx���˫��ʫ����������˪�����ʻ��������������������������������������ʻ�ʻ�����ʪ̫����˺��������������������˪�����f���k��f��fǶW�g���k���̻���f������������������x�������˩f̺�����uw�����w��x�wXx��˪�����������l����l���i��ƹx�f�������������������ʫUW��UUU�UUUX      @   '   :   �                         4     �   ���������J'      ��     �         �      �         �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��   ( ����  �� �� �    � �N ^$   ��B   (  ��   ) ��  � ��     � ��   	 ��   p � ��  � ��  5� �� �� �z  5� �� �$ ^$ �u�  5� ��  � ��  �` ��  ��   ��     ��   � �� ��   �z � �N ^$�� �   �          ��  �� ��  �  �� �� �z  � ��� �$ J �  ��T   �      �      �������2����  g��� 
   �     f ^�          �� ,              �����2�������J����  ��      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                                                  U  T   T   T     T UDUDDUDDDDDDDDDDDDDDDP   E�  DU� DDU�DDDUDDDDDDDDDDDD                UP  E�  E   E                                           ���U�UTD�DDDDDDTDD TDD   �   U_ DEU�DDDUDDDDD��DZT�DDDDDDDDDDDDTDDDDDDDDUTU�����DDDDDDDDDDDEDDDEDDDDTUTU�Ԫ���Z_   P   � �U�UTDUDDDDUTD�DT��D        U_��DEU_DDD_DDDPDDE�DDE  �DD DD DD �DD �UD  �U       DZTDEDDDDE�DDE�DDE�TDDT�DE�TE���DDTU�ZD���������DDTDD��ZT�T���ZTDDE��D��T�T��DUTTT��Z��TQTDDUTD�DDDTDDD�DDDDDDE�DD_TDE�DD_ DDP DDP DD_ DU_ U�  �                                       TE�DDD�UUU                    ���DDDUUUTD  D  D  D  D  U��D�TDDDDEUUDP  DP  DP  DP  UP  TDE�DDDPUUU_                                                    wwwwtDDDt""$t"""t"w"t"w"t"w"t""$wwwwtDGtD"GtD"GtD"GtD"GtD"GtD"GtwwwwDDDD"D"""D"""DD""Gt""Gt""Gt"wwwwDDDD"B"""B""DDD"GwD"GwB$GtB$wwwwDwww$www$wwt$wwtGwwtGwwwwwwwwwwwtDDDD�DLL�D���D�D�D�t�D�t�D�wwwwDDww��Gw��Gww�Gww�Gww�Gww�Gwt"""t"w"t"w"t"w"t"""t""$tDDDwwwwD"GtD"GtD"GtD"DDD""$D""$DDDDwwww"Gt""Gt""Gt""Gt""Gt""Gt"DGtDwwwwGt"DGD"DGB$GGB$DGB""GB""GDDDwwwwwwwwwwwwwwwwDwww$www$wwwDwwwwwwwt�D�t�D�t�D�t�D�t�D�t�DMtDDDwwwww�Gww�Gww�Gww�Gw��Gw��GwDDwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG      w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  " ! " ""  "!  " ! " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  "!  " ! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  " ! " ""  "!  " ! " ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                           �  ��� ݻ� g�� bm� ggz�'w���������������˛������ˊۼ�����˻������H�DH�@U�DPT�E X�T H�P H�@ Ȥ� ̻� ˘ "�� � ���/�"" �""/���               �   �                                                     �  �                      � �                       ���           �                      "  "             ��.�  .                 ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                       �   ���                            �   "                                                                                                                 � ��� ��� ܷz �riwgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �        "   "   "      "   "   "�  �           �   �   �                                                  �               �     "   "                   �     �                    ""�""  ""  / �   �               � � ��      �                                                                                                             �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   U�  U�  EP  L�  ɀ ��  �� �+" �                                                  �� �� ��               �  �  �     "   "                                �  ".��".� ��                        ���                  ""  "".  . �    �                                                                                                                                                       � ̻ �ۼͺ�	ۚ����C�˽T;��UJ��ET�35J�D3T�  ̰ ̻	�̻���w���&��wv��wpʨ� ��� ��� ��  "�� .� "�� ��0 "          .  .  "   "             �  �� ʝ ,��+� "" "��CEJ�D5J� J�  �� 
�� �  �� �+� �"" """����    �         ""�"" �  ��                /���"/�  ��                    �                                                                            �               �     "   "                   �     �                                                                                                                                                                                   "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             �"  �""� "�    �     �                                                                                                                                                                                                  � ��� ��� ܷz �riwgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �        "   "   "      "   "   "�  �           �   �   �                                                  �               �     "   "                            �  �˰ ��� �wp �&                                                                                  �  �  "   "                                                                                  �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp��& ��vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �" �"" �"   �                    .   .   �        �  ��  ��  ww  &'  vv  w                �                        ��"� �"� ����                            �    � �  ��                  ���                � "�"  �    � � �                                                                                                                                   �� ��� ��� ww� &'� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                               " "/ �/� ��     �   "           "   �                    �� �� �� w� b| �"  "  "   �.  �   �                     "  ""  """"""
�                               	�  �       �                            ""  "".  . �    �                                                                                                                                       	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��               �   �   "           �   �   �                                       �  ���          "   "   "                                �   �      ��   �  ��  �  �  �         � ".��".��/����  �                                �   "                                                                                                                 �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp��& ��vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �" �"" �"   �                    .   .   �     .  " "" ��� "                                  �   �                      �".��".  ���    �                    �    � �  ��                  ���                                 ����     �   "  "     "   "   �                           ��   ��                  .  .  "  " ��                                                    
�  	�  �� 	˼ 
�� ���̍��ݻ�	�""�" 4�"#ETUD�DD��D 	�@ 
��  ��  �  �  ""  "!���  ��         ��  ��  ��  w�  b|  gw  w�� ��� �����ɪ��͙�̽�̻����݊���������2,̠",� "*@ B*@ 5�@ 4�  �� ̀  ��  �� �,  "/��"� �!��  ��                  �   �        �   �     �   � �.  .�� �                          "  �"  �         �  ��� ̻� ��� rbp wgz�       �".��".���                                  "  .���"    �     �                   ���������������������  ��  ��  ��  �   �    �          �         �                                                                                                              �� ̻ ��˛��  �� �˚̻���ۚ����I���䘼�^���^�٘�:�^�� ^�� D�( �) �) �) ��) ˹� ț�+��,��,����  �𫒒 ��� �ɍ ��ݨ��ډ�݊�� ��D@ �D�  J�� ݩ� ��� �ۻ �ک �ڹ�ɻ��̸���������� ����������            �   ��  ��  ��  ��  ��                                          .� ".� "/� /�  �                         �   �                        �� ̻ ��          �   �"           �    �         �  �      �           �                        �         �  "� "  �  ��                                                                                                                                                 2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD l � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=GwDGwqwDDwtwwww3333DDDD  � �!�aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( """"����������A��I��I X � �!�aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx""""�����A�DA�I��I� w � �!�aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""��������I���I���I���I��� � � �!�aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(MAMAMMMM�M�M����3333DDDD  � �!�aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�D�����MD��M����3333DDDD m � �!�a�a� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� Sa��m(`���4���4���4���4���4���43334DDDD � � �!�aa � � � �!i!j � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� Sa��(M""""wwwwqqqqwGwGGG � � �!�aa � � � �!m!n � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� Sa�� 
(�""""wwwwwwqqDAwG � u!�!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� S)��(-(�������������������333DDD!�!�!�!�!�!� �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5M��M��D��M����������3333DDDD!�!�!�!�!�!� � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDD��D�M��D����3333DDDD!�!�!�!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���rs��ww""""������DH�H�!�!�!�))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�tu���(+""""�������H�H��D!�!�!�5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�vw��(W(�""""��������H��H��H��H�� !�!�AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���&2�(a(�DD������L��DL����3333DDDD;'(!�AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(�L�A�AAD��DL�����3333DDDD<34!�AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� SA��l(=���4���4���4L��4L��4���43334DDDD  � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� SA��(( """"���������M�MMM X � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� SA��(Xx""""�������A��AA w � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� )��:	9ww��������������333DDD � � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(I��I����������������3333DDDD  � �!�AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((���A���I��I���I�����3333DDDD m � �!�A�A� � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""������������������������  � �!�AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M""""������D�D��� 
 � �!�AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�""""������������������������ - � �!�!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�wqwwqwwwwwqwwwDwwww3333DDDD 69�:���  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5qqwwwDDwtGwwww3333DDDD � � � i i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+www4www4www4www4www4www43334DDDD W � � u u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(�""""wwwwwwqwwwqwqwq a � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(�""""wwwwwwwDwGwA  � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(��A�L�L�L��L���333DDDLDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDDTcW �lc_ � �K/S � K7[ � K8K �K9K � K;S � K<V �	B�e �
B�e �B�M �B�E � B�] � B�L �CJ � CZ �C D � C"L �J�S �J�K � J�R �J�K �J�H �KCc �KF[ � KIb �KJ[ �KLX �ck � cs �K � �  � �!c � � "c� � � #� �$c� � �%c� �&"� � � '"� �(� � �)
� �*"� � � +"� �,"� � �-*� � �."� � � /"� �0� � � 
� �2*� � �3"� � � 4"� �5� � � 
� � 
�(  "Q u  9"B u(  "Q u  ;"C u(  "K u �  "L u �>*m �  "L u3333DDDDAqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD��������������������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ��������������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ��������������������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE��������������������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD��������������������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD��������������������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD��������������������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� ����>�L�L�T�\��=�L�S�H�U�U�L��������>��<���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� ����7�\�J��<�V�I�P�[�H�P�S�S�L�������8�>�7���""""������A�D��I��""""�������D����� ��"��<�V�I�L�Y�[��<�L�P�J�O�L�S�������>��<���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �8�>�7��� ���A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �>��<���#��""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,�����������DDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �����<�L�Z�\�T�L��2�H�T�L����������������� ����4�U�Z�[�H�U�[��<�L�W�S�H�`��������������� ����.�O�H�U�N�L��2�V�H�S�P�L���������������� ������0�K�P�[��7�P�U�L�Z���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            