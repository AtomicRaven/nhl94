GST@�                                                           @m�                                                      O��&                 
      ����e ��	 ʰ����������`���z���        �h      #    z���                                d8<n    �  ?     �����  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    B�jl �   B ��
  �                                                                              ����������������������������������      ��    =b 0Qb 4 114  4c  c  c        	 
      	   
       ��G �� � ( �(                 nnn 	)1         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                  -       �   @  &   �   �                                                                                 '      	n)n1n  �    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE - �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    @4N x@d_�B���|( C��LL^Lc���RZ4�T0 k� �7��;�%�@c  �e1t B  ��    �   �@8N x@d_�B���|( C��LL]Lc���RZ4�T0 k� �7��;�%�@c  �e1t B  ��    �   �@8N t@d_�B���|( C��LL]Lc���RZ4�T0 k� �7��;�%�@c  �e1t B  ��    �   �@8N t@d_�B���|( C��LL]Lc���RZ4�T0 k� �7��;�%�@c  �e1t B  ��    �   �@8M t@d_�B���|( C� LL]Lc���RZ4�T0 k� �7��;�%�@c  �e1t B  ��    �   �@8M t@d_�B���|( S�LP\Lc���RZ4�T0 k� �7��;�%�@c  �e1t B  ��    �   �@8M t@d_�B���|( S�LP\Lc���RZ3��T0 k� �7��;�%�@c  �e1t B  ��    �   �@8M t@d_�B���|( S�LP\Lc��S�RZ3��T0 k� �;��?�%�@c  �e1t B  ��    �   �@8L t@d[�B���|( S�LP\Lc��S�RZ3��T0 k� �;��?�%�@c  �e1t B  ��    �   �@8L t@d[�B���|( S�LP[Lc��S�RZ3��T0 k� �;��?�%�@c  �e1t B  ��    �   �@8L p@d[�B���|( S�K�P[Lc��S�RZ3��T0 k� �;��?�%�@c  �e1t B  ��    �   �@8L p @d[�B���|( S�K�T[Lc��S�RZ3��T0 k� �;��?�%�@c  �e1t B  ��    �   �@8L p @d[�B���|( S�	K�T[Lc��S�RZ3��T0 k� �;��?�%�@c  �e1t B  ��    �   �@<K p @d[�B���|( S�
K�T[Lc��S�RZ3��T0 k� �;��?�%�@c  �e1t B  ��    �   �@<K p @d[�B���|( S�K�TZLc��S�RZ3��T0 k� �;��?�%�@c  �e1t B  ��    �   �@<K p!@d[�B���|( S�K�TZLc��S�RZ3��T0 k� �;��?�%�@c  �e1t B  ��    �   �@<K p!@d[�B���|( c�C�TZLS��S�RZ3��T0 k� �?��C�%�@c  �e1t B  ��    �   �@<K p!@d[�B���|( c�C�TZLS� ��S�RZ3��T0 k� �?��C�%�@c  �e1t B  ��    �   �@<J l"@d[�B���|( c�C�XYLS�!��S�RZ3��T0 k� �?��C�%�@c  �e1t B  ��    �   �@<J l"@d[�B���|( c�C�TYLS�"����RZ3��T0 k� �?��C�%�@c  �e1t B  ��    �   �@<J l"@d[�B���|( c�C�TYLS�#����RZ3��T0 k� �?��C�%�@c  �e1t B  ��    �   �@<J l"@d[�B���|( c�E�TYLS�$����RZ3��T0 k� �?��C�%�@c  �e1t B  ��    �   �@<J l#@d[�B���|( c�E�TYD��%����RZ3��T0 k� �?��C�%�@c  �e1t B  ��    �   �@<I l#@d[�B���|( c�E�TYD��'���RZ3��T0 k� �?��C�%�@c  �e1t B  ��    �   �@<I l$@d[�B���|( c�E�TXD��(���RZ3��T0 k� �?��C�%�@c  �e1t B  ��    �   �@<I h$@d[�B���|( c�E�TXD��)���RZ3��T0 k� �C��G�%�@c  �e1t B  ��    �   �@<H h%@d[�B���|( c�E�TXD��*���RZ3��T0 k� �C��G�%�@c  �e1t B  ��    �   �@<H d&@d[�B���|( s�E�TXLS�+���RZ3��T0 k� �C��G�%�@c  �e1t B  ��    �   �@<H d&@d[�B���|( s�E�TXLS�-���RZ3��T0 k� �C��G�%�@c  �e1t B  ��    �   �@<G `'@d[�B���|( s�E�PXLS�.� ��RZ3��T0 k� �C��G�%�@c  �e1t B  ��    �   �@<G `(@d[�B���|( s�E�PWLS�/� ��RZ3��T0 k� �C��G�%�@c  �e1t B  ��    �   �@<G `(@d[�B���|( s�E�LWLS�0� ��RZ3��T0 k� �C��G�%�@c  �e1t B  ��   �   �@<F \)@d[�B���|( s�E�LWLS�1� ��RZ3��T0 k� �C��G�%�@c  �e1t B  ��    �   �@<F \*@d[�B���|( s� E�HWLS�2� ��RZ3��T0 k� �C��G�%�@c  �e1t B  ��    �   �@<F \*@d[�B���|( s�"C�DVLS�3� ��RZ3��T0 k� �C��G�%�@c  �e1t B  ��    �   �@<E X+@d[�B���|( s�#C�DVLS�5� ��RZ3��T0 k� �G��K�%�@c  �e1t B  ��    �   �@<E X,@d[�B���|( s�%C�@VLS�6�!��RZ3��T0 k� �G��K�%�@c  �e1t B  ��    �   �@<E T,@dW�B���|( s�'C�<VLS�7�!��RZ3��T0 k� �G��K�%�@c  �e1t B  ��    �   �@<D T-@dW�B���|( C�(C�8ULS�8�!��RZ3��T0 k� �G��K�%�@c  �e1t B  ��    �   �@<D T-@dW�B���|( C�*C�4ULS�9�!��RZ3��T0 k� �G��K�%�@c  �e1t B  ��    �   �@<D P.@dW�B���|( C�*C�0ULS�:�!��RZ3��T0 k� �G��K�%�@c  �e1t B  ��    �   �@<C P/@dW�B���|( C�+C�,ULc�;�!��RZ3��T0 k� �G��K�%�@c  �e1t B  ��    �   �@<C P/@dW�B���|( C�-C�,ULc�<�!��RZ3��T0 k� �G��K�%�@c  �e1t B  ��    �   �@<C L0@dW�B���|( Ӑ.C�,TLc�=�"��RZ3��T0 k� �G��K�%�@c  �e1t B  ��    �   �@<C L0@dW�B���|( Ӑ0C�(TLc�?�"��RZ3��T0 k� �K��O�%�@c  �e1t B  ��    �   �@<B L1@dW�B���|( Ӑ1C�(TLc�@�"��RZ3��T0 k� �K��O�%�@c  �e1t B  ��    �   �@<B L1@dW�B���|( Ӑ2C�(TLc�A�"��RZ3��T0 k� �K��O�%�@c  �e1t B  ��    �   �@<B H2@dW�B���|( Ӑ4C�(TLc�B�"��RZ3��T0 k� �K��O�%�@c  �e1t B  ��    �   �@<A H2@dW�B���|( Ӑ5C�(TLc�C�"��RZ3��T0 k� �K��O�%�@c  �e1t B  ��    �   �@<A H3@dW�B���|( ӌ6C�(TLc�D�"��RZ3��T0 k� �K��O�%�@c  �e1t B  ��    �   �@<A D3@dW�B���|( ӌ8C�(TLc�D�"��RZ3��T0 k� �K��O�%�@c  �e1t B  ��    �   �@<A D4@dW�B���|( ӌ9C�$TLc�D�#��SZ3��T0 k� �K��O�%�@c  �e1t B  ��    �   �@<@ D4@dW�B���|( ӌ:C�$TLc�D�#��SZ3��T0 k� �K��O�%�@c  �e1t B  ��    �   �@<@ D5@dW�B���|( ӌ:C�$TLc�E�#��SZ3��T0 k� �K��O�%�@c  �e1t B  ��    �   �@<@ @5@dW�B���|( ӈ;C�$TLc�E�#��SZ3��T0 k� �O��S�%�@c  �e1t B  ��    �   �@<@ @6@dW�B���|( ӈ<C�$TLc�E�#��SZ3��T0 k� �O��S�%�@c  �e1t B  ��   �   �@<@ @6@dW�B���|( �=C�$TLc�E�#��SZ3��T0 k� �O��S�%�@c  �e1t B  ��    �   �@<? <7@dW�B���|( �=D$TLc�E�#��SZ3��T0 k� �O��S�%�@c  �e1t B  ��    �   �@<? <7@dW�B���|( �>D$TLc�E�#��SZ3��T0 k� �O��S�%�@c  �e1t B  ��    �   �@<? <7@dW�B���|( �?D$TLc�E�$��SZ3��T0 k� �O��S�%�@c  �e1t B  ��    �   �@<? <8@dW�B���|( �@D$TLc�E�$��SZ3��T0 k� �O��S�%�@c  �e1t B  ��   �   �@<> 88@dW�B���|( �AD$TLc�E�$��SZ3��T0 k� �O��S�%�@c  �e1t B  ��   �   �@<> 89@dW�B���|( �AD$TLc�E�$��SZ3��T0 k� �O��S�%�@c  �e1t B  ��    �   �@<> 89@dW�B���|( �BD$TLc�E�$��SZ3��T0 k� �S��W�%�@c  �e1t B  ��   �   �@<> 8:@dW�B���|( �|CD$TLc�E�$��SZ3��T0 k� �S��W�%�@c  �e1t B  ��    �   �@<> 8:@dW�B���|( �|DD$TLc�E�$��SZ3��T0 k� �S��W�%�@c  �e1t B  ��    �   �@<= 4:@dW�B���|( �|ED$TLc�F�$��SZ3��T0 k� �S��W�%�@c  �e1t B  ��    �   �@<= 4;@dW�B���|( �|FD$ULc�F�$��SZ3��T0 k� �S��W�%�@c  �e1t B  ��    �   �@<= 4;@dW�B���|( �xGD$ULc�F�$��SZ3��T0 k� �S��W�%�@c  �e1t B  ��    �   �@8= 4;@dW�B���|( �xGD$ULc�F�$��SZ3��T0 k� �S��W�%�@c  �e1t B  ��    �   �@8= 0<@dW�B���|( �xHD$ULc�F�%��SZ3��T0 k� �S��W�%�@c  �e1t B  ��    �   �@8< 0<@dW�B���|( �xID$ULc�F�%��SZ3��T0 k� �S��W�%�@c  �e1t B  ��    �   �@8< 0=@dW�B���|( �tJD$ULc�F�%��SZ3��T0 k� �S��W�%�@c  �e1t B  ��    �   �@8< 0=@dW�B���|( �tKD$ULc�F�%��SZ3��T0 k� �S��W�%�@c  �e1t B  ��    �   �@8< 0=@dW�B���|( �tKD$ULc�F�%��SZ3��T0 k� �W��[�%�@c  �e1t B  ��    �   �@8< 0>@dW�B���|( �tLD$ULc�F�%��SZ3��T0 k� �W��[�%�@c  �e1t B  ��    �   �@8< ,>@dW�B���|( �pMD$ULc�F�%��SZ3��T0 k� �W��[�%�@c  �e1t B  ��    �   �@8; ,>@dW�B���|( �pMD$ULc�F�%��SZ3��T0 k� �W��[�%�@c  �e1t B  ��    �   �@8; ,?@dW�B���|( �pND$ULc�F�%��SZ3��T0 k� �W��[�%�@c  �e1t B  ��    �   �@8; ,?@dW�B���|( �pOC�$ULc�G�%��SZ3��T0 k� �W��[�%�@c  �e1t B  ��    �   �@8; ,?@dW�B���!�( �lPC�$ULc�G�%3�Sbs��T0 k� �W��[�%�@c  �e1t B  ��    �   �@8; (?@dW�B���!�( �lPC�$ULc�G�%3�Sbs��T0 k� �W��[�%�@c  �e1t B  ��    �   �@8; (@@dW�B���!�( �lQC� ULS�G�&3�Sbs��T0 k� �W��[�%�@c  �e1t B  ��    �   �@8; (@@dW�B���!�( �lRC� VLS�G�&3�Sbs��T0 k� �W��[�%�@c  �e1t B  ��    �   �@8: (@@dW�B���!�( �hRL VLS�G�&3�Sbs��T0 k� �[��_�%�@c  �e1t B  ��    �   �@8: (A@dW�B���!�( �hSL VLS�G�&3�Sbs��T0 k� �[��_�%�@c  �e1t B  ��    �   �@8: (A@dW�B���!�( �hSL VLS�G�&3�Sbs��T0 k� �[��_�%�@c  �e1t B  ��    �   �@8: $A@dW�B���!�( �hTL VLS�G�&3�Sbs��T0 k� �[��_�%�@c  �e1t B  ��    �   �@8: $B@dW�B���!�( �hUL VD��G�&3�Sbs��T0 k� �[��_�%�@c  �e1t B  ��    �   �@8: $B@dW�B���!�( �dULVD��G�&3�Sbs��T0 k� �[��_�%�@c  �e1t B  ��    �   �@8: $B@dW�B���!�( �dVLVD��G�&3�Sbs��T0 k� �[��_�%�@c  �e1t B  ��    �   �@89 $B@dW�B���|( �dVLVD��G�&3�SZ3��T0 k� �[��_�%�@c  �e1t B  ��    �   �@89 $C@dW�B���|( �dWLVD��G�&3�SZ3��T0 k� �[��_�%�@c  �e1t B  ��    �   �@89 $C@dW�B���|( �dWLVE�H�&3�SZ3��T0 k� �[��_�%�@c  �e1t B  ��    �   �@89  C@dW�B���|( �`XLWE�H�&C�SZ3��T0 k� �[��_�%�@c  �e1t B  ��    �   �@89  C@dW�B���|( �`YLWE�I�&C�SZ3��T0 k� �_��c�%�@c  �e1t B  ��    �   �@89  D@dW�B���|( �`YLWE�I�'C�SZ3��T0 k� �_��c�%�@c  �e1t B  ��    �   �@89  D@dW�B���|( �`ZL$WE�I�'C�TZ3��T0 k� �_��c�%�@c  �e1t B  ��    �   �@89  D@dW�B���|( �`ZL$WF�I�'C�TZ3��T0 k� �_��c�%�@c  �e1t B  ��    �   �@88  D@dW�B���|( �`[L$WF�I�'C�TZ3��T0 k� �_��c�%�@c  �e1t B  ��    �   �@88  E@dW�B���|( �\[L$WF�J�'C�TZ3��T0 k� �_��c�%�@c  �e1t B  ��    �   �@88 E@dW�B���|( �\\L$WF�K�'C�TZ3��T0 k� �_��c�%�@c  �e1t B  ��    �   �@88 E@dW�B���!�( �\\L$WF�K�'C�Tb���T0 k� �_��c�%�@c  �e1t B  ��    �   �@88 E@dW�B���!�( C\]L$WDӤL�'C�Tb���T0 k� �_��c�%�@c  �e1t B  ��    �   �@88 E@dW�B���!�( C\]L$WDӤL�'C�Ub���T0 k� �_��c�%�@c  �e1t B  ��    �   �@88 F@dW�B���!�( C\^L$WDӤM�'C�Ub���T0 k� �_��c�%�@c  �e1t B  ��    �   �@88 F@dW�B���!�( CX_L$XDӤM�'C�Ub���T0 k� �c��g�%�@c  �e1t B  ��    �   �@88 F@dW�B���!�( CX_L$XDӠM�'C�Ub���T0 k� �c��g�%�@c  �e1t B  ��    �   �@88 F@dW�B���!�( 3X`L$XF�N�'C�Ub���T0 k� �c��g�%�@c  �e1t B  ��    �   �@87 F@dW�B���!�( 3XaL$XF�N�'C�Ub���T0 k� �c��g�%�@c  �e1t B  ��    �   �@87 G@dW�B���!�( 3XbL$XF�N�'C�Vb���T0 k� �c��g�%�@c  �e1t B  ��    �   �@87 G@dW�B���!�( 3XcL$XF�N�'C�Vb���T0 k� �c��g�%�@c  �e1t B  ��    �   �@87 G@dW�B���!�( 3XdL$XF�O�'C�Vb���T0 k� �c��g�%�@c  �e1t B  ��    �   �@87 G@dW�B���|( #XeL$XE��O�'C�VZ3��T0 k� �c��g�%�@c  �e1t B  ��    �   �@87 G@dW�B���|( #XfL$XE��P�(C�WZ3��T0 k� �c��g�%�@c  �e1t B  ��    �   �@87 H@dW�B���|( #XgL$XE��P�(C�WZ3��T0 k� �c��g�%�@c  �e1t B  ��    �   �@87 H@dW�B���|( #\hL$YE��Q�(C�WZ3��T0 k� �c��g�%�@c  �e1t B  ��    �   �@87 H@dW�B���|( #\iL$YE��Q�(C�WZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@87 H@dW�B���|( \jL$YE#�Q�(C�WZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@87 H@dW�B���|( `kL$ YE#�Q�(C�XZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@86 H@dW�B���|( `lL$ YE#�R�(C�XZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@86 I@dW�B���|( dmL$ YE#�R�(C�XZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@86 I@dW�B���|( dnL$ YE#�S�(C�XZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@86 I@dW�B���|( hoL$ YE3�S�(C�XZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@86 I@dW�B���|( �loL$ YE3�T�(C�XZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@86 I@dW�B���|( �lpL$ YE3�U�(C�XZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@86 I@dW�B���|( �pqL$ ZE3�U�(C�XZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@86 J@dW�B���|( �trL$ ZE3�V�(C�XZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@86 J@dW�B���|( �xrL$ ZEC�W�(C�XZ3��T0 k� �g��k�%�@c  �e1t B  ��    �   �@86 J@dW�B���|( �|sL$ ZEC�X�(C�XZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@86 J@dW�B���|( ��sL$$ZEC�Y�(C�YZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@86 J@dW�B���|( ��tL$$ZEC�Z�(C�YZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@86 J@dW�B���|( ��tL$$ZEC�[�(C�YZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@86 J@dW�B���|( ��uL$$ZEC�\�(C�YZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@86 K@dW�B���|( ��uL$$ZEC�]�(C�YZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@85 K@dW�B���|( s�uL$$ZES�^�(3�ZZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@85 K@dW�B���|( s�uL$$ZES�^��(3�ZZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@85 K@dW�B���|( s�uL$$ZES�_��)3�ZZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@85 K@dW�B���|( s�uL$ZES�_��)3�ZZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@85 K@dW�B���|( s�uL$[ES�`��)3�ZZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@85 K@dW�B���|( s�uL$[EC�a��)3�ZZ3��T0 k� �k��o�%�@c  �e1t B  ��    �   �@85 L@dW�B���|( s�uL([EC�b��)3�ZZ3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 L@dW�B���|( s�uL([EC�c��)3�[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 L@dW�B���|( s�uL([EC�c��)3�[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 L@dW�B���|( ��tC�([EC�d��)3�[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 L@dW�B���|( ��tC�([EC�d��)��[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 L@dW�B���|( ��tC�([EC�d��)��[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 L@dW�B���|( ��tC�$[@��d��)��[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 L@dW�B���|( ��sC�$[@��d��)��[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 L@dW�B���|( ��sC�$[@��d��)��[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 M@dW�B���|( ��sC�$[@��c�)��[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 M@dW�B���|( ��rC�$[@��c�)��[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 M@dW�B���|( ��rC�$[@��c�)��[Z3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@85 M@dW�B���|( ��qC�$\@��c�)��ZZ3��T0 k� �o��s�%�@c  �e1t B  ��    �   �@84 M@dW�B���|( ��qC� \@��b�)��ZZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 M@dW�B���|( ��pC� \@��b�)��ZZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 M@dW�B���|( ��pC� \E#�b�)��ZZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 M@dW�B���|( ��oC� \E#�b�)��ZZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 M@dW�B���|( ��nC� \E#�b�)��ZZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( ��mC� \E#�b�)��ZZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( ��lC� \E#�b�)��ZZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( ��kC� \E#�b�)��ZZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( ��jC� \E�b�)��ZZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( ��jC� \E�b�)��ZZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( s�jC� ]E�b�)��YZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( s�jC� \E�b�)��YZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( s�jC� \E�b�)��YZ3��T0 k� �s��w�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( s�iD [B��a�)��XZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( s�iD [B��a�)��XZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( s�iD [B��a�*��XZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 N@dW�B���|( c�hD [B��a�*��XZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 O@dW�B���|( c�hD ZB��`�*��XZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 O@dW�B���|( c�gD ZK��`�*��XZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 O@dW�B���|( c�gD ZK��`�*��XZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 O@dW�B���|( c�gD ZK��`�*��XZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 O@dW�B���|( c�gD YK��`�*��WZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 O@dW�B���|( c�gD YK��_�*��WZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 O@dW�B���|( c�gD YK��_�*3�WZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 O@dW�B���|( c�fD YK��_�*3�WZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �@84 O@dW�B���|( c�fD YK��_�*3�WZ3��T0 k� �w��{�%�@c  �e1t B  ��    �   �D��8  , C��_8(/?�|( �+�E0(E�tQ�
��#Z3� T0 k� �{���%�@c  �e1t B  ��    �   DD��9�0 C��_8*/C�|( �+�E0(E�xQ�
��#Z3� T0 k� �t�x%�@c  �e1t B  ��    �   ED��:�4 C��_8+�C�|( �+�E0(F xQ� �#Z3� T0 k� �p�t%�@c  �e1t B  ��    �   FD��:�8 C��_8,�G�|( �+�E0(F |Q� �#Z3� T0 k� �l�p%�@c  �e1t B  $�    �   GD��;�<C��_8-�G�|( �+�E0(F �Q� �#Z3� T0 k� 0d
�h
%�@c  �e1t B  �    �   HD�=<C��_8/�K�|( �+�E0$F �a#� �#Z3� T0 k� 0h�l%�@c  �e1t B  ��    �   ID�>@ E��_80	?K�|( �+�E $F �a+� �$Z3� T0 k� 0d�h%�@c  �e1t B  ��    �   JD�>D E��_80	?K�|( �+�E $F �a/� �$Z3� T0 k� 0g��k�%�@c  �e1t B  ��    �   KD�?K�E��o81	?O�|( �+�E $F �a3� �$Z3� T0 k� �g��k�%�@c  �e1t B  ��    �   LD�AS�E��o83	?O�|( �/�E $
F �	a?� �%Z3� T0 k� �o��s�%�@c  �e1t B  ��    �   MD�B[�E�o84	OO�|( �/�E $	E��
aG� �%Z3� T0 k� �o��s�%�@c  �e1t B  ��    �   ND�C_�E�o84	OO�|( �/�E $E��aK� �%Z3� T0 k� �s��w�%�@c  �e1t B  ��    �   OD� Dg�E�o85	OO�|( �/�E (E��aS� �&Z3� T0 k� �w��{�%�@c  �e1t B  ��    �   PD�$Ek�E�o86	OS�|( �/�E (E��aW��&Z3� T0 k� �����%�@c  �e1t B  ��    �   QD�,Gw�E�o87	?S�|( �/�E (E��c��'Z3� T0 k� ������%�@c  �e1t B  ��    �   SE 0I{�B��o88	?S�|( 	�/�E,E��k��'Z3� T0 k� ������%�@c  �e1t B  ��    �   UE 8J��B��o88	?S�|( 	�/�E, E��o��(Z3� T0 k� ������%�@c  �e1t B  ��    �   WE <K���B��89	?W�|( 	�/�E3�E��w���(Z3� T0 k� ������%�@c  �e1t B  ��    �   YE @L���B�#�89	?W�|( 	�/�E3�E�����)Z3� T0 k� ������%�@c  �e1t B  ��    �   [E�LN���E�+�8;	OW�|( 	�/�E;�B������*Z3� T0 k� ������%�@c  �e1t B  ��    �   ]E�PO���E�3�8;	OW�|( 	�/�E;�B������*Z3� T0 k� ������%�@c  �e1t B  ��    �   _E�XP���E�7�8<	OT |( 	�/�E?�B������*Z3� T0 k� ������%�@c  �e1t B  ��    �   aE�\Q���E�;�8<	OX|( 	�/�EC�B������+Z3� T0 k� ������%�@c  �e1t B  ��    �   cE�`R���E�?�8=	OX|( 	�/�EG�B������+Z3� T0 k� ������%�@c  �e1t B  ��    �   eE�hS���E�C�8=	?X|( 	�/�EK�B����
��+Z3� T0 k� ������%�@c  �e1t B  ��    �   gB�tU���B�O�8>	?X|( 	�/�ES�B����
� ,Z3� T0 k� ������%�@c  �e1t B  ��    �   jB�|V���B�S�8?	?X|( 	�/�E�W�B���
�-Z3� T0 k� ������%�@c  �e1t B  ��    �   mB��W���B�[�8@	?X|( 	�/�E�[�B���
�-Z3� T0 k� ������%�@c  �e1t B  ��    �   pB��X���B�_�8@	O\|( 	�/�E�_�E���
�-Z3� T0 k� �����%�@c  �e1t B  ��    �   sB��Y���B�c�8A	O\|( 	�/�E�c�E���
�.Z3� T0 k� ����%�@c  �e1t B  ��    �   vI�Y���Ek�8A	O\|( 	�/�E�g�E� ��
�.Z3� T0 k� ����%�@c  �e1t B  ��    �   yI�[��Ew�8B	O\|( 	�/�E�s�E�0��
� /Z3� T0 k� ���#�%�@c  �e1t B  ��    �   |I�[��E{�8C	?\|( 	�/�E�w�E�8��
�$/Z3� T0 k� �'��+�%�@c  �e1t B  ��    �   I�\��E��8C	?\|( 	�/�E�{�E�@��
�(/Z3� T0 k� �3��7�%�@c  �e1t B  ��    �   �I �\�#�E��8C	?`	|( 	�/�E���E�H��00Z3� T0 k� �?��C�%�@c  �e1t B  ��    �   �I �]�+�B���8D	?`	|( 	�/�E���E�P��40Z3� T0 k� �G��K�%�@c  �e1t B  ��    �   �I �]�7�B���8D	?`
|( 	�/�E���E�X��80Z3� T0 k� �O��S�%�@c  �e1t B  ��    �   �I �^�G�B���8E	O`|( 	�/�E���E�h'��D1Z3� T0 k� �_��c�%�@c  �e1t B  ��    �   �I�^O�B���8F	O`|(  3�E���E�l�+��H1Z3� T0 k� �c��g�%�@c  �e1t B  ��    �   �I�_W�I��8F	O`|(  3�E���E�t�3��L1Z3� T0 k� �k��o�%�@c  �e1t B  ��    �   �I�__�I��8G	O`|(  3�E���E�|�;��P1Z3� T0 k� �s��w�%�@c  �e1t B  ��    �   �I�_g�I��8G	Od|(  3�DЯ�E���?��T1Z3� T0 k� �{���%�@c  �e1t B  ��    �   �I�_o�I��8G	?d|(  7�Dз�E���G��\0Z3� T0 k� ������%�@c  �e1t B  ��    �   �I �`{�Ií/8H	?d|( �7�Dл�E���K��`0Z3� T0 k� ������%�@c  �e1t B  ��    �   �I �`��I Ϭ/8I	?d|( �;�D���E���W��h0Z3� T0 k� ������%�@c  �e1t B  ��    �   �I �`��I Ӭ/8I	?h|( �?�D���E���[�l/Z3� T0 k� ������%�@c  �e1t B  ��    �   �I �`��I ׬/<J/h|( �?�D���B��_�p/Z3� T0 k� ������%�@c  �e1t B  ��    �   �B��` !��I ۬/<K/h|( �C�D���B��c�t/Z3� T0 k� ������%�@c  �e1t B  ��    �   �B��` !��I ߬/<K/l|( �G�D���B���k�|.Z3� T0 k� ������%�@c  �e1t B  ��    �   �B��` !��I�<L/l|( �K�D���B���o��.Z3� T0 k� ������%�@c  �e1t B  ��    �   �B��` !��I�@M/p|( �O�D���B���s��.Z3� T0 k� �����%�@c  �e1t B  ��    �   �B��` !��I�@Mp|( �O�D���B���w��-Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`���I�DNt|( �S�D���B���w��-Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`���I ��HOx|( �[�D��B�����,Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`���I ��HP||( �_�D��B������+Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`���I ���LP�||( �c�D��B������*Z3� T0 k� ���#�%�@c  �e1t B  ��    �   �B��`���I ���PQ��|( �k�D�#�B������*Z3� T0 k� �#��'�%�@c  �e1t B  ��    �   �B��`��I ���TQ��|( �o�D�+�E�R����)Z3� T0 k� �'��+�%�@c  �e1t B  ��    �   �B��` r�B����TR��|( �s�D�3�E�R����)Z3� T0 k� �/��3�%�@c  �e1t B  ��    �   �B��` r�B����XR��|( �w�D�;�E� R����(Z3� T0 k� �4�8%�@c  �e1t B  ��    �   �B� ` r#�B���`S��|( ��D�K�E�0R����'Z3� T0 k� �H�L%�@c  �e1t B  ��    �   �B�` r/�B���dT��|( ���D�S�E�8R����'Z3� T0 k� �P�T%�@c  �e1t B  ��    �   �B�` r7�B���hT��|( ���D�[�E�@R����&Z3� T0 k� �X�\%�@c  �e1t B  ��    �   �B�` r?�B���lU��|( ���D�c�E�HR����&Z3� T0 k� �`�d%�@c  �e1t B  ��    �   �B�` rG�B���pU��|( �D�k�E�PR����%Z3� T0 k� �h�l%�@c  �e1t B  ��    �   �B�` rO�B���tV��|(  ��D�s�E�XR����%Z3� T0 k� �p�t%�@c  �e1t B  ��    �   �B� ` rW�B���xV��|(  ��D�{�E�`R����$Z3� T0 k� �x	�|	%�@c  �e1t B  ��    �   �B�,` rW�B���W�|(  ��D��E�p%�����#Z3� T0 k� ��
��
%�@c  �e1t B  ��    �   �B�0`�[�B�#��X�|(  ��F��E�x%����#Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�8`�c�B�'��X�|( ��F��E��%����#Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�<`�g�B�+��Y�|( ��F��E��%����"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�D`�k�B�/��Y� |( ǐF��E��%����"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�L`�o�B�7��Z� |( ˑF��E��%���� "Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�P`�s�B�;���Z��!|( ӒF��E��%����$"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�``�{�B�C���[��"|( �F��PR�%����4"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�d`��B�K���[��"|( �F� PR�%����<"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�l`��B�O���[��"|( �F�PR�%����D"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�t`��B�S���[�"|( ���E��PR�%���	2H"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�|`��B�[���\�"|( ���E��PR�%���	2P"Z3� T0 k� ����%�@c  �e1t B  ��    �   �Bф`��B�_���\�"|( ��E��PR�%���	2X"Z3� T0 k� ����%�@c  �e1t B  ��    �   �Bь`��B�g���\�#|( ��E��Pb�%���	2\"Z3� T0 k� ����%�@c  �e1t B  ��    �   �Bє`��B�k���\�#|( ��E��Pb�%���	2d"Z3� T0 k� ����%�@c  �e1t B  ��    �   �Bќ`��B�s���\�$#|( ��E�Pb�%���	2h"Z3� T0 k� ����%�@c  �e1t B  ��    �   �BѬ`��B����\�4"|( �3�E�Pb�%���	Bt"Z3� T0 k� ����%�@c  �e1t B  ��    �   �BѴ`��B�����\�<"|( �;�E�	Pb�%���	Bx"Z3� T0 k� ����%�@c  �e1t B  ��    �   �BѼ`��B���� [�@"|( �C�E�$
Pb�%���	B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`��B����[�H"|( �K�E�,
Pb�
%���	B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`��B����[�P"|( �W�E�4Pc 
%���	B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`��Bџ��[�X!|( �_�E�<PS	%���2�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`��Bѧ��Z�`!|( �g�E�DPS%���2�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`��Bѯ�� Z�h!|( �s�E�LPS%���2�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`��Bѷ��(Z�p |( �{�E�TPS%���2�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��`��B�ì�8Y�||( �{�E�dPS %��B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�`��B�ˬ�@X��|( ���E�lE�$%��B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�`���B�׬�DX��|( ���E�tE�(%��B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�`���B�߬�LW��|( ���E�|E�,%��B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�`���B���TW��|( ���E��E�0%��B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�$`���B���\V�|( ���E��E�4%��B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�,`���B����dU��|( ���E��IS8%��B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�4`���B����lU��|( ���E��IS<%��B�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�D`���B���xS��|( �ǦE��ISD%��2�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�L`���B����S��|( �ϦE��ISH %��2�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�T`���B����R��|( צE��E�O�%��2�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�\`���B�'��R��|( �E��E�S�%��2�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�h`���B�3��Q��|( �E��E�W��#�2�"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B�p`���B�;��Pp�|( �E��E�[��#���"Z3� T0 k� ����%�@c  �e1t B  ��    �   �B��` r��B�K��Oq |( �E��PSc��'���"Z3� T0 k� � �%�@c  �e1t B  ��    �   �B��` r��B�S���Nq|( �E��PSg��'���"Z3� T0 k� ��%�@c  �e1t B  ��    �   �B` r��B�[���Mq|( �E��PSk��'���#Z3� T0 k� ��%�@c  �e1t B  ��    �   �B` r��B�c���Mq|( �#�E��PSo��'���#Z3� T0 k� ��%�@c  �e1t B  ��    �   �B ` r��B�k���Lq |( �#�E��PSs��+���#Z3� T0 k� ��%�@c  �e1t B  ��    �   �B°`��B�{���Jq,|( �3�E�Pc{��+���$Z3� T0 k� �	�	%�@c  �e1t B  �    �   �@�`��E�����Jq4|( �?�E�Pc��+�"�%Z3� T0 k� ��%�@c  �e1t B  �    �   �@�`��E�����I�<|( G�E�Pc��c+�# %Z3� T0 k� � � %�@c  �e1t B  �    �   �@�`��E�����H�H|( W�E� Pc��c+�#&Z3� T0 k� 3�%�@c  �e1t B  ��    �   �@�`�E���@�G�P|( c�Ps$Pc��c+�#'Z3� T0 k� 3�%�@c  �e1t B  ��    �   �@�`�E���A F�X|( k�Ps(PS��c+�#(Z3� T0 k� 3�%�@c  �e1t B  ��    �   �@�`��E���AE�`|( �w�Ps,PS��S'�#(Z3� T0 k� 3�%�@c  �e1t B  ��    �   �@�`��E���AE�d|( ��Ps4PS��S'�#)Z3� T0 k� 3���%�@c  �e1t B  ��    �   �@�`��E�ǰAD�l|( ���Ps8PS��S'�#*Z3� T0 k� ����%�@c  �e1t B  ��    �   �@�`��@bϰAC�p|( ���Ps<PS��S'�# *Z3� T0 k� ����%�@c  �e1t B  ��    �   �@`�@b߰A$B� |( ���P�D
PS��S#��(,Z3� T0 k� ����%�@c  �e1t B  ��    �   �@`�@b�A,B��|( ���P�H
PS��c��0-Z3� T0 k� ������%�@c  �e1t B  �    �   �@`#�@b�A0A��|( ���P�P
PS��c��4-Z3� T0 k� ������%�@c  �e1t B  �    �   �@`'�@b��A8@��|( ���P�T	PS��c��8.Z3� T0 k� ������%�@c  �e1t B ��    �   �@$`+�@b��A<@��|( ���P�X	PS��c��</Z3� T0 k� ������%�@c  �e1t B ��    �   �@,`+�@c�AD?��|( ���P�\	PS��c��@0Z3� T0 k� ������%�@c  �e1t B ��    �   �@0`/�@c�AH?��|( �ǩP�`	A�����H1Z3� T0 k� ������%�@c  �e1t B ��    �   �@8`3�@c�AL>��|( �ϪP�d	A�����L2Z3� T0 k� ������%�@c  �e1t B ��   �   �@<`7�@c�AT=��|( �۪PshA�����P3Z3� T0 k� ������%�@c  �e1t B ��    �   �@D`;�@c#�AX=��|( ��PslA�����T4Z3� T0 k� �{���%�@c  �e1t B ��    �   �@H`#?�@c+�A\<��|( ��PstA�����\5Z3� T0 k� �k��o�%�@c  �e1t B ��    �   �@P`#C�@c3�Ad<��|( ���PsxEӷ����`6Z3� T0 k� �[��_�%�@c  �e1t B ��    �   �@\`#K�@c?�Al;���|( ���Ps�Eӷ���l8Z3� T0 k� �;��?�%�@c  �e1t B
 ��    �   �@``#O�@cG�Ap:���|( ���EÄEӷ���p9Z3� T0 k� �+��/�%�@c  �e1t B
 ��    �   �@d`#S�@cO�Ax:���|( ��EÄEӷ���t:Z3� T0 k� ����%�@c  �e1t B ��    �   �@l`#W�@cW�A|9���|( ��EÈA�����|;Z3� T0 k� ����%�@c  �e1t B ��    �   �@p`3[�@c_�A�9���|( ��EÌA������<Z3� T0 k� ������%�@c  �e1t B ��    �   �@x`3_�@cg�A�8���|( ��EÐA������=Z3� T0 k� ������%�@c  �e1t B �    �   �@|`3_�@co�A�8���|( �'�EӐA�������?Z3� T0 k� 1�����%�@c  �e1t B ��    �   �@�`3_�@cw�A�7���|( C/�EӔA�������@Z3� T0 k� 1�����%�@c  �e1t B ��    �   �@�`3c�@c�A�7���|( C7�EӘLS������AZ3� T0 k� 1�����%�@c  �e1t B ��    �   �@�`3g�@c��A�6���|( CC�EӘLS������CZ3� T0 k� 1�����%�@c  �e1t B ��    �   �@�`3k�@c��A�5���|( CK�E�LS�����	3�EZ3� T0 k� ������%�@c  �e1t B ��    �   �@�`3k�@c��A�5��|( CS�E�LS�����	3�FZ3� T0 k� ������%�@c  �e1t B ��    �   �@�`3k�@c��A�5��!�( CW�E�LS�����	3�Gb�� T0 k� ������%�@c  �e1t B ��   �   �@�`3o�@c��A�4��!�( C_�E�LS�����	3�Hb�� T0 k� ������%�@c  �e1t B ��    �   �@�`3s�@c��A�4��!�( Cg�E�LS�����	3�Ib�� T0 k� ������%�@c  �e1t B ��    �   �@�`3s�@c��A�3��!�( Ck�A��LS�����	3�Jb�� T0 k� !�����%�@c  �e1t B ��    �   �@�`3w�@c��A�3��!�( Cs�A��LS�����	C�Jb�� T0 k� !�����%�@c  �e1t B ��    �   �@�`3w�@c��A�2��!�( Cw�A��LS�����	C�Kb���T0 k� !�����%�@c  �e1t B
 ��    �   �@�`3{�@cǸA�2�#�!�( S�A��LS�����	C�Lb���T0 k� !�����%�@c  �e1t B
 ��    �   �@�`3{�@c˸A�2�'�!�( S��A��	LS�����	C�Mb���T0 k� !�����%�@c  �e1t B	 ��    �   �@�`3�@cӸA�1�+�!�( S��A�
Lc�����	C�Mb���T0 k� A�����%�@c  �e1t B	 ��    �   �@�`3�@c׹A�1�/�!�( S��A�
Lc��R��	3�Nb���T0 k� A�����%�@c  �e1t B	 ��    �   �@�`3��@c�A�0�3�!�( S��A�Lc��R��	3�Ob���T0 k� A�����%�@c  �e1t B ��    �   �@�`3��@c�A�0�7�|( S��A�Lc��R��	3�OZ3��T0 k� A�����%�@c  �e1t B ��    �   �@�`3��@c�A�/�;�|( S��D��Lc��R��	3�PZ3��T0 k� !�����%�@c  �e1t B ��    �   �@�`3��@c��A�/�?�|( S��D��Lc��R��	C�PZ3��T0 k� !�����%�@c  �e1t B ��    �   �@�`3��@c��A�/�C�|( S��D��Lc��B��	C�PZ3��T0 k� !�����%�@c  �e1t B ��    �   �@�a3��@c��A�.�G�|( S��D��Lc��B��	C�PZ3��T0 k� !�����%�@c  �e1t B ��    �   �@�a3��@d�A�.�K�|( c��D��Lc��B��	C�PZ3��T0 k� !�����%�@c  �e1t B ��    �   �@�a3��@d�A�.�O�|( c��D��Lc��B��	C�PZ3��T0 k� ������%�@c  �e1t B ��    �   �@�a3��@d�A�-�O�|( c��D��Lc��B��	3�PZ3��T0 k� ������%�@c  �e1t B ��    �   �@�a3��@d�A�-�S�|( c��D��Lc�����	3�PZ3��T0 k� ������%�@c  �e1t B ��    �   �@�a3��@d�A�-�W�|( c��D��Lc�����	3�PZ3��T0 k� ������%�@c  �e1t B ��    �   �@�b3��@d#�A�,�_�|( ���D��Lc�����	3�PZ3��T0 k� ������%�@c  �e1t B  ,�    �   �@�b3��@d'�A�,�_�!�( ���D��Lc��ҿ�	C�Pbs��T0 k� ������%�@c  �e1t B  ��    �   �@ b3��@d+�A�,�c�!�( ���D��Lc��һ�	C�Pbs��T0 k� !�����%�@c  �e1t B  ��    �   �@b3��@d3�B +�g�!�( ���D��Lc��ҷ�	C�Pbs��T0 k� !�����%�@c  �e1t B ��    �   �@b3��@d7�B+�k�!�( ���D��Lc��ү�	C�Pbs��T0 k� !����%�@c  �e1t B ��    �   �@c3��@d;�B+�k�!�( ���D��Lc��ҫ�	C�Pbs��T0 k� !����%�@c  �e1t B ��    �   �@c3��@d?�B*�k�!�( ���D��!Lc����	3�Pbs��T0 k� !����%�@c  �e1t B ��    �   �@c3��@dC�B*�k�!�( ���D��#Lc����	3�Pbs��T0 k� �����%�@c  �e1t B ��    �   �@c3��@dG�B*�g�!�( ���D��$Lc����	3�Pbs��T0 k� �����%�@c  �e1t B ��    �   �@c3��@dK�B*�g�!�( ���D��&Lc����	3�Pbs��T0 k� �����%�@c  �e1t B ��   �   �@c3��@dO�B)�g�!�( ��D��(Lc����	3�Pbs��T0 k� �����%�@c  �e1t B ��    �   �@c3��@dS�B)�c�!�( ��D��*Lc��«� ��Pbs��T0 k� ����%�@c  �e1t B ��    �   �@ d3��@dW�B)�_�|( ��D��+Lc��§� ��PZ3��T0 k� ����%�@c  �e1t B ��    �   �@ d3��@d[�B)�[�|( ��D��-Lc��£� ��PZ3��T0 k� ����%�@c  �e1t B ��    �   �@$d3��@d_�B(�W�|( ��E�/Lc��� ��PZ3��T0 k� "���%�@c  �e1t B ��   �   �@(d3��@dc�B (�S�|( 4�E�1Lc��� ��PZ3��T0 k� "���%�@c  �e1t B ��    �   �@(d3��@dg�B$(�S�|( 4�E�3Lc��� ��PZ3��T0 k� "���%�@c  �e1t B ��    �   �@,d3��@dk�B$(�O�|( 4�E�5Lc��� ��PZ3��T0 k� "���%�@c  �e1t B ��    �   �@0d3��@do�B('�K�|( 4�E�7Lc��� ��PZ3��T0 k� "���%�@c  �e1t B ��    �   �@0d3��@ds�B('�G�|( 4�E�9Lc��� ��PZ3��T0 k� ����%�@c  �e1t B ��    �   �@,d3��@dw�B,'�C�|( ��E�;Lc��� ��PZ3��T0 k� ����%�@c  �e1t B ��    �   �@,c3��@d{�B,'�C�|( ��F�=Lc��� ��PZ3��T0 k� ����%�@c  �e1t B ��    �   �@,c3��@d�B0&�?�|( ��F�?Lc�����PZ3��T0 k� ����%�@c  �e1t B ��    �   �@,c3��@d�B0&�;�|( ��F�ALc�����PZ3��T0 k� ����%�@c  �e1t B ��    �   �@,b3��@d��B4&�;�|( ��F�DLc������PZ3��T0 k� ����%�@c  �e1t B ��   �   �@,b3��@d��B4&�7�|( ��F�FLc������PZ3��T0 k� ����%�@c  �e1t B ��    �   �@,b3��@d��B8&�3�|( ��F�HLS���{���PZ3��T0 k� "���%�@c  �e1t B ��    �   �@,b3��@d��B8%�/�|( ��F�JLS���w���PZ3��T0 k� "���%�@c  �e1t B ��    �   �@,a3��@d��B<%�/�|( ��F�LLS���w���PZ3��T0 k� "���%�@c  �e1t B  ��    �   �@,a3��@d��B<%�+�|( ��F�NLS���s���PZ3��T0 k� "���%�@c  �e1t B  ��    �   �@,a3��@d��B@%�+�|( ��F�PLS���o���PZ3��T0 k� "���%�@c  �e1t B  ��    �   �@(a3��@d��B@%�'�|( ��F�RLS���o���PZ3��T0 k� ����%�@c  �e1t B  .�    �   �@(`3��@d��BD$�#�|( ��F�UD����k���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@(`3��@d�BD$�#�|( ��F�WD����g���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@(`3��@d�BH$��|( ��E��YD����g���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@(`3��@d�BH$��|( ��E��[D����c���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@(_3��@d�BL$��|( ��E��]D����c���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@(_3��@d�BL$��|( ��E��_D���_���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@(_3��@d�BL#��|( ��E��aD���[���PZ3��T0 k� ����%�@c  �e1t B  ��   �   �@(_3��@d{�BP#��|( ���E��cD���[���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@(^3��@d{�BP#��|( ���E��eD���W���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@(^3��@d{�BT#��|( ���E��fD���W���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@(^3��@d{�BT#��|( ���E��hD���S���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$^3��@d{�BT#��|( ���E��jD���S���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@d{�BX"��|( ���E��lD���O���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@dw�BX"��|( ���E��mD���O���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@dw�B\"��|( ���E��oD���K���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@dw�B\"��|( ���E��qD���K���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@dw�B\"���|( ���E��rD���G���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@dw�B`"���|( ���E��tD���G���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@dw�B`"���|( ���E��uD���C���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@ds�B`!���|( ���E��vD���C���PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@ds�Bd!���|( ���E��wD���< ��PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@ds�Bd!���|( ���E��yD���<��PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@ds�Bd!���|( ���E��zD���8��PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@ds�Bh!���|( ���E�{D���8��PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@ds�Bh!���|( ���E�zD���8��PZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3��@ds�Bh!���|( ���E�yD���4��OZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$]3� @do�Bl!���|( ���E�yD���4��OZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$\3� @do�Bl ���|( ���E�xD���0��OZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$\3�@do�Bl ���|( ���E�wEc��0��OZ3��T0 k� ����%�@c  �e1t B  ��    �   �@$\3�@do�Bl ���|( ���E�vEc��0��OZ4�T0 k� ����%�@c  �e1t B  ��    �   �@$\3�@do�Bp ���|( ���E�uEc��,��OZ4�T0 k� ����%�@c  �e1t B  ��    �   �@$\3�@do�Bp ���|( ���E�tEc��,��OZ4�T0 k� ���#�%�@c  �e1t B  ��    �   �@$\3�@do�Bp ���|( ���E�sEc��(��OZ4�T0 k� ���#�%�@c  �e1t B  ��    �   �@$\3�@do�Bt ���|( ���E�rEc��(��OZ4�T0 k� ���#�%�@c  �e1t B  ��    �   �@$\3�@do�Bt ���|( ���E�qEc��(��OZ4�T0 k� ���#�%�@c  �e1t B  ��    �   �@$\3�@dk�Bt ���|( ���E�oEc��$	��OZ4�T0 k� ���#�%�@c  �e1t B  ��    �   �@$\3�@dk�Bt���|( ���E�nEc��$	��OZ4�T0 k� ���#�%�@c  �e1t B  ��    �   �@$\C�@dk�Bx���|( ���E� mD3��$
��OZ4�T0 k� ���#�%�@c  �e1t B  ��    �   �@$\C�@dk�Bx���|( ���E� lD3�� 
��OZ4�T0 k� ���#�%�@c  �e1t B  ��    �   �@$[C�@dk�Bx���|( ���E� lD3�� ��OZ4�T0 k� �#��'�%�@c  �e1t B  ��    �   �@$[C�@dk�Bx���|( ���K� kD3�� ��OZ4�T0 k� �#��'�%�@c  �e1t B  ��   �   �@$[C�@dk�B|���|( ���K� kD3����OZ4�T0 k� �#��'�%�@c  �e1t B  ��    �   �@$[C�	@dk�B|���|( ���K� kLS����NZ4�T0 k� �#��'�%�@c  �e1t B  ��    �   �@$ZC�	@dk�B|���|( ���K� kLS�����NZ4�T0 k� �#��'�%�@c  �e1t B  ��    �   �@$ZC�
@dg�B|���|( ���K�$jLS�����NZ4�T0 k� �#��'�%�@c  �e1t B  ��    �   �@(YC�@dg�B����|( ���K�$jLS�����NZ4�T0 k� �#��'�%�@c  �e1t B  ��    �   �@(Y�@dg�B����|( ���K�$iLS�����NZ4�T0 k� �#��'�%�@c  �e1t B  ��    �   �@(Y�@dg�B����|( ���K�(iLS�����NZ4�T0 k� �'��+�%�@c  �e1t B  ��    �   �@(X�@dg�B����|( C��K�(iLS� ���NZ4�T0 k� �'��+�%�@c  �e1t B  ��    �   �@(X�@dg�B����|( C��K�(hLS����NZ4�T0 k� �'��+�%�@c  �e1t B  ��    �   �@(W�@dg�B����|( C��L,hLS����MZ4�T0 k� �'��+�%�@c  �e1t B  ��    �   �@(W�@dg�B����|( C��L,gLS����MZ4�T0 k� �'��+�%�@c  �e1t B  ��    �   �@(V�@dg�B����|( C��L,gLS��C�MZ4�T0 k� �'��+�%�@c  �e1t B  ��    �   �@,V�@dg�B����|( ���L0fLS��C�MZ4�T0 k� �'��+�%�@c  �e1t B  ��    �   �@,U �@dg�B����|( ���L0fLS��C�MZ4�T0 k� �+��/�%�@c  �e1t B  ��    �   �@,U �@dc�B����|( ���L0eLc��C�NZ4�T0 k� �+��/�%�@c  �e1t B  ��    �   �@,T �@dc�B����|( ���L4eLc�C�NZ4�T0 k� �+��/�%�@c  �e1t B  ��    �   �@,T �@dc�B����|( ���L4eLc�C�NZ4�T0 k� �+��/�%�@c  �e1t B  ��    �   �@,T �@dc�B����|( ���L4dLc�C�NZ4�T0 k� �+��/�%�@c  �e1t B  ��    �   �@,T �@dc�B����|( ���L8dLc�C�OZ4�T0 k� �+��/�%�@c  �e1t B  ��    �   �@,T �@dc�B����|( ���L8dLc�	C�OZ4�T0 k� �+��/�%�@c  �e1t B  ��    �   �@,T �@dc�B����|( ���L8cLc�
C�OZ4�T0 k� �+��/�%�@c  �e1t B  ��   �   �@0S �@dc�B����|( ���L8cLc�
C�PZ4�T0 k� �/��3�%�@c  �e1t B  ��    �   �@0S �@dc�B�q��|( C��L<cLc�S�PZ4�T0 k� �/��3�%�@c  �e1t B  ��    �   �@0S �@dc�B�q��|( C��L<bLc�S�QZ4�T0 k� �/��3�%�@c  �e1t B  ��    �   �@0R �@dc�B�q��|( C��L<bLc�S�QZ4�T0 k� �/��3�%�@c  �e1t B  ��    �   �@0R �@dc�B�q��|( C��L<bLc� S�QZ4�T0 k� �/��3�%�@c  �e1t B  ��    �   �@0R �@dc�B�q��|( C��L@aLc� S�RZ4�T0 k� �/��3�%�@c  �e1t B  ��    �   �@0Q �@dc�B�q��|( 3��L@aLc� S�RZ4�T0 k� �/��3�%�@c  �e1t B  ��    �   �@0Q |@d_�B�q��|( 3��L@aLc� S�RZ4�T0 k� �/��3�%�@c  �e1t B  ��    �   �@0Q |@d_�B�q��|( 3��L@`Lc� S�RZ4�T0 k� �3��7�%�@c  �e1t B  ��    �   �@4Q |@d_�B�q��|( 3��LD`Lc��S�RZ4�T0 k� �3��7�%�@c  �e1t B  ��   �   �@4P |@d_�B���|( 3��LD`Lc��S�RZ4�T0 k� �3��7�%�@c  �e1t B  ��    �   �@4P |@d_�B���|( C��LD_Lc��S�RZ4�T0 k� �3��7�%�@c  �e1t B  ��    �   �@4P |@d_�B���|( C��LD_Lc��c�RZ4�T0 k� �3��7�%�@c  �e1t B  ��    �   �@4O x@d_�B���|( C��LH_Lc��c�RZ4�T0 k� �3��7�%�@c  �e1t B  ��    �   �@4O x@d_�B���|( C��LH_Lc��c�RZ4�T0 k� �3��7�%�@c  �e1t B  ��    �   �@4O x@d_�B���|( C��LH^Lc��c�RZ4�T0 k� �3��7�%�@c  �e1t B  ��    �   �@4O x@d_�B���|( C��LH^Lc��c�RZ4�T0 k� �3��7�%�@c  �e1t B  ��    �   �@4N x@d_�B���|( C��LH^Lc���RZ4�T0 k� �7��;�%�@c  �e1t B  ��    �   �                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��D� ]�&�&� � �� 4#�          �۝     4*�۝    ��               
   l �           ��     ���   0	%           O��          � ¹�     O� ���    ��                  �           %0     ���   0
 
         ��v       �    ��u+�                      l �         �     ���   8
           �K   $ $     �|M     �K �x�       3               A��          }P     ���   8         ���h         . c(�    ���h c)V      ��   	            ��          �`     ���   P	           �p  ��	      B�
+�      �p�
+�                              ���              �  ���    P              f�R  V V
    V ��     f�v ��    ��                	 Z �          �b     ��@  8�          Y%� A A 	   j��     YR3��    �d�0               ' Z �         �p�    ��@  (
 
           _k� � �
     ~ ��u     _� ���    ��D                Z �          + �     ��`   8

            *E�  � �    � t�Z     *?g t�     ]��               6 Z �         	 � �  
  ��h   (
            WS�  � �
   � �-b     Ws� �1�    � ��                	 Z �         
 �0�   
  ��`  P
B         ��ȓ��     � ��    ��ȓ �g      ��                      ����             �  ��@    8		 1                   ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��\�  ��        � �ܸ    ��{x ���    �4 "                  x                j  �   �	   �                         ��    ��        � �      ��   �           "                                                �                          � � c�
 � � t � ��� � �           
 	     
   �    �p ��G       &� `m@ 'd n  '� n  �� v  �  v@ &� n  0 k� $� �m@ %� n@ �� v  �  v@ �D n� �d n����J ����X ����X � 
�\ W� (D  q  � u� 
�\ W� �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� �R� � }` 
�\ V� 
� V� 
�\ W ���� � $ `m@ � n   n  �$ �r@ �$ s@ �D s` �d s� Є s� Ф s� �� 0o� �$ `p  �� p� � q  �$ q  �D q@ �� �t� �� u� � u� �$ v  �D v  �d v@ k @`� k� `a@ lD b  ld b  l� b@���� � 
�� W� 
�| W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� �   ���  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    B�j l �  B �
� �  �  
� ����  ��     � �  �    O��  ��     � �       *��  ��     � t          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �      �� � �  ���        �*T ��        �        ��        �        ��        �  	  ��    �n;����        ��                         T�) ,   ��                                     �                  ����           �� x���%��     � 2                 8 Geoff Sanderson y   0:01                                                                        2  2      �C
�Uc� =c� u c�&T c�0D � �C � �C/ 	C"	
B�H �	k~R �k�X �k�X �k� � �k� � �k� � k� � �c�O �c�G � c�G � c�T �c�B �	cVS �c\[ � c`S �kjO � kpG � kqQ �	� � �	� � �� � � � �!J�+ �"K � �#K �1$"�?1 %"�Q!&"�?!'*�N("� )"�,o*�o+
�) � ,!� � � -"H � �." � �/" x0"0 �1*P � 2)�` �  *Hx �  *K� �  *O� �  *R� �7*40 � 8*NP �  *R� �  *R� �  *H� �  *K� x=*$8 x>* P �  *O�
 
�* A"�4
B�
 
�-                                                                                                                                                                                         �� P @       �     @ 
        �     W P E X  ��        	           	 �������������������������������������� ���������	�
��������                                                                                          ��    ��~�q� ��������������������������������������������������������   �4, =  @y���q��%                                                                                                                                                                                                                                                                                                                                                        @f�@�                                                                                                                                                                                                                                              �        � �  D�J    	  E                             ������������������������������������������������������                                                                                                                                           �      �      �                �  �          	  
 	 
 	 	  ��� �� �����������  �������� ���� �������� ��������������������������� ������������������� �������������� �������������������������� ����������   � ������� ������������ �������������������  ��������������������������� ����������������             &                      �    2     �  L�J      
�                             ������������������������������������������������������                                                                                                                                            �    ��      �                ��            	     	 	 ������ ������ � ���� �������� � ���� �������������� ��������������������������������������������������������������� ��������������������������������������������� ��  �������������� �������� �������� �������� ������������ ������ ��� ���������             &                                                                                                                                                                                                                                                                                                               �             


            �   }�         ����������������   1������������    ����������������   '����������������  '�����������������������������                                                          'u                     ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" R > / 	              	                  � \&� �m@                                                                                                                                                                                                                                                                                     	n)n1n  �                a      e      e                        m                                                                                                                                                                                                                                                                                                                                                                                                                  �  >�  J�  (�  (�  Cm�  �̎����� ������8����
����B���˦�������                 ����  � {
        	 �   &  AG� �   h                    �                                                                                                                                                                                                                                                                                                                                      p B I   �        -             !��                                                                                                                                                                                                                            Y   �� �~ ���      �� B 	      ��� �� �����������  �������� ���� �������� ��������������������������� ������������������� �������������� �������������������������� ����������   � ������� ������������ �������������������  ��������������������������� ���������������������� ������ � ���� �������� � ���� �������������� ��������������������������������������������������������������� ��������������������������������������������� ��  �������������� �������� �������� �������� ������������ ������ ��� ���������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     :      9   � ��                       B     �   �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$     `d  �`���6 ��  �`���6 �$ ^$ �d`  �`  �d`   � 
�8 ��   � 
  @     �T w ���5�������� J�Q  @ 
in   ���� ��      m@ &� �� m@ &� �$ O&  ��O &      �  ��   )���� e�����   g���   �     f ^�         ��         )      ��D����2�������J��[���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            "! "   "      ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "! ""! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       "! "   "      ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �    �  �   �   �   �  �         �  �   �   ��  �              ��  �           �   �   �                                                  �               �  �  ��  �   �   �           �     �                   ���������������������  ��  ��  ��  �   �    �          �         �                                                                                              �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   �                         ��  �                             �  �   �   �   �   �  �   ��  ��       �  ��  ��  �   �   �    �  ��  ��  �                    � �� ��  �� ��  �  �  �   �                                                                                                                                                                                                    	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                        ��  ��  �                            �   �    �   �       �   �   �                .      �  �  ��  �   �   �        �   ��  ��  ��  �  �   ��  ��                                                                                                                                                                      �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   �   � �  ��" � �� "��  �                     �   �                                                            �               �  �  ��  �   �   �        ��  �  �  �   �                                                                                                                                                                             �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        ��                          ��  ��  ��  }�  ��  vw� wz� ��� �����        "  ""  ""/ �"� ��          �   �  � �� ��  �                        �   ��  �   ��  ��  �  �  �   �                                 �   ���                            �   �                                                                                                         �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                                                �   �   �  �  �  �  ���������  �U4"+�B�*�����"/���  ��� �� �  � �     �               ۲  �!  "  �� �� �  ��� ��  �� �                          	ʐ ��� ��� ڝ��ݩ��ݩ��ݩ��ک�̪��̪��̪������̽� ��� ��T �C                �   �   ��  ��  ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����            �  �  ��  �   �   �       ���                                                                                                                                                                                              � ���	�˽
ɷw�kk�gg��y ��� "-� �  8  ��  C> D4 D4  3�  ��  �$  ") "  "� �   �       �   �   ٰ  ��  ��  ��  ��  ٩  ��  ��  J�  [�  �  .0  ".  C�� T0�EP �   "   "   ��� �   �   �                        ��  ��                                �  �� �  �  �   �     ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                        � ��                  �  �˰ ��� �wp ���                                                                                                                                                                                     "  "(��ȩ�ܚ��ۊ����� ��  �   �   �   �   �� ��� ̻� ˽� ��� �w� �������������������������� �̻ ���         �   �       �   �   "" �+� Ȼ� ɫ� ɨ� ��                �� �I��3 ��D 
UD 
UD TD  T�  ˸  ��  �� ̰ �+ ��"/ �"/  ����  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �                �������  ���    �                      "  .���"    �     �                                                                                                                                                                                    "  " �" ��" ��- �ۼ w۽��ݹ����� ��� ��  ˼  ��  ˼  ��  H�  �D  J�  J�  �  �  �  �  
�  �  �  �  ,�  " "" �" �"�   ˰  ��  wp ��ډ�v���r�̸��˰��� ��  ��  ��  ��  ̸  ��  ��  DC  C4@ T4@ T40 T30 T30 S;� H�  ��  ��  ��  ""  "  �""� "�/��        �   �   �      �  �   �   �   �   �              �   �   �   �             ���� �                        " "" """ �"  �   �   �                              � ��                  �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                   �w
���̩ۚ,���+��   �   �   �   �  �  9  D3  D2 T2 DB DB �@ ��  ��  ��  �  "" ""�"!��" ��       �                w�  ��� ��� ��� ˼����ɀ�؊�˽ـ��˰��̰�̻@"���"+H�"$X�"$�@"E� U� E� D� ,˸  ��  ��  ,� "" �"" """�"!���� � �              �         �           �       �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                ���                                                                                                                                                                                                                     �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �               � � ����� ��                                                                                                                                                                                               �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��           	 
          
        ((((((( 
	(((( ����������������             ! " # $ % & '   ( $ % ) ! " # * ('(&(%($(#("(! (((���������������� + , -   . / 0 1  	 2         3       4 (((((((2	10/(.(-(,(+���������������� 5 6   7   8 9 1 :   $ % ) ! " #   ; ) ! " # $ % ) (#("(!()(%($ :198(((7(6(5����������������    <     = 8 0 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>108(=((( (<���������������� L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L����������������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7����������������  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(������������������D" � j  "  B   J jF� ����
��� �����
���� ����
��� �����
��� 0 q����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
�Uc� =c� u c�&T c�0D � �C � �C/ 	C"	
B�H �	k~R �k�X �k�X �k� � �k� � �k� � k� � �c�O �c�G � c�G � c�T �c�B �	cVS �c\[ � c`S �kjO � kpG � kqQ �	� � �	� � �� � � � �!J�+ �"K � �#K �1$"�?1 %"�Q!&"�?!'*�N("� )"�,o*�o+
�) � ,!� � � -"H � �." � �/" x0"0 �1*P � 2)�` �  *Hx �  *K� �  *O� �  *R� �7*40 � 8*NP �  *R� �  *R� �  *H� �  *K� x=*$8 x>* P �  *O�3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������B�[�X�O��5�N�S�_�R�K�\� � � � � � � � �,�>�0�����������������������������������������!��9�G�Z��6�G�0�U�T�Z�G�O�T�K� � � � � � �,�>�0�����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $������������������������     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %������������������������ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 