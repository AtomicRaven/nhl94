GST@�                                                            \     �                                               � ���      �  �           ����e ����ʲ������������������        �g      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    "�j* ,  �����
�"     �j@ �    ��
  �                                                                              ����������������������������������       ��    a= bQ0 4 411 c  cc  cc   	     
    	   
         Gg� �� (	� (�                 nYE 11         8:�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             nn  )          == �����������������������������������������������������������������������������                                ��     �  Y�   @  #   �   �                                                                                '   5  1n1YE  n)n    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��AS��Ak���  !���7��lKü\��s��p|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��kK��\��s��o|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��kK��[��s��o|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��kK��[��s��o|8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��jK��[��s��o|8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��jK��[��s��o|8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��iK��[��s��o|8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��hK��Z��s��o|8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��hK��Z��r��o|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��gK��Z��r��o|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��fK��Z��q��o|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��Ak���  s��7��fK��Z��q��n|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��Ak���  !���7��eK��Z��q��n|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��Ak���  !���7��dK��Y��p��n|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ak���  !���7�� cK��Y��p��n|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  !���7�� cK��Y��o��n|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  !���7�� bK��Y��o��n|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  !���7�� bK��Y��n��n|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  !���7�� aK��Y��ns�n|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  !���7�� aK��X��ns�n|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  !���7�� aK��X��ms�n|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  !���;��aK��X��ms�m|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  !���;��aK��X��ms�m|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��aK��X��ms�m|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��aK��W��mӀm|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��W��mӀm|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��W��lӀm|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��W��lӀm|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��W��lӀl|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��W��kӀl|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��V��kӀl|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��V��jӀk|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��V��jӀk|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��V��jӀj|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��V��jӀj|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��`K��VS�jӄi|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;��`K��US�j�i|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;��`K��US�j�h|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;��`K��US�i�h|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;��`K��US�i�g|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;��`K��US�i�f|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;��`K��US�h��f|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;��`K��US�h��e|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�T`K��TS�h��e|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�T`K��TS�h��e|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�T`K��TS�h��d|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�d;�T`K��TS�h��d|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�d;�T`K��TS�h��d|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�d;�T`K��TS�h��c|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�d;�T`K��Tc�h��b|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�d;�T`K��Tc�h��b|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�d;�T`@c�Tc�h��a|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�d;�T`@c�Tc�h��a|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�d;�T`@c�Tc�h��`|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�d;�T`@c�Tc�h��_!�8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�T_@c�Tc�h��_!�8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�T_@c�Tc�h��_!�8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�d_@c�Tc�h��_!�8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�d_@c�Sc�h��^!�8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�d_@c�Sc�h��^!�8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�d_@c�Sc�g��^!�8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�d_@c�Sc�g��^!�8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�d_@c�Sc�g��]!�8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�d_@c�Sc�g��]!�8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;�d_@c�Sc�g��]!�8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d_@c�Sc�g��]|8T0 k� �C�#t� %Q8D"!6�0d   �    � $ ���AS��Ao���  s��;�d_@c�Sc�g��]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d_@c�Sc�g��]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d_@c�Sc�g��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d_@c�Sc�gà]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d_@c�Sc�gà]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gà]|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;�d^@c�Rc�gà]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gà]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gä]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gä]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gä]!�8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gä]!�8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gä]!�8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gä]!�8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gӤ]!�8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gӤ]!�8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gӤ]!�8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^@c�Rc�gӤ]!�8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^K��Rc�gӤ]!�8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^K��Rc�gӤ]!�8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^K��Rc�g �]!�8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^K��Rc�g �]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d^K��Rc�g �]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d]K��Rc�g �]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d]K��RS�g �]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d]K��RS�g��]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d]K��RS�g��]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d]K��RS�g��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d]K��RS�g��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d]K��RS�g��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d]K��R��g��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�d]K��R��g��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T]K��R��g��]|8T0 k� �C�$� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T ]K��R��g��]|8T0 k� �C�$� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T ]K��R��g��]|8T0 k� �C�$� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T ]K��Q��f��]|8T0 k� �C�$� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T ]K��Q��f��]|8T0 k� �C�$� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T ]K��Q��f��]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� ]K��Q��e��]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� ]K��Q��e��]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� ]K��Q��e��]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��$\K��Q��e��]|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;��$\K��Q��d��]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T$\K��Q��d��]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T$\K��P��d��]|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;�T$\K��P��d��]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T$[K��P��d �]|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;�T [K��P��d �]|8T0 k� �C�#d� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��P��d �]|8T0 k� �C�#d� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��P��d �]|8T0 k� �C�#d� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��P��d �]|8T0 k� �C�#d� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��P��d��]|8T0 k� �C�#d� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��P��d��]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��P��d��]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��O��d��]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��O��d��]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T [K��O��d��]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T [K��O��d��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T [K��O��e��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T [K��O��e��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T [K��O��e��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�T [K��O��e��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��O��e��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��O��e��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��O��e��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��O��e��]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��N��e �]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��N��e �]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��N��e �]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��N��e �]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��N��e �]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��N��e �]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��N��eC�]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��N��eC�]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��N��eC�]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��N��eC�]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [K��N��eC�]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [K��N��eC�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [K��N��eC�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [K��NS�eC�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [K��NS�eC�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [@c�NS�eC�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [@c�NS�eC�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [@c�NS�eC�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [@c�NS�e�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [@c�NS�e�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [@��NS�e�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��NS�e�]|8T0 k� �C�$� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��NS�e�]|8T0 k� �C�$� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��NS�eS�]|8T0 k� �C�$� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��NS�eS�]|8T0 k� �C�$� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��NS�eS�]|8T0 k� �C�$� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��NS�eS�]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��Nc�eS�]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��Nc�eS�]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��Nc�eS�]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��Nc�eS�]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�d;�$ [@��Nc�eS�]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�d;�$ [@��Nc�eS�]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�d;�$ [@��Nc�eS�]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�d;�$ [@��Nc�eS�]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�d;�$ [@��Nc�eS�]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�d;�$ [@��Nc�eS�]|8T0 k� �C�#T� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�d;�$ [@��Nc�ec�]|8T0 k� �C�#T� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�d;�$ [@��Nc�ec�]|8T0 k� �C�#T� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�d;�$ [@��Nc�ec�]|8T0 k� �C�#T� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [@��Nc�ec�]|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s�T;�$ [@��Nc�ec�]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [K��Nc�ec�]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [K��Nc�ec�]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [K��Nc�ec�]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [K��Nc�ec�]|8T0 k� �C�#t� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s�T;�$ [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�$ [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;� [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��Nc�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��Nc�ec�]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� [K��Nc�ec�]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� ZK��Nc�ec�]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�� ZK��Nc�ec�]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��Nc�ec�]|8T0 k� �C�#İ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��Nc�ec�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��Nc�ec�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��NS�ec�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��NS�ec�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��NS�ec�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��NS�ec�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��NS�ec�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��NS�ec�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��NS�ec�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��NS�ec�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��NS�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��NS�ec�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��ZK��N��eS�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��eS�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��eS�]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��eS�]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��eS�]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��eS�]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��e�]|8T0 k� �C�#4� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��e�]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��e�]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��e�]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��e�]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��N��e�]|8T0 k� �C�#D� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�ZK��M��e�]|8T0 k� �C�#T� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�YK��M��e�]|8T0 k� �C�#T� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�YK��M��e�]|8T0 k� �C�#T� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�YK��M��e�]|8T0 k� �C�#T� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�YK��M��e�]|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;�YK��M��e�]|8T0 k� �C�#d� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�YK��M��e�]|8T0 k� �C�#d� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�TYK��M��e�]|8T0 k� �C�#d� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�TYK��M��e�]|8T0 k� �C�#d� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�TYK��L��e�]|8T0 k� �C�#d� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�TYK��L��e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�TYK��L��e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�TYK��L��e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�TYK��L��e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YK��L��e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA�L��e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA�L��e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA�L��e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA�L��e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA�LS�e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA�LS�e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YAS�LS�e�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YAS�LS�f�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YAS�LS�f�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YAS�LS�f�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YAS�LS�f�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA��LS�f�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��XA��LS�f�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��XA��LS�fS�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��XA��LS�fS�]|8T0 k� �C�#�� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA��LS�fS�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA��LS�fS�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA��LS�gS�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA��Lc�gS�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA��Lc�gS�]|8T0 k� �C�#԰ %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;��YA��Lc�gS�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�TYD��Lc�gS�]|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ao���  s��;�TYD��Mc�gS�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�TYD��Mc�gS�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ���AS��Ao���  s��;�TYD��Mc�gS�]|8T0 k� �C�#� %Q8D"!6�0d   ��    � $ ��/�AS?�A+��'�  ,S������W�Tr��T!$|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ��/�ASC�A/��#�  ,S������[�Tr��T!#,	|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ��+�ASC�A/��#�  ,S������[�Tr��X!#0|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ��+�ASG�A/��#�  ,S������[�Tr��X!#4|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ��+�ASG�A/��#�  s������[�Tr��X!#<|8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ��+�ASK�A3��#�  s������[�Tr��\"#@|8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ��+�ASK�A3��#�  s������[�Tr��\"�H|8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ��+�ASO�A3��#�  s������[�Tr��\"�L|8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ��+�ASO�A3��#�  s������[�Tr��`"�T|8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ��'�ASO�A3��#�  s������[�Tr��`"�X|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ��'�ASS�A7��#�  s������[�Tr��d"�`|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ��'�ASS�A7��#�  s������[�Tr��d"�d|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ��'�ASW�A7��#�  s�����[�Tr��d"�l|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ��'�ASW�A7��#�  s�����[�Tr��d"�p|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ��'�AS[�A7��#�  s�����_�Tr��h"�x|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ��'�AS[�A;��#�  s�����_�Tr��h"�||8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ��'�AS[�A;��#�  s�����_�Tr��l"��|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ��'�AS_�A;��#�  s�����_�Tr��l"ӈ|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ��#�AS_�A;���  s�����_�T���l"ӌ!|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ��#�ASc�A;���  s�����_�T���p"Ӕ"|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ��#�ASc�A?���  s�����_�T���t#Ә$|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ��#�ASc�A?���  s�����_�T���t#Ӝ%|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ��#�ASg�A?���  s�����_�T���x#Ӡ&|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ��#�ASg�A?���  s����D_�T���|$Ө'|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ��#�ASg�A?���  s����D_�T���|$Ӭ)|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ��#�ASk�A?���  s����Dc�T���$Ӱ*|8T0 k� �C�#D� %Q8D"!6�0d   ��  � $ ��#�ASk�AC���  s����Dc�T���%Ӵ+|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ��#�ASk�AC���  s����Dc�Ub��%Ӽ,|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���ASo�AC���  s����Dg�Ub��&��-|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���ASo�AC���  s����Dg�Ub��&��/|8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���ASo�AC���  s����Dg�Ub��'��0|8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���ASs�AC���  s����Dk�Ub��'��1|8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���ASs�AG���  s����Dk�Ub��(��2|8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���ASs�AG���  s����Dk�Ub��)��3|8T0 k� �C�#d� %Q8D"!6�0d   ��   � $ ���ASw�AG���  s����Dk�Ub��)��4|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���ASw�AG���  s����To�Ub��*��5|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���ASw�AG���  s��T�To�E���+��6!�8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS{�AG���  s��T�To�E���,��7!�8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS{�AG���  s��T�Ts�E���,��8!�8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS{�AK���  s��T�Ts�E���-��9!�8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS{�AK���  s��T�Ts�E���.��:!�8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS�AK���  s��T�Ts�E���/��;!�8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS�AK���  s��T�Tw�E���0��<!�8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS�AK���  s��T�Tw�E���1��=!�8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS�AK���  s��T�Tw�E���2� >!�8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��AK���  s��T�Tw�E���3�?!�8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��AK���  s��d�d{�F��4�@!�8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��AO���  s��d�d{�F��5�A|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��AO���  s��d�d{�F��6�A|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��AO���  s��d�d{�F��7�B|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��AO���  s��d�d�F��8�C|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��AO���  s��d�d�D�� �9�D|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��AO���  s��d�d�D�� �;�E|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��AO���  s��d�d�D��!<� F|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��AO���  s��d�d��D��!=�$F|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��AO���  s��T�d��D��">�$G|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��AS���  s��T�d��D��#?�(H|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��AS���  s��T�t��D��#@�,I|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��AS���  s��T�t��D��$ A�0I!�8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��AS���  s��T�t��D��%(B�0J!�8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ���AS��AS���  s��T�t� D��&0C�4K!�8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ���AS��AS���  s��T�t�D��'�8D�8K!�8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ���AS��AS���  s��T�t�D� '�<E�8L!�8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ���AS��AS���  s��T�ĄD�(�DF�<M!�8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ���AS��AS���  s����ĄD�)�LG�@N!�8T0 k� �C�#� %Q8D"!6�0d   ��  � $ ���AS��AS���  s����ĄD�*�TH�@N!�8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��AW���  s����Ĉ
D�+�XI�DO!�8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��AW���  s����ĄD�,�`I�HO!�8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��AW���  s����ĄD�-�hJ�HP!�8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��AW���  s���#�ĄD�.�pK�LQ|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ���AS��AW���  s���#�ĄD� /�xL�PQ|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ���AS��AW���  s���#�ĄD�$0��M�PR|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ���AS��AW���  s���#�ĄD�(1��N�TS|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ���AS��AW���  s���#���D�,2��N�TS|8T0 k� �C�$� %Q8D"!6�0d   ��   � $ ���AS��AW���  s���#���D�04��O�XT|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��AW���  s���#���D�45��P�XT|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��AW���  s���#���D�86��Q�\U|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��AW���  s���#��|D�<7��Q�`V|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���#��|D�D8	�R�`V|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���#��x!D�H:	�R�dW|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���#��x"D�L;	�S�dX|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��t$D�P<	�S�hY|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��t&D�X=	�T�hZ|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��p(D�\?	#�T�h[|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��p*Ls`@	#�U�l\|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��l,LsdA	#�U�l]|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��h.LslB	#�U�l^|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��h0LspD	#�U�p_|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��d2LstE	�U�p`|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��`3LsxF	�V�pa|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��\5Ls|G	�V�pb|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��A[���  s���'��X7Ls�H	�V�pc|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���'��X9Ls�I	�V�lc|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���'��T;Ls�K	#�V�hd|8T0 k� �C�#t� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���'��P=Ls�L	#�V�he|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+��L?Ls�M	#�V�de|8T0 k� �C�#�� %Q8D"!6�0d   ��  � $ ���AS��A_���  s���+��HALs�N	#�V�`f|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+��DCLs�O	#�V�\f|8T0 k� �C�#�� %Q8D"!6�0d   ��  � $ ���AS��A_���  s���+��@EL��P	�V�Xg|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+��@GL��Q	 V�Tg|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+��<IL��R	 V�Ph|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+�	t8JL��S	 V�Lh|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+�	t4LL��T	 V�Hi|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+�	t4ML��U	#�V�Di|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+�	t4NL��V	#�W�@j|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+�	t4OL��V	#�W�8j|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+�	�4OL��W	#�X�4k|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+�	�4PL��W	#�Y�0k|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��A_���  s���+�	�8PL��X��Z�(l|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���+�	�8QL��Y� [�$l|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���+�	�8RL��Z� \� l|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���+��8RL��[� \�l|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���+��8SL��\� ]�m|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���/��4TL��\� ]�m|8T0 k� �C�#İ %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���/��4TL��\� ^�n|8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���/��4TL��]��^�o|8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���/��4UL��]��_� o|8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���/��4UL��^��_��p|8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���/��4VL��^��_��p|8T0 k� �C�#԰ %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���/��4VL��^��`��q|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���/��4VL��_��`��q|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���/��4WL��`��a��q|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s���/�4WL��`��a��q|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s� �/�4XL��a��b��r|8T0 k� �C�#� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s� �/�4XL��b��b��r|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s� �/�4YL��b��c��r|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s� �/�4ZL��b��c��r|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s� �/�4ZL��b��c��r|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s� �/�4[L��b�d��s|8T0 k� �C�#�� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s� �/�0[L��b�d��s|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s� �/�0[L��b�e�s|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ac���  s� �/�0\L��b�e�s|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� �/�0\L��b�e�s|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� �/�0]L��c�f�s|8T0 k� �C�#4� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� �/�$0]L��c�f�t|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� �/�$0^L��c�f�t|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� �3�$0^L��c�g�t|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� �3�$0_L��c�g�t|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� �3�$0_L��c�h�s|8T0 k� �C�#D� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� �3�$0`Ls�c�h�s|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� �3�$,`Ls�c�h�s|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� �3�$,`Ls�c�iӠs|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� T3�$,aLs�c�iӠs|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� T3�$,aLs�c�iӠs|8T0 k� �C�#T� %Q8D"!6�0d   ��   � $ ���AS��Ag���  s� T3�