GST@�                                                            \     �                                               � ���  ��                    ���2����
 J���������������z���        �h     #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    "�j��,  " ��
  ��                                                                              ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������o=  0  o4   1  +      '           �                    	�  7�  V�  	�                    
          : �����������������������������������������������������������������������������                                �d      C  ��   @  #   �   �                                                                                '       )n)n1n  
    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    K��{BC�L��M,[�w|( �_�A�LE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K� {BC�L��M,[��w|( �_�A�HE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K� {BC�@�M,[��w|( �_�A�HE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K� {BC�@�M0[��w|( �_�A�HE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�{BC�@�M0[��x|( �_�A�HE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�zBC�@�M0[��x|( �_�A�HE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�zBC�@�M0[��x|( �_�A�HE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�zBC�BA�M0[��x|( �_�A�HE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�z2C�BA�M4[��w|( �_�A�HE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�z2C�BA�M4[��w|( �_�A�HE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�z2C�BA�M4\��w|( �_�A�HE_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��   �  }K�y2C�BA�N4\Q�w|( �_�A�HE_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�y2C�D��N8\Q�w|( �_�A�HE_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�y2C�D��N8\Q�v|( �_�A�HE_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�y�C�D��N�8\Q�v|( �_�A�HE_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�y�C�D��O�8\Q�v|( �_�A�HE_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�y�C�D��O�8\Q�v|( �_�A�HE_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�y�C�D��O�<\Q�u|( �_�A�HE_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�x�C�D��O�<\Q�u|( �_�A�HF_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�x�C�D��O�<\Q�u|( �_�A�HF_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�x�C�D��O�<\Q�u|( �_�A�HF_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�x�C�D��OR<\Q�u|( �_�A�HF_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�x�C�D��OR<\Q�t|( �_�A�HF_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�x�C�D��OR<]Q�t|( �_�A�HF_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K�x�C�D��OR<]Q�t|( �_�A�DF_�B�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }A^�S���F�F l3� ���8$��pA�S��P0_xT3�T0 k� ��W��W%�0d  U89D"!   ��"    � �FA^�S���F�G l3� ���8$��qA�S��P,_tT3�T0 k� ��X��X%�0d  U89D"!   ��"    � �FA^�S���F�I l7� ���8$��rA�W��P(_pU3�T0 k� ��X��X%�0d  U89D"!   ��"    � �FA^�S���F|K l;� ���<$��sA�W���P$_lU3�T0 k� ��Y��Y%�0d  U89D"!   ��"    � �FA^�S���F|L l;� ���<$��tA�W���P _hV3�T0 k� ��Z��Z%�0d  U89D"!   ��"    � �FA^�S���F|N l?� ���<$� uA�[���P_dV3�T0 k� ��[��[%�0d  U89D"!   ��"    � �FA^�S���FxP l?� ���<$�vA�[���P_`W3�T0 k� ��]��]%�0d  U89D"!   ��"    � �FA^�S���FxQ lC� ��<$|vA�_���P _\W3�T0 k� ��_��_%�0d  U89D"!   ��"    � �FA^�S���FxS lC� ��<$|wA�_���P _XW3�T0 k� ��`��`%�0d  U89D"!   ��"    � �FA^�S���FxU lG� ��<$|wA�c���P!_TX3�T0 k� ��b��b%�0d  U89D"!   ��"    �  �FA^�S���FxV lG� ��<$|xA�c���P!_PX3�T0 k� ��d��d%�0d  U89D"!   ��"    � !�FA^�S���FxX lK� ��<$| xA�g���P"_LY3�T0 k� ��f��f%�0d  U89D"!   ��"    � "�FA^�S���FxZ lO� ��<$|$yA�g���P"_HY3�T0 k� ��g��g%�0d  U89D"!   ��"    � #�FA^�S���H�x\ lO� ��<$|(yA�g���P#_HY3�T0 k� ��j��j%�0d  U89D"!   ��"    � $�FA^�S���H�x] lS� ��@$|,yA�k���P #_DZ3�T0 k� ��l��l%�0d  U89D"!   ��"    � %�FA^�S���H�x_ lS� ��@$|0zA�k���_�$_@Z3�T0 k� ��n��n%�0d  U89D"!   ��"    � &�FA^�S���H�xa lW� ��@$|4zA�o���_�$_<[3�T0 k� ��p��p%�0d  U89D"!   ��" 
   � '�FA^�S���H�xb lW� ��@$l8zA�o���_�%_8[3�T0 k� ��r��r%�0d  U89D"!   ��" 
   � (�FA^�S���H�xd lW� ��@$l<zA�l ��_�%_4[3�T0 k� ��t��t%�0d  U89D"!   ��" 
   � )�FA^�S���H�xe l[� ��@#l@zA�p��_�&_4\3�T0 k� ��u��u%�0d  U89D"!   ��" 
   � *�FA^�S���H�xg l[� ��@#lDzA�p��_�&_0\3�T0 k� ��w��w%�0d  U89D"!   ��" 
   � +�FA^�S���H�xh l_� ��@#lDyA�p��_�'_,\3�T0 k� ��x��x%�0d  U89D"!   ��" 
   � ,�FA^�S���H�xj l_� ��@#,@wA�t��_�'_(]3�T0 k� ��z��z%�0d  U89D"!   ��" 
   � -�FA^�S���H�xk lc� ��@#,@vA�t��_�(_(]3�T0 k� ��x��x%�0d  U89D"!  �" 
   � .�MA^�S���H�xm lc� ��@#,@uA�t��_�(_$^3�T0 k� ��w��w%�0d  U89D"!  ��/ 
   � /�TA^�S���H�xm lg� ��@#,<tA�x��_�(_ ^3�T0 k� ��u��u%�0d  U89D"!  ��/ 
   � 0�[A^�S���H�xn lg� ��D#,8sA�x��_�)_^3�T0 k� ��t��t%�0d  U89D"!  ��/ 
   � 1�bA^�S���H�|o lg� ��D#�8rA�x��_�)__3�T0 k� ��r��r%�0d  U89D"!  ��/ 
   � 2�iA^�S���H�|p lk� ��D#�4rA�|��_�*__3�T0 k� ��q��q%�0d  U89D"! 	 ��/ 
   � 3�oA^�S���I|q lk� ��D#�0qA�|��_�*__3�T0 k� ��o��o%�0d  U89D"! 
 ��/ 
   � 4�uA^�S���I�s lo� ��D#�0pA�|	��_�+__3�T0 k� �n�n%�0d  U89D"!  ��/ 
   � 5�{A^�S���I�t lo� ��D#�,oA��	��_�+_`3�T0 k� �m�m%�0d  U89D"!  ��/ 
   � 6��A^�S���I�u lo� ��D#�,nA��
��_�+_`3�T0 k� �$k�(k%�0d  U89D"!  ��/ 
   � 7��A^�S���I�t ls� ��D#�(mA��
��_�,_`3�T0 k� �4j�8j%�0d  U89D"!  ��/ 
   � 8��A^�S���I�t ls� ��D#�$mA����_�,_a3�T0 k� �Dh�Hh%�0d  U89D"!  ��/ 
   � 9��A^�S���I�t lw� ��D#�$lA����_�,_a3�T0 k� �Tg�Xg%�0d  U89D"!  ��/ 
   � :��A^�S���I�t lw� ��D#� kA����_�-_a3�T0 k� �de�he%�0d  U89D"!  ��/ 
   � ;��A^�S���I�s lw� ��D#� jA����_�-_ b3�T0 k� �td�xd%�0d  U89D"!  ��/ 	   � <��A^�S���I�s l{� ��D#�iA����_�-_ b3�T0 k� ��b��b%�0d  U89D"!  ��/ 	   � <��A^�S���I�s l{� #��D#�iA����_�.^�b3�T0 k� ��a��a%�0d  U89D"!  ��/ 	   � <��A^�S���I�s l{� #��D#�hA����_�.^�b3�T0 k� ��_��_%�0d  U89D"!  ��/ 	   � <��A^�S���I�r l� #��H#�gA����_�/^�c3�T0 k� ��^��^%�0d  U89D"!  ��/ 	   � <��A^�S���I�r l� #��H#�gA����_�/^�c3�T0 k� ��]��]%�0d  U89D"!  ��/ 	   � <��A^�S���I�r l� #��H#�fA����_�/^�c3�T0 k� ��[��[%�0d  U89D"!  ��/ 	   � <��A^�S���I�r l�� '��H#�eA���_�0^�c3�T0 k� ��Z��Z%�0d  U89D"!  ��/ 	   � <��A^�S���I�r l�� '��H#�eA���_�0^�d3�T0 k� ��X��X%�0d  U89D"!  ��/ 	   � <��A^�S���I�q l�� '��H#�dA��{�_�0^�d3�T0 k� �W�W%�0d  U89D"!  ��/ 	   � <��A^�S���I�q l�� '��H#�cA��{�_�0^�d3�T0 k� �U�U%�0d  U89D"!  ��/ 	   � <��A^�S���I�q l�� '��H#�cA��w�_�1^�d3�T0 k� �$T�(T%�0d  U89D"!   ��/ 	   � <��A^�S���I�q l�� '��H#�bA��w�_�1^�e3�T0 k� �4R�8R%�0d  U89D"! ! ��/ 	   � <��A^�S���BL�q l�� +��H#�aA��s�_�1^�e3�T0 k� �DQ�HQ%�0d  U89D"! ! ��/ 	   � <��A^�S���BL�p l�� +��H#�aA��s�_�2^�e3�T0 k� �TO�XO%�0d  U89D"! " ��/ 	   � <��A^�S���BL�p l�� +��H#� `A��o�_�2^�e3�T0 k� �dN�hN%�0d  U89D"! # ��/ 	   � <��A^�S���BL�p l�� +��H#� _A��o�_�2^�e3�T0 k� �tL�xL%�0d  U89D"! $ ��/ 	   � <��A^�S���BL�p l�� +��H#� _A��k�_�2^�f3�T0 k� ��K��K%�0d  U89D"! % ��/    � <��A^�S���BL�p l�� +��H#��^A��k�_�3^�f3�T0 k� ��J��J%�0d  U89D"! % ��/    � <��A^�S���BL�p l�� +��H#��]A��g�_�3^�f3�T0 k� ��H��H%�0d  U89D"! & ��/    � <��A^�S���BL�o l�� /��H#��\A��g�_�3^�f3�T0 k� ��G��G%�0d  U89D"! ' ��/    � < A^�S���BL�o l�� /��H#��\A��g�_�4^�g3�T0 k� ��E��E%�0d  U89D"! ' ��/    � < A^�S���BL�o l�� /��L#��[A��c�_�4^�g3�T0 k� ��D��D%�0d  U89D"! ( ��/    � < 	A^�S���BL�o l�� /��L#��ZA��c�_�4^�g3�T0 k� ��B��B%�0d  U89D"! ( ��/    � < A^�S���BL�o l�� /��L#��ZA��_�_�4^�g3�T0 k� ��A��A%�0d  U89D"! ) ��/    � < A^�S���BL�o l�� /��L#��YA��_�_�5^�g3�T0 k� � ?�?%�0d  U89D"! * ��/    � < A^�S���BL�n l�� /��L#��XA��[�_�5^�g3�T0 k� �>�>%�0d  U89D"! * ��/    � < A^�S���BL�n l�� 3��L#��XA��[�_�5^�h3�T0 k� � <�$<%�0d  U89D"! + ��/    � < A^�S���BL�n l�� 3��L#��WA��[�_�5^�h3�T0 k� �0;�4;%�0d  U89D"! + ��/    � < !A^�S���BL�n l�� 3�!�L#��VA��W�_�5^�h3�T0 k� �@9�D9%�0d  U89D"! + ��/    � < %A^�S���BL�n l�� 3�!�L#��VA��W�_�6^�h3�T0 k� �P8�T8%�0d  U89D"! , ��/    � < )A^�S���BL�n l�� 3�!�L#��UA��W�_�6^�h3�T0 k� �`7�d7%�0d  U89D"! , ��/    � < -A^�S���BL�n l�� 3�!�L#��TA��S�_�6^�i3�T0 k� �p5�t5%�0d  U89D"! - ��/    � < 1A^�S���BL�m l�� 3�!�L#��TA��S�_�6^�i3�T0 k� ��4��4%�0d  U89D"! - ��/    � < 5A^�S���BL�m l�� 3�!�L#��SA��O�_�7^�i3�T0 k� ��2��2%�0d  U89D"! - ��/    � < 9A^�S���BL�m l�� 7�!�L#��SA��O�_�7^�i3�T0 k� ��1��1%�0d  U89D"! - ��/    � < =A^�S���BL�m l�� 7�!�L"��RA��O�_�7^�i3�T0 k� ��/��/%�0d  U89D"! . ��/    � < AA^�S���BL�m l�� 7�!�L"��RA��K�_�7^�i3�T0 k� ��.��.%�0d  U89D"! . ��/    � < EA^�S���BL�m l�� 7�!�L"��QA��K�_�7^�j3�T0 k� ��,��,%�0d  U89D"! . ��/    � < IA^�S���BL�m l�� 7�!�L"��PA��K�_�8^�j3�T0 k� ��+��+%�0d  U89D"! . ��/    � < MA^�S���BL�m l�� 7��L"��PA��G�_�8^�j3�T0 k� ��)��)%�0d  U89D"! . ��/    � < QA^�S���BL�l l�� 7��L"��OA��G�_�8^�j3�T0 k� � (�(%�0d  U89D"! / ��/    � < UA^�S���BL�l l�� 7��L"��OA��G�_�8^�j3�T0 k� �'�'%�0d  U89D"! / ��/    � < YA^�S���BL�l l�� 7��L"��NA��C�_�8^�j3�T0 k� � %�$%%�0d  U89D"! / ��/    � < ]A^�S���BL�l l�� ;��L"��NA�� C�_�9^�j3�T0 k� �0$�4$%�0d  U89D"! / ��/    � < aA^�S���BL�l l�� ;��L"��MA�� C�_�9^�k3�T0 k� �@"�D"%�0d  U89D"! / ��/    � < eA^�S���BL�l l�� ;��P"��MA�� C�_�9^�k3�T0 k� �P!�T!%�0d  U89D"! / ��/    � < iA^�S���BL�l l�� ;��P"��LA��!< _�9^�k3�T0 k� �`�d%�0d  U89D"! / ��/    � < mA^�S���BL�l l�� ;��P"��LA��!< _�9^�k3�T0 k� �p�t%�0d  U89D"! / ��/    � < qA^�S���BL�l l�� ;��P"��KA��!< _�9^�k3�T0 k� ����%�0d  U89D"! . ��/    � < uA^�S���BL�k l�� ;��P"��KA��!8 _�:^�k3�T0 k� ���%�0d  U89D"! . ��/    � < yA^�S���BL�k l�� ;�!�P"��KA��"8 _�:^�k3�T0 k� ���%�0d  U89D"! . ��/    � < }A^�S���BL�k l�� ;�!�P"��JA��"8 _�:^�l3�T0 k� ���%�0d  U89D"! . ��/    � < �A^�S���BL�k l�� ;�!�P"��JA��"8 _�:^�l3�T0 k� ���%�0d  U89D"! . ��/    � < �A^�S���BL�k l�� ?�!�P"��IA��"4 _�:^�l3�T0 k� ����%�0d  U89D"! . ��/    � < �A^�S���BL�k l�� ?�!�P"��IA��#4_|:^�l3�T0 k� ����%�0d  U89D"! - ��/    � < �A^�S���BL�k l�� ?�!�P"��HA��#4_|;^�l3�T0 k� ����%�0d  U89D"! - ��/    � ; �A^�S���BL�k l�� ?�!�P"��HA��#4_|;^�l3�T0 k� ��� %�0d  U89D"! - ��/    � : �A^�S���BL�k l�� ?�!�P"��HA��#0_|;^�l3�T0 k� ��%�0d  U89D"! , ��/    � 9 �A^�S���BL�k l�� ?�!�P"��GA��$0_|;^�l3�T0 k� �� %�0d  U89D"! , ��/    � 8 �A^�S���BL�k l�� ?�!�P"��GA��$0_x;^�l3�T0 k� �,�0%�0d  U89D"! , ��/    � 7 �A^�S���BL�j l�� ?�!�P"��FA��$0_x;^�m3�T0 k� �<�@%�0d  U89D"! + ��/    � 6 �A^�S���BL�j l�� ?��P"��FA��$0_x;^�m3�T0 k� �L	�P	%�0d  U89D"! + ��/    � 5 �A^�S���BL�j l�� ?��P"��FA��%,_x<^�m3�T0 k� �\�`%�0d  U89D"! * ��/    � 4 �A^�S���BL�j l�� ?��P"��EA��%,_x<^�m3�T0 k� �l�p%�0d  U89D"! * ��/    � 3 �A^�S���BL�j l�� ?��P"��EA��%,_t<^�m3�T0 k� �|��%�0d  U89D"! ) ��/    � 2 �A^�S���BL�j l�� C��P"��EA��%,_t<^�m3�T0 k� ���%�0d  U89D"! ) ��/    � 1 �A^�S���BL�j l�� C��P"��DA��%(_t<^�m3�T0 k� ���%�0d  U89D"! ( ��/    � 0 �A^�S���BL�j l�� C��P"��DA��&(_t<^�m3�T0 k� ���%�0d  U89D"! ( ��/    � / �A^�S���BL�j l�� C��P"��DA��&(_t<^�m3�T0 k� �����%�0d  U89D"! ' ��/    � . �A^�S���BL�j l�� C��P"��CA��&(_t<^�n3�T0 k� ������%�0d  U89D"! & ��/    � - �A^�S���BL�j l�� C��P"��CA��&(_p=^�n3�T0 k� ������%�0d  U89D"! & ��/    � , �A^�S���BL�j l�� C��P"��CA��&$_p=^�n3�T0 k� ������%�0d  U89D"! % ��/    � + �A^�S���BL�j l�� C��P"��BA��'$_p=^�n3�T0 k� �����%�0d  U89D"! $ ��/    � * �A^�S���BL�i l�� C��P"��BA��'$_p=^�n3�T0 k� ����%�0d  U89D"! # ��/    � ) �A^�S���BL�i l�� C��P"��BA��'$_p=^�n3�T0 k� ���#�%�0d  U89D"! # ��/    � ( �A^�S���BL�i l�� C��P"��AA��'$_p=^�n3�T0 k� �/��3�%�0d  U89D"! " ��/    � ' �A^�S���BL�i l�� C��P"��AA��'$_p=^�n3�T0 k� �?��C�%�0d  U89D"! ! ��/    � & �A^�S���BL�i l�� C��P"��AA��( _l=^�n3�T0 k� �O��S�%�0d  U89D"!   ��/    � % �A^�S���BL�i l�� C��P"��AA��( _l=^�n3�T0 k� �_��c�%�0d  U89D"!  ��/    � $ �A^�S���BL�i l�� C��T"��@A��( _l>^�n3�T0 k� �o��s�%�0d  U89D"!  ��/    � # �A^�S���BL�i l�� G��T"��@A��( _l>^�o3�T0 k� �����%�0d  U89D"!  ��/    � " �A^�S���BL�i l�� G��T"��@A��( _l>^�o3�T0 k� �����%�0d  U89D"!  ��/    � ! �A^�S���BL�i l�� G��T"��?A��( _l>^�o3�T0 k� �����%�0d  U89D"!  ��/    �   �A^�S���BL�i l�� G��T"��?A��)_l>^�o3�T0 k� �����%�0d  U89D"!  ��/    �  �A^�S���BL�i l�� G��T"��?A��)_h>^�o3�T0 k� �����%�0d  U89D"!  ��/    �  �@�x �P"�F pX b|  �`@�`xStF ��T X� T0 k� �8F�<F%�0d  U89D"!  ��/    �  @�x �P"�F pX b|  �`@�`xStF ��T X� T0 k� �8F�<F%�0d  U89D"!   /�/    �  �@�x �P"�F pX b|  �`@�`xStF ��T X� T0 k� � J�$J%�0d  U89D"!   ��/    �  �@�x �@�F pX b|  �`@�`x�tF ��T X� T0 k� �L�L%�0d  U89D"!   ��/    �   �@�x �@�F pX b|  �`@�`x�pF ��T X�T0 k� �M�M%�0d  U89D"!   ��/    � ! �@�x �@�F pX b|  �`@�`x�pF ��T X�T0 k� �N�N%�0d  U89D"!   ��/    � " �@�x �@�F tX b|  �`@�`x�pF ��T X�T0 k� �O�O%�0d  U89D"!   ��/    � # �@�x �@�F tX b|   �`@�`x�hF ��T X�T0 k� ��P� P%�0d  U89D"!   ��/    � $ �CCxSBB�F�tX|  S`C�`x�`F ��T X�T0 k� ��Q��Q%�0d  U89D"!   ��/    � % �CCwSBB�F�tX|$ S`C�\w�XF�� X�T0 k� ��S��S%�0d  U89D"!   ��/    � & �CCwSBB�F�xX|$ S`C�\w�PF�� X�T0 k� ��T��T%�0d  U89D"!   ��/    � ' �CCvSBB�F�xX|$ S`C�\w�HF�� X�T0 k� ��U��U%�0d  U89D"!   ��/    � ( �CCvSBB�F�|X|( S`C�\w�@F���X�T0 k� ��V��V%�0d  U89D"!   ��/    � ) �CCu�BB�F�|XR|( �`C�Xv�@F���X�T0 k� ��W��W%�0d  U89D"!   ��/    � * �CCu�BB�F��XR|( �`C�XvS@FS�3�W�T0 k� ��X��X%�0d  U89D"!   ��3    � + �CCt�BB�F��XR|( �`E3TuS<FS�3�W�T0 k� �X��X%�0d  U89D"!   ��3    � , �E#t�F�F��XR|( �`E3TuS8FS�3�W�	T0 k� �X��X%�0d  U89D"!   ��3    � - �E#s�F�F��XR|( �`E3TtS4FS�3�W�
T0 k� �X��X%�0d  U89D"!   ��3    � . �E#r�F�F��X�|( �`E3TtS0FS�3�V�T0 k� �R��R%�0d  U89D"!   ��3    � / �E#q�F�F��X�|( �`E3TsS,F��3�V�T0 k� �N��N%�0d  U89D"!   ��3    � 0 �E#p�E��F��X�|( �`E3TsS,F��3�U�T0 k� �K��K%�0d  U89D"!   ��3    � 0 �E#o�E��F��W�|( �`E3TrS(F��C�U�T0 k� �G��G%�0d  U89D"!   ��3    � 0 �Eo�E��F��W�|( �`E3TqS(F��C�T�T0 k� �E��E%�0d  U89D"!   ��3    � 0 �En�E��F��W2|( �`E3TpS(F��C�T�T0 k� �D��D%�0d  U89D"!   ��3    � 0 �El�@b�FR�V2|( �`CCTnS$F3�C�S�T0 k� ��D��D%�0d  U89D"!   ��3    � 0 �El�@b�FR�V2|( �`CCTmS F3�C�R�T0 k� ��@��@%�0d  U89D"!   �3    � 0 �Ek�@b�FR�U2|( �`CCTlS F3�c�Q�T0 k� ��<��<%�0d  U89D"!   ��?    � 0 �Ej�@b�FR�U� |( c`CCTkS F3�c�Q�T0 k� ��9��9%�0d  U89D"!   ��?    � 0 �Ei�E�E�T��|( c\E�TkSF3�c�O�T0 k� ��1��1%�0d  U89D"!   ��?    � 0 �E�h�E�E�T��|( c\E�TjSF3�c�O�T0 k� ��.��.%�0d  U89D"!   ��?    � 0 �E�h�E�E�T��|( cXE�TiSFC�S�N�T0 k� ��*��*%�0d  U89D"!   ��?    � 0 �E�h�E�E�T��|( cXE�XgSFC�S�N�T0 k� ��&��&%�0d  U89D"!   ��?    � 0 �E�g�E�D��T��|( cXE�XfSFC�S�M�T0 k� ��#��#%�0d  U89D"!   ��?    � 0 �E�f�E�D��T��|( cTE�XdSFC�S�L�T0 k� ����%�0d  U89D"!   ��?    � 0 �D�e�B��C��T��|( SPE�XbS FC���K�T0 k� ����%�0d  U89D"!   ��?    � 0 �D�e�B��C��T��|( SPE�XaS FC��K3�T0 k� ����%�0d  U89D"!   ��?    � 0 �D�e�
B��C��T��
|( SPE�X`S FC��J3�T0 k� ����%�0d  U89D"!   ��?    � 0 �D�e�	B��B��T��	|( SLC�X]S FS��I3�
T0 k� � 	�	%�0d  U89D"!   ��?    � 0 �E�d�	E��A��T��|( �L
C�X[S ES�	��I3�	T0 k� ��%�0d  U89D"!   ��    � / �E�d�E��A��T�|( �H	C�XZS ES�	��I3�T0 k� ��%�0d  U89D"!   ��    � . �E�c�E��A��T�|( �H	C�TWS FS�
	��H3�T0 k� ����%�0d  U89D"!   ��    � . �E� c�E��@��S�|( �HC�TUS FS�
	��H3�T0 k� ����%�0d  U89D"!   ��    � . �E� b�E��?��S�|( �DC�TTS FS�
	��G3�T0 k� ����%�0d  U89D"!   ��    � . �E�$b� E��>��S�|( �@C�PQ� FS�	��G3�T0 k� ����%�0d  U89D"!   ��    � . �E�(a��E��=��S��|( �<C�PQ� ES|	��G3� T0 k� ����%�0d  U89D"!   ��    � - �E�(a�� E��=��S��|( �<C�PP�ES|	��G3��T0 k� ����%�0d  U89D"!   ��    � , �E�,`r��E��;��S��|( �8C�PM�ES|	��G3��T0 k� ����%�0d  U89D"!   ��    � + �E�,`r��E��:��S��|( �4E�PM�ESx	��F3��T0 k� ����%�0d  U89D"!   ��    � * �E�0`r��E��9��S���|( �0E�PM�ESx	��F3��T0 k� ����%�0d  U89D"!   ��    � * �E�0`r��E��8��S���|( �0E�PL�DSt	��F3��T0 k� ����%�0d  U89D"!   ��    � ) �E�0_r��E��5��S���|( �+�E�PL�DSl	��F3��T0 k� ����%�0d  U89D"!   ��    � ( �E�0_r��E��4��S���|( �+�E�PK�CSh	��F3��T0 k� ����%�0d  U89D"!   ��    � ' �E�0_r��E��3��S���|( �'�E�LK�CCd	��F3��T0 k� ����%�0d  U89D"!   ��    � & �E�4_r��E��1��S���|( �#�E�HI� BC\	��F3��T0 k� �����%�0d  U89D"!   ��    � % �E�4_r��E��/��S���|( ��E�DH��ACX��F3��T0 k� ������%�0d  U89D"!   ��    � $ �E�4_r��E��.��S���|( ��E�DF��ACX��F3��T0 k� ������%�0d  U89D"!   ��    � # �E�4_r��E��+r�S���|( ��E�<D��@CP��F3��T0 k� ������%�0d  U89D"!   ��    � " �E�4_r��E��*s R	��|( ��E�8C��?CL��F3��T0 k� ������%�0d  U89D"!   ��    � ! �E�4_r��E��)s R	��|( ��E�4B��?CH��F3��T0 k� ������%�0d  U89D"!   ��    � ! �@c4_r��E��'sR	��|( ��E�4A��>CD�F3��T0 k� ������%�0d  U89D"!   ��    �   �@c4_r��E��%%�Q	��|( ��E�,@��=3<�F3��T0 k� ������%�0d  U89D"!   ��    �  �@c4_r��E��#%�P	��|( ��E�$?�=38�F3��T0 k� ������%�0d  U89D"!   ��    �  �@c4_r��E��"%�P	!��|( ��E� >�<34�F3��T0 k� ������%�0d  U89D"!   ��    �  �@c4_r��C��%�O	!��|( ���C�<�<3,��E3��T0 k� ������%�0d  U89D"!   ��    �  �@c4_���C��%�O	!��|( ���C�;�;3(��E3��T0 k� ������%�0d  U89D"!   ��    �  �@c4_���C��%�O	!��|( ���C�:�;3$��D3��T0 k� ������%�0d  U89D"!   ��    �  �@�4_���C��%�N	��|( ���C�8�:3��C3��T0 k� ������%�0d  U89D"!   ��    �  �@�4_���C��%�N	��|( ���E��7�:3��C3��T0 k� ������%�0d  U89D"!   ��    �  �@�4_	���C��%�M	��|( ���E��7�9#��B3��T0 k� ������%�0d  U89D"!   ��    �  �@�4_	���C��%�M	��|( ���E��6�9#��B3��T0 k� ������%�0d  U89D"!   ��    �  �@�4_	���C�%� L	!��|( ���E��4�8#��@3��T0 k� ������%�0d  U89D"!   ��    �  �@�4_	���C�%� L	!��|( ���E��3�8#��?3��T0 k� ������%�0d  U89D"!   ��    �  �A4_b��C�%�$L	!��|( ���E��3|7���?3��T0 k� ������%�0d  U89D"!   ��    �  �A4_bϿC�%�$K	!��|( ���E��2t7���>3��T0 k� ������%�0d  U89D"!   ��    �  �A4_bϻC�%�(K	��|( ���E��0d6� 
��<3��T0 k� �����%�0d  U89D"!   ��    �  �A4_b˹C�%�(J	��|( ���EҼ0\6� ��;3��T0 k� �����%�0d  U89D"!   ��    �  �A4_b˷C�%�,J	��|( ���E�/T5"���:3��T0 k� �����%�0d  U89D"!   ��    �  �AS4_bǵC�%�,J	��|( ���E�.L5"���93��T0 k� �����%�0d  U89D"!   ��    �  �AS4_bǴC�%�,I	��|( ���E�.D5"���73��T0 k� �����%�0d  U89D"!   ��    �  �AS0_bðD�	%�0I	!��|( ���E�-�44"���53��T0 k� �����%�0d  U89D"!   ��    �  �AS0_b��D|%�4I	!��|( ���E�,�,4���43��T0 k� �����%�0d  U89D"!   ��    �  �C�0_b��Dt%�4H	!��|( ���E�,�(3���33��T0 k� �����%�0d  U89D"!   ��    �  �C�0_b��Dp%�4H	!��|( ���E�|+� 3���13��T0 k� �����%�0d  U89D"!   ��    �  �C�,_b��Dh%�8H	!��|( ���E�t+�3���03��T0 k� �����%�0d  U89D"!   ��    �  �C�,_b��D`s8H a��|( ���D2l+�3���/3��T0 k� �����%�0d  U89D"!   ��    �  �C�(_b��D\s8G a��|( ���D2d+�2���-3��T0 k� �����%�0d  U89D"!   ��    �  �C�(_���DTs<G a��|( ���D2\*� 2���,3��T0 k� �����%�0d  U89D"!   ��    �  �C�$_���DLs<F a��|( ���D2T*��2����*3��T0 k� �����%�0d  U89D"!   ��    �  �C�$_���DHs<F a��|( ���D2L*��1����)3��T0 k� �����%�0d  U89D"!   ��    �  �C� _���D@ c<E ���|( ���D2D*��1����'3��T0 k� �����%�0d  U89D"!   ��    �  �C�_���D;�c@E ���|( ���D2<*��1����&3��T0 k� �����%�0d  U89D"!   ��    �  �C�_���D3�c@D ���|( ���D24*��1����$3��T0 k� �����%�0d  U89D"!   ��    �  �C�_���D/�c@D ���|( ���D2(*��0� ��"3��T0 k� �����%�0d  U89D"!   ��    �  �C�_���D'�c@C ���|( ���D2 +��0s ��!3��T0 k� �����%�0d  U89D"!   ��    �  �C�_���D��@B��|( ���D2+�0s��3��T0 k� �����%�0d  U89D"!   ��    � 
 �C�_���D��<A��|( ���DB+	��0s	ӌ3��T0 k� �����%�0d  U89D"!   ��    � 
 �C�_���D��<A��|( ���DB +	��0s	ӌ3��T0 k� �����%�0d  U89D"!   ��    � 
 �C� _���D���<@��|( ���DA�,	��0s	ӌ3��T0 k� �����%�0d  U89D"!   ��    � 	 �C��_���D���<@��|( ���DA�,	��0s	ӌ3��T0 k� �����%�0d  U89D"!   ��    � 	 �D�_���C����8?���|( ���DA�-	��0s	ӌ3��T0 k� �����%�0d  U89D"!   ��    � 	 D�_���C����8?���|( ���E��-	��0s	ӌ3��T0 k� �����%�0d  U89D"!   ��    �  ~D�_���C����4>���|( ���E��-	��0s	�3��T0 k� �����%�0d  U89D"!   ��    �  }D�_���C����0=���|( ���E��-	��0�	�3��T0 k� �����%�0d  U89D"!   �    �  }D�_���E���S0=��|( ���E��.	�|0�	�3��T0 k� �����%�0d  U89D"!   �    �  }D�_���Eѿ�S,<��|( ���E��.	�t0�	�3��T0 k� �����%�0d  U89D"!   ��    �  }D�_���Eѷ�S(<��|( ���E��.	�l0��3��T0 k� �����%�0d  U89D"!   ��    �  }D�_���Eѯ�S$;��|( ���E��/	�h0��3��T0 k� �����%�0d  U89D"!   ��    �  }D�_���Eѧ�S$;��|( ���E�/	�`0��3��T0 k� �����%�0d  U89D"!   ��    �  }L�_���Eџ�S :���|( ���A��/	�\0��
3��T0 k� �����%�0d  U89D"!   ��    �  }L�_���Eї�C:���|( ���A��0	�T0��	3��T0 k� �����%�0d  U89D"!   ��    �  }L�_���Eя�C:���|( ���A��0	�P0��3��T0 k� �����%�0d  U89D"!   ��   �  }L�_���Eч�C9���|( ���A��0	�H0��3��T0 k� �����%�0d  U89D"!   ��    �  }L�_���E��C9���|( ���A��1	�D0��3��T0 k� �����%�0d  U89D"!   ��    �  }L�_���E�w�C9���|( ���A��1	�<0��3��T0 k� �{���%�0d  U89D"!   ��    �  }L�_���E�k��9���|( ���A��1Q80��3��T0 k� �{���%�0d  U89D"!   ��    �  }L�_���E�c��9���|( ���A��2Q00��3��T0 k� �{���%�0d  U89D"!   ��    �  }L�_���E�[�� 8���|( ���A��2Q,0� �3��T0 k� �{���%�0d  U89D"!   ��    �  }L�_���E�S���8���|( ���A��2Q(0� �3��T0 k� �w��{�%�0d  U89D"!   ��    �  }L�_���E�K���8��|( ���A��3Q 0� � 3��T0 k� �w��{�%�0d  U89D"!   ��    �  }L�_���E�C���8��|( ���A�x3Q0� ��3��T0 k� �w��{�%�0d  U89D"!   ��    �  }L�_��E�;���9��|( ���A�t3Q0�$��3��T0 k� �w��{�%�0d  U89D"!   ��    �  }L|_��E�3���9��|( ���A�p3Q0�$��3��T0 k� �s��w�%�0d  U89D"!   ��    �  }L"x_��E�+���9��|( ���A�l4Q0�$��3��T0 k� �s��w�%�0d  U89D"!   ��    �  }L"t_�{�E����9��|( ���A�h4Q0�$��3��T0 k� �s��w�%�0d  U89D"!   ��    �  }L"p_�{�E����9��|( ���A�`4Q0�(��3��T0 k� �s��w�%�0d  U89D"!   ��    �  }L"l_�{�E����9��|( ���A�\4Q 0�(��3��T0 k� �o��s�%�0d  U89D"!   ��    �  }L"h_�{�E����:��|( ���A�X5P�0�(��3��T0 k� �o��s�%�0d  U89D"!   ��    �  }L"d_�w�E�����:��|( ���A�T5P�0�(��3��T0 k� �o��s�%�0d  U89D"!   ��   �  }L"`_�w�E�����:��|( ���A�P5P�0�(��3��T0 k� �o��s�%�0d  U89D"!   ��    �  }L"\_�w�E�����:��|( ���A�L5P�0�,��3��T0 k� �k��o�%�0d  U89D"!   ��    �  }L"X_�w�E����:��|( ���A�H6P�0�,��3��T0 k� �k��o�%�0d  U89D"!   ��    �  }L"P_�w�E����:��|( ���A�D6P�0�,��3��T0 k� �k��o�%�0d  U89D"!   ��    �  }L"L_�s�E����;��|( ���A�@6P�0�,��3��T0 k� �k��o�%�0d  U89D"!   ��    �  }L"L_�s�E����;��|( ���A�86P�0�,��3��T0 k� �k��o�%�0d  U89D"!   ��    �  }L"H_�s�F ���;��|( ���A�47P�0�0��3��T0 k� �g��k�%�0d  U89D"!   ��    �  }L"D_�s�F ���;��|( ���A�07P�0�0��3��T0 k� �g��k�%�0d  U89D"!   ��    �  }L"@_�o�F ���;��|( ���A�,7P�0�0��3��T0 k� �g��k�%�0d  U89D"!   ��    �  }L"<_�o�F ���;��|( ���A�,7P�0�0��3��T0 k� �g��k�%�0d  U89D"!   ��    �  }L"8_�o�F ���<��|( ���A�(8P�1�0��3��T0 k� �g��k�%�0d  U89D"!   ��    �  }L"4_�o�F ���<��|( ���A�$8P�1�4��3��T0 k� �c��g�%�0d  U89D"!   ��    �  }L"0_�o�F ���<��|( ���A� 8P�1�4��3��T0 k� �c��g�%�0d  U89D"!   ��    �  }L",_�k�F ���<��|( ���A�8P�1�4��3��T0 k� �c��g�%�0d  U89D"!   ��    �  }L"(_�k�F ���<��|( ���A�8P�1�4��3��T0 k� �c��g�%�0d  U89D"!   ��    �  }L"(_�k�DЗ��<��|( ���A�9P�1�4��3��T0 k� �c��g�%�0d  U89D"!   ��    �  }L"$_�k�DГ��<��|( ���A�9P�1�4��3��T0 k� �_��c�%�0d  U89D"!   ��    �  }L" _�k�DЏ��=��|( ���A�9P�1�8��3��T0 k� �_��c�%�0d  U89D"!   ��    �  }L"_�k�DЋ��=��|( ���A�9P�1�8��3��T0 k� �_��c�%�0d  U89D"!   ��    �  }L"_�g�DЇ�|=��|( ���A�9P�1�8��3��T0 k� �_��c�%�0d  U89D"!   ��    �  }L"_�g�DЃ�x=��|( ��A�:P�1�8��3��T0 k� �_��c�%�0d  U89D"!   ��    �  }L"_�g�D��t=��|( ��A� :P�1�8��3��T0 k� �_��c�%�0d  U89D"!   ��    �  }L"_�g�D�{�t=��|( ��A��:P�1�8��3��T0 k� �[��_�%�0d  U89D"!   ��    �  }L"_�g�D�w�p=��|( ��A��:P�1�<��3��T0 k� �[��_�%�0d  U89D"!   ��    �  }L"_�g�D�w�l>��|( ��A��:P�1�<��3��T0 k� �[��_�%�0d  U89D"!   ��    �  }L"_�c�D�s�h>��!�( ��A��:P�1�<��"���T0 k� �[��_�%�0d  U89D"!   ��    �  }L"_�c�Mpo�h>��!�( �{�A��;P�1�<��"���T0 k� �[��_�%�0d  U89D"!   ��    �  }L" _�c�Mpo�d>��!�( �{�A��;P�1�<��"���T0 k� �[��_�%�0d  U89D"!   ��    �  }L" _�c�Mpk�`>��!�( �{�A��;P�1�<��"���T0 k� �[��_�%�0d  U89D"!   ��    �  }L!�_�c�Mpg�\>��!�( �{�A��;P�1�<��"���T0 k� �W��[�%�0d  U89D"!   ��    �  }L!�_�c�Mpg�\>��!�( �{�A��;P�1�@��"���T0 k� �W��[�%�0d  U89D"!   ��    �  }L!�_�c�Mp` X>���!�( �{�A��;P�1�@��"���T0 k� �W��[�%�0d  U89D"!   ��    �  }L!�_�_�Mp` T>���!�( �{�A��<P�1�@��"���T0 k� �W��[�%�0d  U89D"!   ��    �  }L!�_�_�Mp\T?���!�( �{�A��<P|1�@��"���T0 k� �W��[�%�0d  U89D"!   ��    �  }L!�_�_�MpXP?���!�( �w�A��<Px1�@��"���T0 k� �W��[�%�0d  U89D"!   ��    �  }L�_�_�MpXL?���!�( �w�A��<Px1�@��"���T0 k� �W��[�%�0d  U89D"!   ��    �  }L�_�_�M�TL?���|( �w�A��<Pt1�@��3��T0 k� �W��[�%�0d  U89D"!   ��    �  }L�_�_�M�TH?��|( �w�A��<Pt1�@��3��T0 k� �S��W�%�0d  U89D"!   ��    �  }L�_�_�M�PD?��|( �w�A��<Pp1�D��3��T0 k� �S��W�%�0d  U89D"!   ��    �  }L�_�[�M�PD?��|( �w�A��=Pl1�D��3��T0 k� �S��W�%�0d  U89D"!   ��    �  }L�_�[�M�L@?��|( �w�A��=Pl1�D��3��T0 k� �S��W�%�0d  U89D"!   ��    �  }C��_�[�M�H@?��|( �w�A��=Ph1�D��3��T0 k� �S��W�%�0d  U89D"!   ��    �  }C��_�[�M�H<?1��|( �s�A��=Ph1�D��3��T0 k� �S��W�%�0d  U89D"!   ��    �  }C��_�[�M�D	8@1��|( �s�A��=Pd1�D��3��T0 k� �S��W�%�0d  U89D"!   ��    �  }C��_�[�M�D	8@1��|( �s�A��=P`1�D��3��T0 k� �S��W�%�0d  U89D"!   ��    �  }C��_�[�Mp@
4@1��|( �s�A��=P`1�D��3��T0 k� �S��W�%�0d  U89D"!   ��    �  }C��_�[�Mp@4@1��|( �s�A��=P\1�D��3��T0 k� �O��S�%�0d  U89D"!   ��    �  }C��_�[�Mp<0@1��!�( �s�A��>P\1�H��"s��T0 k� �O��S�%�0d  U89D"!   ��    �  }C��_�W�Mp<0@1��!�( �s�A��>PX1�H��"s��T0 k� �O��S�%�0d  U89D"!   ��    �  }C��_�W�Mp<,@1��!�( �s�A��>PX1�H��"s��T0 k� �O��S�%�0d  U89D"!   ��    �  }C��_�W�Mp8,@1��!�( �s�A��>PT1�H��"s��T0 k� �O��S�%�0d  U89D"!   ��    �  }C��_�W�Mp8�(@A��!�( �s�A��>PT1�H��"s��T0 k� �O��S�%�0d  U89D"!   ��    �  }C��_�W�Mp4�(@A��!�( �o�A��>PP1�H��"s��T0 k� �O��S�%�0d  U89D"!   ��    �  }C��_�W�Mp4�$@A��!�( �o�A��>PP1�H��"s��T0 k� �O��S�%�0d  U89D"!   ��    �  }C�_�W�D�0�$AA��!�( �o�A��>PL1�H��"s��T0 k� �O��S�%�0d  U89D"!   ��    �  }C�_�W�D�0� AA��!�( �o�A��?PL1�H��"s��T0 k� �O��S�%�0d  U89D"!   ��    �  }C�_�W�D�0� AA��!�( �o�A��?PH1�H��"s��T0 k� �K��O�%�0d  U89D"!   ��    �  }C�_�W�D�,�AA��!�( �o�A��?PH1�L��"s��T0 k� �K��O�%�0d  U89D"!   ��    �  }C�_�S�D�,�AA��|( �o�A��?PD1�L��3��T0 k� �K��O�%�0d  U89D"!   ��    �  }C�_�S�D�,�AA��|( �o�A��?PD1�L��3��T0 k� �K��O�%�0d  U89D"!   ��    �  }C�_�S�D�,�AA��|( �o�A��?P@1�L��3��T0 k� �K��O�%�0d  U89D"!   ��    �  }C�_�S�D�,�BA��|( �o�A��?P@1�L��3��T0 k� �K��O�%�0d  U89D"!   ��    �  }C�_�S�F ,BBA��|( �o�A��?P@1�L��3��T0 k� �K��O�%�0d  U89D"!   ��    �  }C�_�S�F ,BBQ��|( �o�A��?P<1�L��3��T0 k� �K��O�%�0d  U89D"!   ��    �  }D�_�S�F ,BCQ��|( �k�A��?P<1�L��3��T0 k� �K��O�%�0d  U89D"!   ��   �  }D�_�S�F ,BCQ��|( �k�A��@P81�L��3��T0 k� �K��O�%�0d  U89D"!   ��    �  }D�_�S�F ,BDQ��|( �k�A��@P81�L��3��T0 k� �K��O�%�0d  U89D"!   ��    �  }D�_�S�F ,2DQ��|( �k�A��@P81�L��3��T0 k� �K��O�%�0d  U89D"!   ��    �  }D�_�S�E�,2 EQ��|( �k�A��@P41�L��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }A��_�S�E�,2 EQ��|( �k�A��@P41�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }A��_�O�E�01�FQ��|( �k�A��@P01�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }A��_�O�E�01�GQ��|( �k�A��@P01�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }A��_�O�E�0A�GQ�|( �k�A��@P01�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }A��_�O�B�4 A�HQ�|( �k�A��@P,1�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }A�_2O�B�4!A�Ha�|( �k�A��@P,1�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }A�_2O�B�4!A�Ia�|( �k�A��@P,1�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }A�_2O�B�4!A�Ia�|( �k�A��@P(2�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }A�_2O�B�8!A�Ja�	|( �k�A��AP(2�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }A�_2O�B�8"A�Ja�|( �g�A��AP$2�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }BA�_2O�B�<"A�Ja�|( �g�A��AP$3�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }BA�_2O�B�@#A�Ja�|( �g�A��AP$3�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }BA�_2O�B�@#Q�Ka�|( �g�A��AP 3�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }BA�_2O�B�D$Q�Ka�|( �g�A��AP 3�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }BA�_2O�B�H$Q�K1�|( �g�A��AP 4�P��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }K��_2O�B�L%Q�K1�|( �g�A��AP4�T��3��T0 k� �G��K�%�0d  U89D"!   ��    �  }K��_2K�B�P%Q�L1�|( �g�A��AP4�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_2K�B�T%Q�L1�|( �g�A��AP4�T��3��T0 k� �C��G�%�0d  U89D"!   ��   �  }K��_2K�B�X&Q�L1�|( �g�A��AP5�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�B�\&Q�M1�|( �g�A��AP5�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�E�`'Q�M1� |( �g�A�|AP5�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�E�d'Q�N1�"|( �g�A�|AP5�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�E�h(Q�O1�%|( �g�A�|BP5�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�E�l)a�O1�'|( �g�A�|BP6�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�E�p)a�P!�)|( �g�A�xBP6�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�E�t*a�Q!�+|( �g�A�xBP6�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�E�x+a�Q!�-|( �g�A�xBP6�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�D�|+a�R!�/|( �g�A�xBP7�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�DЀ,a�S!�2|( �g�A�tBP7�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�DЈ-a�S!�4|( �g�A�tBP7�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�DЌ.a�T!�6|( �c�A�tBP7�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�DА/a�T!�8|( �c�A�tBP7�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�E��/a�T!�:|( �c�A�pBP8�T��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��_BK�E��0a�T!�=|( �c�A�pBP8�X��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��`BK�E��1q�T�?|( �c�A�pBP8�X��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��`BK�E��1q�T�A|( �c�A�pBP8�X��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��`BK�E��2q�T�C|( �c�A�pBP8�X��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��`BK�E��3q�U�E|( �c�A�lBP9�X��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��`BG�E��3q�U�H|( �c�A�lCP9�X��3��T0 k� �C��G�%�0d  U89D"!   ��    �  }K��`BG�B��4q�U!�J|( �c�A�lCP 9�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��`BG�B��5q�U!�L|( �c�A�lCP 9�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��`BG�B��5 ��U!�N|( �c�A�lCP 9�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��`BG�B��6 ��U!�N|( �c�A�hCP 9�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��`BG�B��7 ��U!�P|( �c�A�hC_�:�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��`BG�E��8 ��U!�P|( �c�A�hC_�:�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��aBG�E��8 ��U!�Q|( �c�A�hC_�:�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��bBG�E��9 ��U!�R|( �c�A�hC_�:�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��cBG�E��: ��U�S|( �c�A�hC_�:�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��dBG�E��; ��U�T|( �c�A�dC_�:�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��dBG�E��< ��U�T|( �c�A�dC_�;�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��eBG�E�= ��U�T|( �c�A�dC_�;�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��gBG�D�? ��U��V|( �c�A�dC_�;�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��hBG�D�@ ��U��W|( �c�A�dC_�;�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��iBG�D�@ ��U��X|( �c�A�`C_�;�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��iBG�D�$A ��U��Y|( �c�A�`C_�;�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��jBG�D�,B ��U��Y|( �c�A�`C_�<�X��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��kBG�E�4C ��U��Z|( �c�A�`C_�<�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��lBG�E�<D ��U��[|( �c�A�`C_�<�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��lBG�E�DE ��U��\|( �c�A�`C_�<�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��m2G�E�LF ��U��\|( �c�A�\D_�<�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��n2G�E�TF ��U��]|( �c�A�\D_�<�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��n2G�E�XG�U��^|( �c�A�\D_�<�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��o2G�B�`H�U��^|( �_�A�\D_�<�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��p2G�B�hI�U��_|( �_�A�\D_�=�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��p2G�B�pI�U��`|( �_�A�\D_�=�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��q�G�B�xJ�U��`|( �_�A�\D_�=�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��r�G�B��K�U��a|( �_�A�\D_�=�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��r�G�I�K�U��b|( �_�A�XD_�=�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��s�G�I�L�U��b|( �_�A�XD_�=�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��t�G�I�L�U��c|( �_�A�XD_�=�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��t2G�I�M�U��d|( �_�A�XD_�=�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��u2G�I�M�U��d|( �_�A�XD_�>�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��u2G�I!�M��U��e|( �_�A�XD_�>�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��v2C�I!�N��U��e|( �_�A�XD_�>�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }K��w2C�I!�N��U��f|( �_�A�XD_�>�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }B��w2C�I!�N��U��g|( �_�A�XD_�>�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }B��x2C�I!�N��U��g|( �_�A�TD_�>�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }B��x2C�I�O��U��h|( �_�A�TD_�>�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }B��y2C�I�O��U��h|( �_�A�TD_�>�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }B��y2C�I�O��V��i|( �_�A�TD_�>�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }B��zBC�I�O� V��i|( �_�A�TD_�>�\��3��T0 k� �?��C�%�0d  U89D"!   ��    �  }B��zBC�I�O� V��j|( �_�A�TD_�?�\��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }B��{BC�L��N�V��j|( �_�A�TD_�?�\��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��{BC�L��N�V��k|( �_�A�TD_�?�\��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��|BC�L��N�W��k|( �_�A�TD_�?�\��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��|BC�L��N�W��l|( �_�A�TD_�?�\��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��}BC�L��NW��l|( �_�A�PD_�?�\��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��}BC�L��NW��m|( �_�A�PD_�?�\��3��T0 k� �;��?�%�0d  U89D"!   ��   �  }K��~BC�L��NW��m|( �_�A�PD_�?�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��~BC�L��NW��n|( �_�A�PE_�?�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��BC�L��NW��n|( �_�A�PE_�?�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��BC�L��NX��o|( �_�A�PE_�?�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��BC�L��NX��o|( �_�A�PE_�?�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K���BC�L��NX��p|( �_�A�PE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��BC�L��NX��p|( �_�A�PE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��BC�L��NX��p|( �_�A�PE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��BC�L��NX��q|( �_�A�PE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��BC�L��NY��q|( �_�A�PE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��BC�L��NY��r|( �_�A�LE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��~BC�L��MY��r|( �_�A�LE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��~BC�L��MY��r|( �_�A�LE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��~BC�L��MY��s|( �_�A�LE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��~BC�L��M Y��s|( �_�A�LE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��}BC�L��M Y��t|( �_�A�LE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��}BC�L��M Y��t|( �_�A�LE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��}BC�L��M$Z��t|( �_�A�LE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��}BC�L��M$Z��u|( �_�A�LE_�@�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��}BC�L��M$Z��u|( �_�A�LE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��|BC�L��M$Z��u|( �_�A�LE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��|BC�L��M(Z�v|( �_�A�LE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��|BC�L��M(Z�v|( �_�A�LE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��|BC�L��M(Z�v|( �_�A�LE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }K��|BC�L��M,Z�w|( �_�A�LE_�A�`��3��T0 k� �;��?�%�0d  U89D"!   ��    �  }                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��	0 ]�$$ p �� x#H  � �
 	   � ��     xA; ��    �=�               Z }           ��    ���   0	%          ���>     
    � �j�    ���� �j�     8��             k  Z }         Q      ���   0
 	          Oô  I I      }��     Oô }��                    K	 Z }         �     ���  8

           ]n     	    ���     ]h ��     �P               [ Z }          ,��   
  ���  8          t�&   � �	   . u~     t�' u7�    �"              
 Z }          ��  (  ���   P	           Ӏ  ��     B�
��      Ӏ�
��           	                ���x                 ���    P             ��PQ    	     V �M$    ��PQ �M$                            �         w�     ��H  (	          FZ   	   j �     F *     @�w                   Y��          �p     ��@   8�           B�Y          ~��`�     B����k�     ��U              	 1��          ��     ��@   0
9
          _�         � ��-     _� ���       5               �� �         	 �p     ��@   H	$
         �Ȗc        � �P6    �Ȝ �P6    ��                    	   �         
 �     ��@   H
	!         ��I� ��     � �$t    ��I� �$t                              ���M                ��@                   ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��7  ��        � ��    ��7 ��         "                  x                j  �       �                         ��    ��        � �      ��   �           "                                                 �                          � � } � u�
 � �� � � ��� � �  
               	
  -   � �I �)�s       / ``� /� a� /� a� 0 a� �� �c@ �� d@ �d _@���. ����< ����J ����X ����  ����. ����< ����J ����X � �� u� 
�\ V� 
� V� 
�| W  
�< W� 
�\ W� � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0� ���� � � }`���� ����� � 
�� V� 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� }  ����  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    "�j�� , " �
� �  �  
� ��    ��     � �      ����  ��     � �      ��    ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �      �� � � ���        �!T ���        �        ��        �        ��        �    ��     <�� <��        ��                         �w� $  %��                                     �                  ����            �� ����%��    }�� F � $          16 Pat Verbeek son y   2:51                                                                        0  0     �cc~2� c�:Ekj3] krC �C.h �C2h �C4P �C7H � 	C;` � 
C<O �K@ � KI � KP � K> �J�i �J�a �J�a � � � �CM � C"U � � � �B� � � B� � �cV � � c^ � ~c� � c� � sc� � � c� � _c� � gc� � d c� � l !c�  J	"� � J	#� � Z$� � Z%�	 �&"� � � '"� � �(� � �)
� � �*"� } � +"� � �,"� } �-*� � �."� � � /"� � �0� � � 
� � �2� � � 
� � �4� � � 
� � � 
� � �7*6� �8*:� �9)��:*<�<;*:�\ )��?=*:_ )� �  *P�                                                                                                                                                                                                                         �� R @      �     @         �     Y P E ]  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��    ��g�� ��������������������������������������������������������   �4, 7  @� �v��                                                                                                                                                                                                                                                                                                                                                              �"@	�@                                                                                                                                                                                                                                     
     �    /    ��  D�J    	  	�  	                           ������������������������������������������������������                                                                         	                                                                 �      �                      �  �          	  
 	 
 	 	 ���������������������� ���������������������������� � ���� ���������������� ����� ������������������ ���� ������������ ���� � ����� ��� ��� �������� ������ ����������� ������� ��������  ��� �� �� ���� �������������� �������� ��                         	     '          ��  H�J                                    ������������������������������������������������������                                                                           	                                                            
       � �(          ]        �    ��              
 	  
	 
 	 	 �����  ��������� ������� ����������������� ������� ����� �������� ����� �� ��� � �  �� ��� ������������ ������������������ ������������������ ������������������������������� ���������� ���� �������� ����� ����� ��� ������� ��              �                                                                                                                                                                                                                                                                                                              �             


            �   }�                                                                                          ��������   ��������   ������������   ����������������   0��������������������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 0 I =               	                  � }�[� �\                                                                                                                                                                                                                                                                                        )n)n1n  
                            k      m            m      c                                                                                                                                                                                                                                                                                                                                                                                                                 > �  >�  J�  (�  @�  EZmX �����̎����� � �N \�̞�t����������������f�                ���� �+��        	 �   & AG� �   u                 �                                                                                                                                                                                                                                                                                                                                      p B C   �                       !��                                                                                                                                                                                                                            Y   �� �~ ��      �� B 	     ���������������������� ���������������������������� � ���� ���������������� ����� ������������������ ���� ������������ ���� � ����� ��� ��� �������� ������ ����������� ������� ��������  ��� �� �� ���� �������������� �������� �������  ��������� ������� ����������������� ������� ����� �������� ����� �� ��� � �  �� ��� ������������ ������������������ ������������������ ������������������������������� ���������� ���� �������� ����� ����� ��� ������� ��              ���������������������������������������������������f��ff�fff�ff���������l�ff�ffffl��ff˼fllf������l��̼�ʗ���˹�ffjz�fkyl�l��fƨ�����������������������̼��̉������������������������������f���f�fff�ff�ffl�ff�flfl�l��xl�wwl���l̻�����˺��fl����l�xx��w��̻���l�f�f�ƻ�fl�����ffl�ffffffff���f���̚���ffflffflfffffffffflfffff������������������������l���l������f����������������������������l��lf��f�fff�f��l˪���ww��w�����flflffffffff�̼̙��fww��w��fx�̻�llffff�ffff���fl���f�l�l�˶����fffl��fflfll����ff��ff��lfl�lf��l���l�����������l�������l�������ʼ�j˚��̩��ʨ��ɘ���xxxȈ��ɉ�x���̇�̺������www��ww��xw���x��xk�����������wx��������������x����l�ƈ��Ƈ���w��Ɨ��̩z�̩yf̪�f�������������������������������̙i���ɖ�yɌ��ˌȉ̚ə̩���ə��Ɉ����x�̹x�̹�����������ƺ�������������������ˈ������˙������̫��̺�������˪�������������̸��̗�����̇��̇�����������������������̈���xx����x���w���ɉ��̨���k���̛̻�������������l��Ʀl�Ɗl�l���̻�lk��̺�f̩�l��f�ɫ�ˉ�lɊ�˙���ʚ���˙�˫̼���ɬ�̚��̼�����̼���̬������̼�����˻������������f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff���m�    >      /     ��                       B     �   �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �f ��       p���� ��  p���� �$ ^h  ��  p  � ���                 �� �   6   
���(��   �    ����� ��   ����� �$ ^$  9   �  �� K 
]�  ����p ��  � �  � ��� �� � ��� �$  � �  �� �  �      �      �������2����   g���        f ^�         ��              ��	����2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                                    �����   �   �   �   ����                                     	�  		  	 � 	 	 	   	   	   	   	  ��                  ��   	   	   	   	   	   	 	 	 � 		  	�                 �   	    �   	    �   	    �   	   	   �  	   �  	   �  	   �                                      
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           " """ "!   " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "! ""! " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      " """ "!   " ""  !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                       ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                      ��  ��  ���     �     �                                                                                                                                                                                    �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��        �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                                   � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        k}z�gg��j�� 
�� 	�� �� �� 
�� �� ��̻�"+��" 4"  4   D   H   H   �  +  ""    ��       ��  �٠ �ڛ ̸� ̻� �̽ �̀ �ɀ ��0 ��C 4�T H�T H�D �T@ �T  �C  �0  ɚ  ��� ��� �" �"  �"�                 �� �� �� {�             �   �� � � ��� � �  ��                                        �   �   �   "   "   "  !�    ��                             �  �  �     �   �  �  �                  �   �   �   �  �  �  �  �      �     �                                                                                                                                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                  �   ��   �                            � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                                                                                                                                                                    �  ��� ݻ� g�� bm� ggz�'w���������������˛������ˊۼ�����˻������H�DH�@U�DPT�E X�T H�P H�@ Ȥ� ̻� ˘ "�� � ���/�"" �""/���               �   �                                                     �  �                      � �                       ���           �                      �  �  �          ����  �   �             ����                         � "            � "�",�"+� ",                       "  .���"    �     �                              �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                         �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �          �  � � �� ��     �         �  ���ݼ�������ک����   �   �           �   ̰  �˰                                                                                                                                                                                                  �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������              �   �   �   �  �  �  �  �                                                                                                                                                                                                   �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                 ����                                                                                                                                                                                                       	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  ��  ��  �                                �  ��  �  �  ��  �   "   "   "  �� ��                   ����������             �EU �E  
�   �               �"�!/"�  �                                     �   ���                            �   �                                                                                                  �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �   �   "   "   "  !�    ��                              �                        ���� ��� ����        �   �  ���� �   �             �   ��  ��  ��  �  �   ��  ��                                                                                                                                                                �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                          �    � �� �  �� 	  
  �  ",  ""  �"   "                      ��  ��  �          ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                                          �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqcc~2� c�:Dkj3\ krC �C.h �C2h �C4P �C7H � 	C;` � 
C<O �K@ � KI � KP � K> �J�i �J�a �J�a � � � �CM � C"U � � � �B� � � B� � �cV � � c^ � ~c� � c� � sc� � � c� � _c� � gc� � d c� � l !c�  J	"� � J	#� � Z$� � Z%�	 �&"� � � '"� � �(� � �)
� � �*"� } � +"� � �,"� } �-*� � �."� � � /"� � �0� � � 
� � �2� � � 
� � �4� � � 
� � � 
� � �7*6� �8*:� �9)��:*<�<;*:�\ )��?=*:_ )� �  *P�3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������<�K�G�T��,�[�X�Q�K� � � � � � � � � � �2�0�.�����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.�����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������/�.�7� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 