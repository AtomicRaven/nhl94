GST@�                                                           �`�                                                      �   5                       ���2�����	 ʳ����������8�������        i      #    ����                                d8<n    �  ?     2�����  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    $�j� � �$  ��
  �                                                                               ����������������������������������      ��    bb= QQ0 4 111 44            		 

                     ��� �   � �                 nn ))
         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                B  B   �  ��   @  #   �   �                                                                                'w w  )n)n
  �    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E r �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��,O{s�Q{��������� ��Q���CKץ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��*L[w�Q{��������� ��Q���CKפ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��)L[w�Q{��������� ��Q���CKף���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��'L[w�Q{��������� ��Q���CKף���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��%L[w�Q{��������� ��Q���CKע���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��#L[w�Q{��������� ��Q���CKע���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��!L[w�Q{��������� ��Q���CKס���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8�� L[w�Q{��������� ��Q���E;Ӡ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��L[w�Q{��������� ��Q���E;ӟ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��L[w�Q{��������� ��Q���E;Ӟ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��L[w�Q{���������� ��Q���E;ӝ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��L[w�Q{���������� ��Q���E;Ϝ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��L[w�Q{���������� ��Q���E;Ϝ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��L[w�Q{���������� ��Q���E;ϛ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��L[w�Q{���������� ��Q���E;Ϛ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\�Lkw�Q{���������� ��Q���E;˙���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\�Lkw�Q{���������� ��Q���I[˘���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\�Lkw�Q{���������� ��Q���I[˗���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\�
Lkw�Q{���������� ��Q���I[˖���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\�Lkw�Q���|������� ��Q���I[˕���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\�Lkw�Q��|������� ��Q���I[˕���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\�Lkw�Q��|������� ��Q���Aϕ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\�Lkw�Q��|������� ��Q���Aϕ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\�Lkw�Q��|������� ��Q���Aӕ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\��Lkw�Q��|������� ��Q���Aӕ���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\��Lkw�Q���������� ��Q���Aו���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\��Lkw�Q���������� ��Q���E�ו���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\��Lkw�Q���������� ��Q���E�ە���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8\��Lkw�U,��������� ��Q���E�ە���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�U,��������� ��Q���E�ە���^|53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�U,�|������� ��Q���E�ߕ��^|53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�U,�|������� ��Q���A[ߕ��^x53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�U,�|������� ��Q���A[ߕ�{�^x53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�U,�|��{���� ��Q���A[ߕ�{�^t53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�U,�|��{���� ��Q���A[ߕ�w�^t53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�U,�|��{���� ��Q���A[ߕ�w�^p53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�U,#�}�{���� ��Q���A�ߕ�w�^p53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E,#�}�{���� ��Q���A�ߕ�s�^l53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E,'�}�{���� ��Q���A�ߕ�s�^l53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E,'�}�{���� ��Q���A���o�^h53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E,+���{���� ��Q���A���o�^h53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E,/���{���� ��Q���A���k�^d53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E/�������� ��Q���A���k�^d53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E3�������� ��Q���A���k�^d53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E7�������� ��Q���A���g�^`53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E;�}������ ��Q���A���g�^`53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E;�}������ ��Q���A���g�^\53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E?�}������ ��Q���A���c�^\53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E�C�}������ ��Q���A���c�^X53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E�G�}������ ��Q���A���c�^X53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��Lkw�E�K�}����� ��Q���A���_�^X53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��Lkw�E�O�}����� ��Q���A���_�^T53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��Lkw�E�S�m�|��� ��Q���A���_�^T53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��Lkw�E�W�m�|��� ��Q���A���[�^T53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��Lkw�E�[�m�|��� ��Q���A���[�^P53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��Lkw�E�_�m#�|��� ��Q���A���[�^P53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��L[w�E�c�m#�|��� ��Q���A���W�^L53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��L[w�D�g�m#�|��� ��Q���A���W�^L53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��L[w�D�o�m#�|��� ��Q���A���W�^L53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��L[w�D�s�m#�|��� ��Q���A���S�^H53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��L[w�D�w�m#�|��� ��Q���A���S�^H53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��L[w�D�{�m#�|��� ��Q���A���S�^H53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8l��A�w�D��m#�|��� ��Q���A���S�^D53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8l��A�w�D܇�]#�|��� ��Q���A���O�^D53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8l��A�w�D܋�]�|��� ��Q���A���O�^D53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8l��A�w�D܏�]�|��� ��Q���A���O�^D53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8l��A�w�Dܓ�]����� ��Q���A���K�^@53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8l��A�w�Dܛ�]����� ��Q���A���K�^@53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8l��A�w�Dܟ�]����� ��Q���A���K�^@53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8l��A�w�L|��]����� ��Q���A���K�^<53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8\��A�w�L|��]����� ��Q���A���G�^<53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8\��A�w�L|��]����� ��Q���A���G�^<53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8\��A�w�L|��]����� ��Q���A���G�^853�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8\��A�w�L|��]����� ��Q���A���G�^853�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8\��A�w�L|��]��#��� ��Q���A���C�^853�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8\��A�w�L|Ö]��#��� ��Q���A���C�^853�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8���A�w�L|ǖM��#��� ��Q���A���C�^453�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8���A�w�L|ǖM��'��� ��Q���A���C�^453�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8���A�w�L|ǖM��'��� ��Q���A���C�^453�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8���A�w�L|ǖM��'��� ��Q���A���?�^453�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8���A�w�L|ǗM��'��� ��Q���A���?�^053�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8|��A�w�L|ǗM��+��� ��Q���A���?�^053�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8|��A�w�L|ǗM��+��� ��Q���A���?�^053�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8|��A�w�L�ǗM��+�"�� ��Q���A���?�^053�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8|��A�w�L�ǘM��+�"�� ��Q���A���;�^053�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8|��A�w�L�ǘ=��+�"�� ��Q���A���;�^,53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8l��A�w�L�ǘ=��/�"�� ��Q���A���;�^,53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8l��A�w�L�ǘ=��/�"�� ��Q���A���;�^,53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8l��A�w�L�ǘ=��/�"�� ��Q���A���;�^,53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8l��A�w�L�Ǚ=��/�"�� ��Q���A���7�^(53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ǚ=��3�"�� ��R��A���7�^(53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ǙM��3�"�� ��R��A���7�^(53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ǙM��3�"�� ��R��A���7�^(53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ÚM��3��� ��R��A���7�^$53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ÚM��7��� ��R��A���3�^$53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ÚM��7��� ��R��A���3�^$53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ÚM��7��� ��R��A���3�^$53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ÚM��7��� ��R��A���3�^$53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ÚM��7��� ��UK��A���3�^$53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ÛL���;��� ��UK��A���3�^ 53�T0 k� �k��o�U2d  I$1u'2Q  ��   ����8	���A�w�L�ÛL���;��� ��UK��A���/�^ 53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ÛL���;��� ��UK��A���/�^ 53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�ÛL���;��� ��UK��A���/�^ 53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Û\���;��� ��UK��A���/�^ 53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Û\���?�"�� ��UK��A���/�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ü\���?�"�� ��UK��A���/�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ü\��|?�"�� ��UK��A���/�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ü\��|?�"�� ��A��A���+�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ü���|?�"�� ��A��A���+�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ü���|?�"�� ��A��A���+�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ü���|?�"�� ��A��A���+�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ü���|C�"�� ��A��A���+�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ü����C�"�� ��A��A���+�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ü����C�"�� ��A��A���+�^53�T0 k� �k��o�U2d  I$1u'2Q  ��   ����8	���A�w�L�Ü����C�"�� ��A��A���+�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8	���A�w�L�Ü����G��� ��A��A���'�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L�Ü����G��� ��A��A���'�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L�Ü����G��� ��A��A���'�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L�Ü����K��� ��A��A���'�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L�Ü����K��� ��A��A���'�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L�Ü����O��� ��A��A���'�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L�Ý����O��� ��A��A���'�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L�Ý����S��� ��A��A���'�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L|Ý����S��� ��A��A���'�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L|Ý����W��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L|������W��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L|������[��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�L|������_��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�L|������c��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�Dܿ����c��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�Dܿ����g��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�Dܿ����k��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�Dܿ����o��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�D�Þ���s��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�D�Þ����s��� ��A��A���#�^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�D�ß����w��� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�D�ß����{��� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�D�ß������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�D�ß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�D�ß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�BLß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�BLß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�BLß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�BLß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�BLß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ß�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ß�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ß�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ�������� ��A��A����^5"��T0 k� �k��o�U2d  I$1u'2Q  ��   ����8L��A�w�A�Þ�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ�������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�Þ������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��   ����8L��A�w�A�Þ������� ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ÞM������ ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ÞM������ ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8L��A�w�A�ÞM������ ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�A�ÞM������ ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8<��A�w�A�ÞM������ ��A��A����^53�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8 �|AP��E�(H�,X
G�!�(	��Op(iB���R��
��5"s�T0 k� ��� �U2d  I$1u'2Q  ��    � < / �|C೫E�,H�0X
-G�!�(	��Op(iB���b�
��5"s�T0 k� ��� �U2d  I$1u'2Q  ��    � < . �}C௫E�,H�4X
-C�!�(	��Op(hB���b�
��5"s�T0 k� ��� �U2d  I$1u'2Q  ��    � < - �~C௫E�0H�8W
-C�!�(	��Op(hB���b�
��5"s�T0 k� ��� �U2d  I$1u'2Q  ��    � < + �~C௫E�0H�<W
-?�!�(	��Op(hB���b�
��5"s�T0 k� ��� �U2d  I$1u'2Q  ��    � < ) �C૫E�0H�@W
-?�!�(	��Op(gB���b�
� 5"s�T0 k� ��� �U2d  I$1u'2Q  ��    � < ' ��C૫AP0H�DW
-;�!�(	.��Op(gB���b�
� 5"s�T0 k� ��� �U2d  I$1u'2Q  ��    � < % ��C৫AP4H�HW
-;�!�(	.��Op(gB���b��
�5"s�T0 k� ��� �U2d  I$1u'2Q  ��    � < # �C৫AP4H�LV
-;�|(	.��Op(gB��b��
�53�T0 k� ��� �U2d  I$1u'2Q  ��    � < ! �C�AP4H�PV
-;�|(	.��Op(fB��b��
�53�T0 k� ��� �U2d  I$1u'2Q  ��    � <  �C�AP4H�TU
-;�|(	.��Op$fB��b��
�53�T0 k� ��� �U2d  I$1u'2Q  ��    � <  �C�AP4H�XU
-7�|(	��Op$fB��b��
�53�T0 k� ��� �U2d  I$1u'2Q  ��    � <  �~C�AP4H|\T
7�|(	��Op$fB��r��
�53�T0 k� ��� �U2d  I$1u'2Q  ��    � <  �~C�AP0H|`T
7�|(	��Op$eB�#�r��
�53�T0 k� ��� �U2d  I$1u'2Q  ��    � <  �~EP��AP0H|dS
7�|(	��A�$eB�'�r��
� 53�T0 k� �|�|U2d  I$1u'2Q  ��    � <  �~EP��AP0H|hS
7�|(	��A�$eB�/�r��
�(53�T0 k� �y�yU2d  I$1u'2Q  ��    � <  �}EP��C�0H|lR
7�|(	.��A�$eB�7�r��
�,53�T0 k� �w�wU2d  I$1u'2Q  ��    � <  �}EP��C�,HpQ
7�|(	/�A�$eB�;�r��
�053�T0 k� �u�uU2d  I$1u'2Q  ��    � <  �}EP��C�,HtQ
7�|(	/�A�$eB�C�r��
�853�T0 k� �t�tU2d  I$1u'2Q  ��    � <  �}EP�C�(HxP
7�|(	/�A�$eB�K�r��
�<53�T0 k� �r�rU2d  I$1u'2Q  ��    � <  �}E@{�C�(H�O
7�|(	/�A�$eB�S�r��
�@53�T0 k� �p�pU2d  I$1u'2Q  ��    � < 	 �}E@w�C�$H�N
7�|(	�A�$eB�W�r��
�H53�T0 k� �o�oU2d  I$1u'2Q  ��    � <  �}E@s�C�$H�M
7�|(	�A�$eB�_�r��
�L53�T0 k� �n�nU2d  I$1u'2Q  ��    � <  �}E@o�C� H�L
7�|(	�A�$eB�g�B��
�T53�T0 k� �m�mU2d  I$1u'2Q  ��    � <  �}E@k�C�H�L
7�|(	�AP$eB�o�B��
�X53�T0 k� ��j� jU2d  I$1u'2Q  ��    � <  �}C�c�C�H�K�7�|(	�AP$eB�w�B��
�`53�T0 k� ��h��hU2d  I$1u'2Q  ��    � <�� �}C�_�C�H��J�7�|(	/�AP$eB��B��
�h53�T0 k� ��f��fU2d  I$1u'2Q  ��    � <�� �}C�[�C�G��I�;�|(	/�AP$eB���B��
�l53�T0 k� ��e��eU2d  I$1u'2Q  ��    � <�� �}C�W�C�G��H�;�|(	/�AP$eB���	R��
�t53�T0 k� ��d��dU2d  I$1u'2Q  ��    � <�� �}C�S�C�G��G�;�|(	/�A $eI��	R��
�|53�T0 k� ��`��`U2d  I$1u'2Q  ��    � <����}IpO�C�G��F�;�|(	/�A $dI��	R��
�53�T0 k� ��]��]U2d  I$1u'2Q  ��    � <����}IpK�C�G��E�?�|(	�A $dI��	R��
�53�T0 k� ��[��[U2d  I$1u'2Q  ��    � <��� }IpK�C� G��D�?�|(	#�A  dI��	R��
�53�T0 k� ��Y� YU2d  I$1u'2Q  ��'    � <��� }IpG�E��G��D�C�|(	#�A  dI��	R��
�53�T0 k� ��X� XU2d  I$1u'2Q  ��'    � <���}IpC�E��G��C�C�|(	#�A dI��	b��
�53�T0 k� ��V��VU2d  I$1u'2Q  ��'    � <���}I�C�E��G��B�G�|(	#�A cI.��	b��
�53�T0 k� ��U��UU2d  I$1u'2Q  ��'    � <���}I�?�E��G��A�G�|(	/#�AcI.÷	b��
Ұ53�T0 k� ��T��TU2d  I$1u'2Q  ��'    � <���}I�;�E��G��@�K�|(	/#�AcI.Ƿ	b��
Ҹ53�T0 k� ��R��RU2d  I$1u'2Q  ��'    � <���}I�;�E��G��@�O�|(	/#�AbI.Ϸ	b��
��53�T0 k� ��Q��QU2d  I$1u'2Q  ��'    � <���}I�7�E��G��?�S�|(	/#�AbI.ӷ	R��
��53�T0 k� ��Q��QU2d  I$1u'2Q  ��'    � <���}C�7�E��G��>�S�|(	/#�AaI׷	R��
��53�T0 k� ��P��PU2d  I$1u'2Q  ��'    � <���}C�3�E��G��=�W�|( #�AaI۷	R��
��53�T0 k� ��P��PU2d  I$1u'2Q  ��'    � <���}C�/�E��G��=�[�|( #�A `I�	R��
��53�T0 k� ��O��OU2d  I$1u'2Q  ��'    � <���}C�+�E��G�<�_�|( #�A `I�	R��
��53�T0 k� ��N��NU2d  I$1u'2Q  ��'    � <���}C�+�E��G�;�c�|( #�A _I�	b��R�53�T0 k� ��N��NU2d  I$1u'2Q  ��'    � <���}C�'�E��H�;�g�|( #�A ^E��	b��R�53�T0 k� ��M��MU2d  I$1u'2Q  ��'    � <�� }C�#�E�H�:�k�|( #�A ^E���	b��S 53�T0 k� ��L��LU2d  I$1u'2Q  ��'    � <�� }C��E�H�$9�o�|( #�A ]E���	b��S53�T0 k� ��L��LU2d  I$1u'2Q  ��'    � <�� }C��E�H�,9�s�|( o#�A \E���	b��S53�T0 k� ��K��KU2d  I$1u'2Q  ��'    � <�� }C��E�H�08�w�|( o#�A  \E��	R��S53�T0 k� ��J��JU2d  I$1u'2Q  ��'    � <�� }C��E�I�87�{�|( o#�A/�[E��	R��S53�T0 k� ��I��IU2d  I$1u'2Q  ��'    � <��A}C��E�I�@7��|( o#�A/�ZE��	R� S$53�T0 k� ��H��HU2d  I$1u'2Q  ��'    � <��A}C��E�I�H6̓�|( o#�A/�YE��	R�S(53�T0 k� ��H��HU2d  I$1u'2Q  ��'    � <��A}C��E�I�P6	��|( o#�A?�XE��	R�S053�T0 k� ��F��FU2d  I$1u'2Q  ��'    � <��A}C��E�I�X5	��|( o#�A?�WE��2�S453�T0 k� ��D��DU2d  I$1u'2Q  ��'    � <��A}C��A��I�`4	��|( o#�A?�VE�'�2�S<53�T0 k� ��C��CU2d  I$1u'2Q  ��'    � <���}C��A��J�h4	��|( o#�A?�UE�+�2�S@53�T0 k� ��B��BU2d  I$1u'2Q  ��'    � <���}C��A��J�l3	��|( o#�A?�TE�/�2�SD53�T0 k� ��A��AU2d  I$1u'2Q  ��'    � <���}C��A�|J�t3	-��|( o#�E��SE�3�2�SH53�T0 k� ��E��EU2d  I$1u'2Q  ��'    � <���}C���A�xJ�|2	-��|( o#�E��RE�;�"�SL53�T0 k� ��H��HU2d  I$1u'2Q  ��'    � <���}C���A�tJ��2	-� |( �#�E��RE�?�"�SP53�T0 k� ��J��JU2d  I$1u'2Q  ��'    � <���}C���A�pJ��1	-� |( �#�E��QE�C�"�ST53�T0 k� ��K��KU2d  I$1u'2Q  ��'    � <���}C���EolK��1	-� |( �#�E��PE�G�"�	SX53�T0 k� ��L��LU2d  I$1u'2Q  ��'    � <���}C���EodK��0�� |( �#�E��OE�K�"�
S\53�T0 k� ��L��LU2d  I$1u'2Q  ��'    � <���}C���Eo`K��0�� |( �#�E��NE�O��S`53�T0 k� ��M��MU2d  I$1u'2Q  ��'    � <���}C���Eo\K��0�� |( �#�E߼ME�S��Sd53�T0 k� ��L��LU2d  I$1u'2Q  ��'    � <��1|C���EoXK��/��|( �#�EߴLE�W��Sh53�T0 k� ��K��KU2d  I$1u'2Q  ��'    � <��1|C��E_PL��/��|( �#�E߰LE�[��Sh53�T0 k� ��K��KU2d  I$1u'2Q  ��'    � <��1|C��E_LL��/��|( �#�EߨKE�_��Sl53�T0 k� ��J��JU2d  I$1u'2Q  ��'    � <��1|C��E_HL��/��|( �#�EߤJE�_��Sp53�T0 k� �|I��IU2d  I$1u'2Q  ��'    � <��1{C��E_@L��.��|( �#�EߜIE�c��Sp53�T0 k� �tI�xIU2d  I$1u'2Q  ��'    � <��a{C��E_<L��.��|( �#�EߔIE�g��St53�T0 k� �lH�pHU2d  I$1u'2Q  ��'    � <��azC��E_4L��.��|( �#�EߐHE�k��Sx53�T0 k� �hG�lGU2d  I$1u'2Q  ��'    � <��azC��E_0M��.M�|( �#�E߈GE�k��S|53�T0 k� �`F�dFU2d  I$1u'2Q  ��'    � <��azC��EO(M��.M�|( �#�E߀FE�o��S|53�T0 k� �XF�\FU2d  I$1u'2Q  ��'    � <��a yC�ߢEO$M��.M�|( �#�E�xFE�o��S�53�T0 k� �PE�TEU2d  I$1u'2Q  ��'    � <��Q yC�ۡEOM� /M�|( �#�E�tEE�s��S�53�T0 k� �LD�PDU2d  I$1u'2Q  ��'    � <��P�xE�ۡEOM�/M�|( �#�E�lDE�s��S�53�T0 k� �HI�LIU2d  I$1u'2Q  ��'    � <��P�xE�נEOM�/M�	|( �#�E�dDE�s��S�53�T0 k� �@L�DLU2d  I$1u'2Q  ��'    � <��P�wE�ӠEOM�/M�	|( �#�E�\CE�s��S�53�T0 k� �8O�<OU2d  I$1u'2Q  ��'    � <��P�wE�ϠEOM� 0M�
|( �#�E�TCE�w��S�53�T0 k� �0P�4PU2d  I$1u'2Q  ��'    � <����vE�˟EN�M�$0]�|( �#�E�LBE�w��S�53�T0 k� �(R�,RU2d  I$1u'2Q  ��'    � <����vE�ǟEN�L�,1]�|( �#�E�DBE�w��S�53�T0 k� � R�$RU2d  I$1u'2Q  ��'    � <����vE�ÞEN�L�41]�|( �#�E�<BE�w��S�53�T0 k� �S�SU2d  I$1u'2Q  ��'    � <����uC￞E>�L�82]�|( �#�E�8AE�w��S�53�T0 k� �T�TU2d  I$1u'2Q  ��'    � <����uC﷞E>�L�@2]�|( �#�E�0AE�w��S�53�T0 k� �T�TU2d  I$1u'2Q  ��'    � <����tC﷞E>�K�D3��|( �#�A�(AE�s��S�53�T0 k� � R�RU2d  I$1u'2Q  ��'    � <����tC﷞E>�K�L3��|( �#�A� AE�s��S�53�T0 k� ��Q��QU2d  I$1u'2Q  ��'    � <����tCﳞE>�J�P4��|( �#�A�AE�o��S�53�T0 k� ��P��PU2d  I$1u'2Q  ��'    � <�~��sCﯞE>�J�T5��|( �#�A�AE�o��S�53�T0 k� ��O��OU2d  I$1u'2Q  ��'    � <�|��sC﫞E>�I�X6��|( �#�A�AE�k��S�53�T0 k� ��N��NU2d  I$1u'2Q  ��'    � <�z��rC吏E>�I�\6��|( �#�A� AE�g�� S�53�T0 k� ��N��NU2d  I$1u'2Q  ��'    � <�w��rCCN�H�d7��|( �#�A��AE�g��!S�53�T0 k� ��N��NU2d  I$1u'2Q  ��'    � <�u�rCCN�G�h8��|( �#�A��AE�c��!S�53�T0 k� ��N��NU2d  I$1u'2Q  ��'    � <�s�qCCN�F�l:��|( �#�A��AE�_��#S�53�T0 k� ��N��NU2d  I$1u'2Q  ��' 
   � <�r�qC���CN�E�p:��|( �#�A��AE�[��#S�53�T0 k� ��M��MU2d  I$1u'2Q  ��' 
   � <�q�pC���CN�E�p:�� |( �#�A��AE�W��$S�53�T0 k� ��M��MU2d  I$1u'2Q  ��' 
   � <�o�pC���CN�F�p:��"|( �#�A��AE�W��$S�53�T0 k� ��M��MU2d  I$1u'2Q  ��' 
   � <�m�pC���CN�F�p:��$|( �#�A��AE�S��%S�53�T0 k� ��M��MU2d  I$1u'2Q  ��' 
   � <�m�oC��CN�F^l:��%|( �#�A��AE�O��%S�53�T0 k� ��M��MU2d  I$1u'2Q  ��' 
   � <�l�oC�{�CN�G^l:��'|( �#�A��@D�O��&S�53�T0 k� ��M��MU2d  I$1u'2Q  ��' 
   � <�k��oC�w�E>�G^h:��(|( �#�A��@D�K��'S�53�T0 k� ��M��MU2d  I$1u'2Q  ��' 
   � <�j �nC�w�E>�G^h:��*|( �#�E^�@D�G��'S�53�T0 k� ��F��FU2d  I$1u'2Q  ��' 
   � <�i |nC�s�E>�G^d9��,|( �#�E^�@D�G��(S�53�T0 k� ��B��BU2d  I$1u'2Q  ��' 
   � <�h tnC�o�E>�G�d9��-|( �#�E^�@D�C��(S�53�T0 k� ��?��?U2d  I$1u'2Q  ��' 
   � <�g lnC�k�E>�G�`9��/|( �#�E^�?D�?��)S�53�T0 k� ��<��<U2d  I$1u'2Q  ��' 
   � <�f dmDk�E>�G�`8��0|( �#�E^�?D�;��)S�53�T0 k� ��9��9U2d  I$1u'2Q  ��' 
   � <�e `mDg�E��G�\8��2|( �#�E^�?D�;��*S�53�T0 k� ��8��8U2d  I$1u'2Q  ��' 
   � <�d XmDc�E�|G�X8��3|( �#�E^�?D�7��*S�53�T0 k� ��7��7U2d  I$1u'2Q  ��' 
   � <�c PlD_�E�xG�X7��5|( �#�E^�?D�3��+S�53�T0 k� ��6��6U2d  I$1u'2Q  ��' 
   � <�b HlDW�E�tG>T7��6|( �#�E^�?D�/��+S�53�T0 k� ��6��6U2d  I$1u'2Q  ��' 
   � <�a @lDS�E�pG>P6��7|( �#�E^�?D�/� +S�53�T0 k� ��6��6U2d  I$1u'2Q  ��' 
   � <�` 8lDS�E�hG>P6��9|( �#�EN�>Eo+� ,S�53�T0 k� ��2��2U2d  I$1u'2Q  ��' 
   � <�_0kDO�E�dG>L5��:|( �#�EN�>Eo'� c ,��53�T0 k� �|0��0U2d  I$1u'2Q  ��' 
   � <�^(kDK�E�`G>H5��;|( �#�EN�=Eo#� c -��53�T0 k� �x.�|.U2d  I$1u'2Q  ��' 
   � <�] kDC�E�\F^D4��=|( �#�EN�=Eo� c -��53�T0 k� �p,�t,U2d  I$1u'2Q  ��' 
   � <�\kD?�E�XF^@4��>|( �#�EN�<Eo� c .��53�T0 k� �l+�p+U2d  I$1u'2Q  ��' 
   � <�[jD3�C�LF^83��@|( �#�EN�;Eo��/��53�T0 k� �`)�d)U2d  I$1u'2Q  ��' 
   � <�Y jD3�C�HE^42��B|(#�A|;Eo��0��53�T0 k� �P(�T(U2d  I$1u'2Q  ��' 	   � <�W�jD/�C�@E^,2��C|(#�Ax:Eo��1��53�T0 k� �H'�L'U2d  I$1u'2Q  ��' 	   � <�U�iD'�C�<E�(2��D|(#�Ap9Eo��2��53�T0 k� �<'�@'U2d  I$1u'2Q  ��' 	   � <�S�iD#�C�4E�$1��E|(#�Al9D?��2��53�T0 k� �4&�8&U2d  I$1u'2Q  ��' 	   � <�Q�iD�C�0E� 1��E|(#�Ad8D>���3��53�T0 k� �,%�0%U2d  I$1u'2Q  ��' 	   � <�O��iD�EN(D�0��F|(_#�A`7D>���4��53�T0 k� �$$�($U2d  I$1u'2Q  ��' 	   � <�M��iD�EN$D�0��G|(_#�AX6D>���5��53�T0 k� � #�$#U2d  I$1u'2Q  ��' 	   � <�K��hD�END^0��H|(_#�AP5D>���6��53�T0 k� �#�#U2d  I$1u'2Q  ��' 	   � <�I�hD��ENC^/�H|(_#�AL5D>��7��53�T0 k� �"�"U2d  I$1u'2Q  ��' 	   � <�G�hC��ENC]�.��J|(��A<3D>��9��53�T0 k� � � U2d  I$1u'2Q  ��' 	   � <�FߤhC��ENB]�.��J|(��A<3D>�� :�53�T0 k� ��� U2d  I$1u'2Q  ��' 	   � <�EߜgC��EN B]�.��K|(��A.82D>ߓ� ;�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�DߔgC�ۥEM�A]�-��K|(��A.01D>ה� <�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�CߌgC�ӥEM�AM�-��K|(��A.,0D>Ӕ��<�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�B߄fC�˦EM�@M�-��K|(��A.$/DNϕ��=�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�A�xfC�ǦEM�@M�,��L|(��A..DNϕ��>�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�@�pfCE=�?M�,��L|(��A.-DN˕��?�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�?�`eCE=�>M�,��L|(��A.+DN����A�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�>�XdCE=�=M�,��L|(��Gn )DN����A�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�=?PdCE=�<M�,��L|(��Gm�(DN����B�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�<?HdC���E=�<M�+m�L|,���Gm�'DN����C�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�;?@cC���E=�<M�+m�L|,���Gm�&DN����D�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�:?8cC���E=�;M�+m�K|,���Gm�%DN����E�53�T0 k� ����U2d  I$1u'2Q  ��' 	   � <�9?(aC�w�CM�;M�*m|K|0���Gm�#DN����F|53�T0 k� ����U2d  I$1u'2Q  ��'    � <�8? aENo�CM�:=�*mxK|0���G]�"D^����Gx53�T0 k� ����U2d  I$1u'2Q  ��'    � <�8?`ENg�CM�:=x)mtJ|4���G]�!D^����Ht53�T0 k� ����U2d  I$1u'2Q  ��'    � <�8?`ENc�CM�9=p)mpJ|4��G]� D^����Hl53�T0 k� ����U2d  I$1u'2Q  ��'    � <�8?_EN[�CM�8=h)mhJ|4��G]�D^���Id53�T0 k� ����U2d  I$1u'2Q  ��'    � <�8>�^ENK�CM�7�X)m`I|8��G]�D^s���JX53�T0 k� ����U2d  I$1u'2Q  ��'    � <�8N�]ENC�CM�6�P)=\H|8��GM�D^s�2�JT53�T0 k� ����U2d  I$1u'2Q  ��'    � <�8N�]EN7�CM�5�H)=XH|8��GM�D^k�2�KL53�T0 k� ����U2d  I$1u'2Q  ��'    � <�8N�\EN/�CM�4�@)=TG|<��GM�D^g�2�KD53�T0 k� ��
��
U2d  I$1u'2Q  ��'    � <�8N�[EN'�CM�3�8)=PG|<��GM�D^_�2�K<53�T0 k� �x	�|	U2d  I$1u'2Q  ��'    � <�8N�[C��CM�2�0)=HF|<��GM�D^[�2�L853�T0 k� �t�xU2d  I$1u'2Q  ��'    � <�8N�YC��C]x0� )=@E|<��GM�DnK�2�L(53�T0 k� �h�lU2d  I$1u'2Q  ��'    � <�8N�YC��C]t/�)=<D|@��GM�DnG�2�L� 53�T0 k� �d�hU2d  I$1u'2Q  ��'    � <�8N�XC��C]l.�)=4C|@��GM�Dn?�B�L�53�T0 k� �`�dU2d  I$1u'2Q  ��'    � <�8N�WEM��C]h-�*=0C|@��GM�Dn7�B�M�53�T0 k� �\�`U2d  I$1u'2Q  ��'    � <�8N�VEM�C]d*� *=,B|@��G]|Dn3�B�M�53�T0 k� �T�XU2d  I$1u'2Q  ��'    � <�8^�VEM�C=`'<�*=$A|D��G]xDn+�B�M� 53�T0 k� �P�TU2d  I$1u'2Q  ��'    � <�8^�TEM۱C=X"<�+M?|Ds�G]pDn�BxM��53�T0 k� �H�LU2d  I$1u'2Q  ��'    � ;�8^�SEMӱC=X"<�,M>|Dk�G]lDn�BtL��53�T0 k� �D �H U2d  I$1u'2Q  �'    � :�8^xREM˱C=P <�-M=|Dc�GmhDn�BlL��53�T0 k� �C��G�U2d  I$1u'2Q  ��'    � 9�8�pQEMñO=L<�-M<|D[�GmdD>�BhL��53�T0 k� �?��C�U2d  I$1u'2Q  ��'    � 8�8�hQEͻ�O=HL�.M;|HS�GmdD>�B`L��53�T0 k� �?��C�U2d  I$1u'2Q  ��'    � 7�8�XOEͫ�O=<L�0�;|H�C�Gm\
D=�BTK�53�T0 k� ����U2d  I$1u'2Q  �'    � 5�8�TNEͣ�O=8L�0� :|H�;�G}X	D=�RPK�53�T0 k� �����U2d  I$1u'2Q  ��/    � 3�8�LME͛�O=0L�1��9|H�3�G}XD=�RHK�53�T0 k� ������U2d  I$1u'2Q  ��/    � 1�8�DLE͓�O=,<�1��8|H�+�G}TD=߷RDJ�53�T0 k� ������U2d  I$1u'2Q  ��/    � /�8�4JE̓�O= <�3��6|H��G}LD=ϹR4J�53�T0 k� ������U2d  I$1u'2Q  ��/    � .�8n,JE�{�O=<�3��5|H��G�LD=˺R0I�53�T0 k� ������U2d  I$1u'2Q  ��/    � -�8n$IE�s�O=<�4��4�H��G�HD=üR(I�53�T0 k� ������U2d  I$1u'2Q  ��/    � ,�8nHE�k�O=<�4��3�H	���G�D D=��R I�x53�T0 k� �o��s�U2d  I$1u'2Q  �/    � +�8nGE�c�O=<|5��2�H	���G�G�DM��RI�p53�T0 k� �o��s�U2d  I$1u'2Q  ��/    � *�8nFE�[�O=
<x6��1�H 	���G�C�DM��RH�h53�T0 k� �k��o�U2d  I$1u'2Q  ��/    � )�8nEE�S�O=	<p7��/�H 	���G�?�DM��RH�`53�T0 k� �k��o�U2d  I$1u'2Q  ��/    � (�8m�CE�G�O<�,`8��-�D 	���G�;�DM����GP53�T0 k� �g��k�U2d  I$1u'2Q  ��/    � &�8m�BE�?�O<�,\9��+�D 	���G�7�Em����GH53�T0 k� �c��g�U2d  I$1u'2Q  ��/    � %�8m�AE�7�O<�,T:��*�D 	���G�7�Em����G@53�T0 k� �c��g�U2d  I$1u'2Q  ��/    � $�8]�@E�/�O<�,P;��(�G�	���G�3�Em����G453�T0 k� �c��g�U2d  I$1u'2Q  ��/    � #�8]�?E�'�O<�,H<��'�G�	���G�/�Em���F,5"s�T0 k� �_��c�U2d  I$1u'2Q  ��/    � "�8]�=E��O<��,<>��$�G�	���G�+�Emo���F5"s�T0 k� �[��_�U2d  I$1u'2Q  ��/    �  �8]�<E��O<��,8?��"�G�	���G�+�Emk���F5"s�T0 k� �[��_�U2d  I$1u'2Q  ��/    � �8]�;E��O<��,4@�� �G�	���G�'�Emc��E5"s�T0 k� �W��[�U2d  I$1u'2Q  ��/    � �8]�:E���E<��,0A���G�	���G�'�E][��E5"s�T0 k� �W��[�U2d  I$1u'2Q  ��/    � �8]�9E���E<��,(B���G�	���G�#�E]W��E�5"s�T0 k� �S��W�U2d  I$1u'2Q  ��/    � �8]�9E��E<��,$C���G�	���G��E]O��E�5"s�T0 k� �S��W�U2d  I$1u'2Q  ��/    � �8]�7E�߫E<��,E���G�	���G��E]?��D�5"s�T0 k� �O��S�U2d  I$1u'2Q  ��/    � �8]�6E�׫E<��F���C�	���E��E];��D�5"s�T0 k� �K��O�U2d  I$1u'2Q  ��/    � �8]�5E�ϫE<��G���C�	���E��E]3��D�53�T0 k� �K��O�U2d  I$1u'2Q  ��/    � �8M|4E�ǫE<��H���C�	���E��E]+��|C�53�T0 k� �G��K�U2d  I$1u'2Q  ��/    � �8Mt4E쿪E<��I���C�	���E��C�#��pC�53�T0 k� �G��K�U2d  I$1u'2Q  ��/    � �8Md2E쯪E<��K���C�	�{�E��C�#��`B�53�T0 k� �C��G�U2d  I$1u'2Q  ��/    � �8M\2E짪E,��L��
�C�	�w�E��C���XB�53�T0 k� �C��G�U2d  I$1u'2Q  ��/    � �8MT1E쟫E,��M���C�	�w�E���C���PB�53�T0 k� �?��C�U2d  I$1u'2Q  ��/    � �8ML1E엫E,��N���C�	�s�E���C���HA�53�T0 k� �?��C�U2d  I$1u'2Q  ��/    � �8MD0E���E,��O���C�	�o�E���C���@A�53�T0 k� �;��?�U2d  I$1u'2Q  ��/    � �8M4/E���E,���Q�� �C�	�k�C���C���10@�|53�T0 k� �7��;�U2d  I$1u'2Q  ��/ 	   � �8M,/E�{�E,���R����C�	�k�C���C���1(?�t5"��T0 k� �7��;�U2d  I$1u'2Q  ��/ 	   � �8M$/E�s�E,���S����C�	�g�C���C���1 ?�l5"��T0 k� �3��7�U2d  I$1u'2Q  ��/ 	   � �8=/E�k�E,���S���|C�	�g�C���C���1>�d5"��T0 k� �3��7�U2d  I$1u'2Q  �/ 	   � 
�8=/E�c�Q\���T���|?�	�c�C���C���1>�\5"��T0 k� �3��7�U2d  I$1u'2Q  ��/ 	   � 	�8=.E�W�Q\���U��|?�	�_�C���O\��1=�L5"��T0 k� �/��3�U2d  I$1u'2Q  ��/ 	   � �8<�.E�O�Q\���V��|?�	�_�Cܻ�O\��0�<�D5"��T0 k� �+��/�U2d  I$1u'2Q  ��/ 	   � �8<�/E�G�Q\�|V�{��;�	�_�Cܻ�O\��0�<�85"��T0 k� �+��/�U2d  I$1u'2Q  �/ 	   � �8<�/E�C�Q\w�|W�w��;�	�_�Cܳ�O\��0�;�05"��T0 k� �'��+�U2d  I$1u'2Q  ��/ 	   � �8<�/E�;�Q\s�|W�o��7�	�[�Cܯ�O\��0�:�(5"��T0 k� �'��+�U2d  I$1u'2Q  ��/ 	   � �8<�/F/�Q\g�|X�c��3�	�[�O\��O\��0�9�5"��T0 k� �3��7�U2d  I$1u'2Q  ��    ����8<�0F'�Ql_�|X�_��3�	�[�O\��O\��@�8�53�T0 k� �7��;�U2d  I$1u'2Q  ��    ����8<�0F#�Ql[��X�W��/�	�[�O\��O\��@�8�53�T0 k� �;��?�U2d  I$1u'2Q  ��    ����8<�0F�QlW��X�S��+�	�[�O\��O\��@�7� 53�T0 k� �;��?�U2d  I$1u'2Q  ��    ����8<�1@��QlK��X�G��'�	�[�O\��O\��@�6��53�T0 k� �#��'�U2d  I$1u'2Q  ��    ����8,�2@��QlG��X�?��#�	�[�O\��O\��@�5��53�T0 k� ����U2d  I$1u'2Q  ��    ����8,�2@��Ql?��W�;���	�[�O\��O\��@�5 �53�T0 k� ����U2d  I$1u'2Q  ��    ����8,�3@���Q|;��W�3���	�[�O\�O\��@�4 �53�T0 k� �����U2d  I$1u'2Q  ��    ����8,�3@���Q|7��W�/���	�[�O\{�O\��@�3 �53�T0 k� ������U2d  I$1u'2Q  ��   ����8,�5I[�Q|+��V�#����[�O\s�O\w�@�2 �53�T0 k� ����U2d  I$1u'2Q  ��    ����8,�5I[�Q|'��V�����[�O\o�O\s�Px1 �53�T0 k� ����U2d  I$1u'2Q  ��    ����8,�6I[�Q|#��U�����[�O\k�O\o�Pp0 �53�T0 k� ����U2d  I$1u'2Q  ��    ����8,�7I[�Q|��U�����[�O\g�O\k�Ph0 �53�T0 k� �ߨ��U2d  I$1u'2Q  ��    ����8,|8I[߸Q|��T�����[�O\_�O\g�P`/ �53�T0 k� �ר�ۨU2d  I$1u'2Q  ��    ����8,t9E�׸Q|��S�����[�O\W�O\_�PP- �53�T0 k� �˦�ϦU2d  I$1u'2Q  ��    ����8,p:E�ϸQ|��R�����[�O\S�O\[�PH-�53�T0 k� �å�ǥU2d  I$1u'2Q  ��    ����8l;E�˸Q|��Q�����[�O\S�E\W�PD,�53�T0 k� ����äU2d  I$1u'2Q  ��    ����8h<E�ǸQ|��P�����[�O\O�E\S�P<+x53�T0 k� ������U2d  I$1u'2Q  ��    ����8d=E���Q|��N����M[�O\G�E\K�P,)h53�T0 k� ������U2d  I$1u'2Q  ��    ����8`>E˻�Q{���M�����M[�C�;�E\G�`$)`53�T0 k� ������U2d  I$1u'2Q  ��    ����8\?E˷�Q{���L�����M[�C�3�E\C�`(X53�T0 k� ������U2d  I$1u'2Q  ��    ����8\@E˯�Q{���K�����M[�C�3�E\?�`'P53�T0 k� ������U2d  I$1u'2Q  ��    ����8\AE˫�Q{��J�����M[�C�+�E\?�`&H53�T0 k� ������U2d  I$1u'2Q  ��    ����8XBE;��Q{��H������[�O\�E\7�` $853�T0 k� ������U2d  I$1u'2Q  ��    ����8�XCE;��Q{��G������[�O\�E\7�o�$�,53�T0 k� ������U2d  I$1u'2Q  ��    ����8�XDE;��Q{�E������_�O\�E\3�o�#�$53�T0 k� ������U2d  I$1u'2Q  ��    ����8�TDE;��Q{�D������_�O\�E\/�o�"�53�T0 k� ������U2d  I$1u'2Q  ��    ����8�TFI[��Q{۴B������c�O[��E\'�o� �53�T0 k� ������U2d  I$1u'2Q  ��    ����8�TGI[��Q{۴@������c�O[��E\'�?��53�T0 k� ������U2d  I$1u'2Q  �    ����8XGI[��Q{׳�?����� c�O[��E\#�?�_�53�T0 k� ������U2d  I$1u'2Q  �    ����8XHI[��Q{Ӳ�>����� g�O[��E\�?�_�53�T0 k� ������U2d  I$1u'2Q  ��   ����8XIIk�Q{ϰ�;����� k�O[��E\�?�_�53�T0 k� ������U2d  I$1u'2Q  ��    ����8\JIk{�Q{˰� 9����� k�O[��E\���_�53�T0 k� �����U2d  I$1u'2Q  ��    ����8\KIk{�Q{ǯ� 8����� o�O[��A\���_�53�T0 k� �����U2d  I$1u'2Q  ��    ����8�\KIkw�Q{ˮ�$6����� o�O[��A\���_�53�T0 k� �{���U2d  I$1u'2Q  ��    ����8�`LIks�Q{˭�(5����� s�O[��A\���_�53�T0 k� �w��{�U2d  I$1u'2Q  ��    ����8�`LI[o�Q{˭�,3����� s�O[��A\���_�53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8�dMI[o�Q{ˬ�,2����� s�O[��A\���_�53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8�dMI[o�Q{˫�00����� w�O[��A\���_�53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8�hNI[o�Q{ϫ�4/����� w�O[��A[����_�53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8�lNA[s�Q{ϩ�8,����� {�O[��A[���x_�53�T0 k� �c��g�U2d  I$1u'2Q  ��    ����8|pNA[s�Q{ϩ�<*����� {�O[��A[���t_�53�T0 k� �W��[�U2d  I$1u'2Q  ��    ����8|tOA[s�Q{Ө�@(����� �O[��A[��l_�53�T0 k� �O��S�U2d  I$1u'2Q  ��    ����8|tOA[s�Q{ӧ�D'����� �O[��A[��h_�53�T0 k� �G��K�U2d  I$1u'2Q  ��    ����8|xOA[s�Q{ӧ�H%����� �EK��A[��d_�53�T0 k� �?��C�U2d  I$1u'2Q  ��    ����8|xOA�s�Q{Ӧ�L#����� ��EK��A[��\_|53�T0 k� �C��G�U2d  I$1u'2Q  ��    ����8||NA�s�Q{ץ|P"����� ��EK��A[��X_t53�T0 k� �K��O�U2d  I$1u'2Q  ��    ����8�|NA�s�Q{ץ|T ����� ��EK�A[��P_p53�T0 k� �O��S�U2d  I$1u'2Q  ��    ����8��NA�s�Q{פ|X����� ��EK{�A[��L_h53�T0 k� �O��S�U2d  I$1u'2Q  �    ����8��NA�s�Q{פ|\����� ��EKw�A[��H_d53�T0 k� �O��S�U2d  I$1u'2Q  ��    ����8��NA�s�Q{ף|`����� ��C�w�A[ߺ�D_`53�T0 k� �S��W�U2d  I$1u'2Q  ��    ����8��MA�s�Q{ۣ|d����� ��C�w�A[ߺ�<_X53�T0 k� �W��[�U2d  I$1u'2Q  ��    ����8��MA�s�Q{ۢ|h����� ��C�w�A[��8_T53�T0 k� �W��[�U2d  I$1u'2Q  ��    ����8��LA�o�Q{ۡ|h����� ��C�w�A[��4_L53�T0 k� �[��_�U2d  I$1u'2Q  ��    ����8��LA�o�Q{ۡ|l����� ��C�w�A[��0_H53�T0 k� �_��c�U2d  I$1u'2Q  ��    ����8��KD{o�Q{۠|p����� ��NKs�A[��,_D53�T0 k� �_��c�U2d  I$1u'2Q  ��    ����8��KD{o�Q{۠|t����� ��NKw�A[��$
_<53�T0 k� �c��g�U2d  I$1u'2Q  �    ����8��JD{o�Q{ߟ|x����� ��NKw�E[�� 	_853�T0 k� �g��k�U2d  I$1u'2Q  ��    ����8��ID{k�Q{ߟ||����� ��NKw�E[��	_453�T0 k� �g��k�U2d  I$1u'2Q  ��    ����8��ID{k�Q{ߞ||����� ��NK{�E[��_053�T0 k� �k��o�U2d  I$1u'2Q  ��    ����8��HO{k�Q{ߞ������� ��Q�{�E[��_(53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��GO{k�Q{ߝ������� ��Q�{�E[��_$53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8��FO{k�Q{���
����� ��Q��EK��_ 53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8��EO{k�Q{���	����� ��Q��EK��_53�T0 k� �w��{�U2d  I$1u'2Q  ��    ����8��DO{o�Q{�������� ��Q��EK��_53�T0 k� �w��{�U2d  I$1u'2Q  ��   ����8��CO{o�Q{�������� ��Q��EK�� _53�T0 k� �{���U2d  I$1u'2Q  ��    ����8��BO{o�Q{�������� ��Q��EK���_53�T0 k� �����U2d  I$1u'2Q  ��    ����8��AO{o�Q{�������� ��Q��EK���_53�T0 k� �����U2d  I$1u'2Q  ��    ����8��@O{s�Q{�������� ��Q��E;߳��_53�T0 k� ������U2d  I$1u'2Q  ��    ����8��?O{s�Q{�������� ��Q��E;߲��_ 53�T0 k� ������U2d  I$1u'2Q  ��    ����8��=O{s�Q{�������� ��Q��E;߱��^�53�T0 k� ������U2d  I$1u'2Q  ��    ����8��<O{s�Q{��� ����� ��Q���E;߰��^�53�T0 k� ������U2d  I$1u'2Q  ��    ����8��;O{s�Q{��������� ��Q���E;߯��^�53�T0 k� ������U2d  I$1u'2Q  ��    ����8��9O{s�Q{��������� ��Q���E;ۯ��^�53�T0 k� ������U2d  I$1u'2Q  ��    ����8��8O{s�Q{��������� ��Q���E;ۮ��^�53�T0 k� ������U2d  I$1u'2Q  ��    ����8��7O{s�Q{��������� ��Q���E;ۭ��^�53�T0 k� ������U2d  I$1u'2Q  ��    ����8��5O{s�Q{��������� ��Q���E;۬�� ^�53�T0 k� ������U2d  I$1u'2Q  ��    ����8��4O{s�Q{��������� ��Q���CK۫�� ^�53�T0 k� ������U2d  I$1u'2Q  ��    ����8��2O{s�Q{��������� ��Q���CK۪�� ^�53�T0 k� �{���U2d  I$1u'2Q  ��    ����8��1O{s�Q{��������� ��Q���CKש���^�53�T0 k� �w��{�U2d  I$1u'2Q  ��    ����8��/O{s�Q{��������� ��Q���CKר���^�53�T0 k� �s��w�U2d  I$1u'2Q  ��    ����8��.O{s�Q{��������� ��Q���CKק���^�53�T0 k� �o��s�U2d  I$1u'2Q  ��    ����8                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��A ]�,�,� � ����\   � �
    ��?��    ��H��?��     M          V	���8           � �    ���  0
 	         ��@4    	  ����U    ��@4���U                   ���8         l�  �  ���   0
% 
          ��Qv        �0�n    ��Y�0��                  		���8�        �     ���  8	          ��   4 4   �@�    ���x�@��    &{           ���8          � �     ���   8         ���   � �
     .�(�    ��֜�(�     C�             ���8           ��    ���  P
	
         ��8  ��       B�X�    ��8�X�                         	  �p���              �  ���    P             ��|�          V�w^�    ��|��wX�       W              
 �� �          �     ��@   (
I  
         ��͔        j��`    ������Yq    �� c                 � 7         �     ��@   8	           ���_       ~����    ��������     R )                ��        ]�  �  ��H   P	
          ���          ���Ա    ������.    ���S             ���l         	 �     ��@   Pw           5�3        �����     5�3����      �7             	   ��         
 r0     ��@    
2	          �w ��	     � ���     �w ���                              ���E               ��@      5                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         �� �  ��        ����    �� ����         "               x                j  �       �                         ��    ��       ���      ��  ��           "                                                 �                         �?���0�@�(��w�������� ������� 	   
             
  �  V_ �?�H       �d �`� �d a� Ƅ �[� Ǆ  \� �� ]  �� ]  �  ]@���X � �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ���� � � }`���� ����� ����� � � a� � �h@ �  i@���� � <� s  <�  s@ � �o� �  p�   q  ä }@ � `[� d \� �  \� �  \� GD `t� H 0u� Hd u� H� v  3� �^@ 4� _@ $� �j� %� k� #� `m@ $d n  
�\ U� 
�� V  
�| V  
�\ V� 
�� V� 
�| W                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �����8������ �  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    $�j � ��$  �
� �  �  
� ��    ��     ���      ��    ��     ���      ����  ��     ���          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �%%      �� �T ���        � �T ���        �        ��        �        ��        �   (�    5���"��        ��                         ���   �� �                                    �                 ����             �������%��  ���8                 6 Adam Burt apski e   4:03                                                                        3  3     �G � �F � �4J� �I J� �kj �5kr ���"	k~ �. 
k� � CB �CC � �C. � �C4 � �C8 � �K � � K � �B� � �B� � � B� � � B� � �B� � �C � � C � �C � � C! � �cV �c�P � c�X �c� � c� �V "� �V !"� �F"� �F#
� �V$"� �V %"� �F&"� �F'*� �8("� �8 )"� �(*� �(+
� � � ,"& s  -"D { ."R {  /" s@  "H �P 1"R �X  "K �8 3"L �P 4"R �X  "K �X  "H �X  "K �X  "K �X  "G �X  "K �X  "K �X  "K �X  "G �X  "K �X  "G �                                                                                                                                                                                                                         �� R         �    @ 
        �     f P E f  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��    �m�� ��������������������������������������������������������   �4, \� 0@���@��@��A��M�w�������                                                                                                                                                                                                                                                                                                                          ;� �@՜�m����                                                                                                                                                                                                                             f    3      �  D�J    	  "                             �������������������������������������������������������                                                                                                                                     m     ]      "                � �          	  
 	 
 	 	 ����������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� �������������������            �                   �         � �  	f�J      "  	                           ������������������������������������������������������                                                                                                                                      �  �      �        a          �S 3   �          	   	 	 �������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ����              �                                                                                                                                                                                                                                                            
                                                 �             


           �   }�                       +           R�              R�                                      ��������  'r������������  R�����������������    ��������������������  '|  'r�����������������������������ww�ww333wwwwwwww�ww�ww�ww�ww333wwww 0 I =               	                  � ��<Y �`�       �$C�T+P�4$`!                                                                                                                                                                                                                                                           )n)n
  �        c      e      `      a                        m                                                                                                                                                                                                                                                                                                                                                                                                        � � �  � ��  � @��  � 2��  � 2��  EZmR  �N b�����v�����v�����"����������D�����\������                 y � : h |        	 	 �   & AG� �  �   
              �                                                                                                                                                                                                                                                                                                                                      p B L   �     p    
             !��                                                                                                                                                                                                                            Y��   �� � ���      �� B 	     ����������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� ��������������������������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ����             $��ƺ�̼���k�̼̻�����������l���ƪ��̩��̩��̪���ʫ�k���ɻ��̼��fl�������������f�ffǶ�f�ff�{ff����l���̺���i�ff̩ffffffffff�f�f�l����������������ʩ��fl��ff��f�˻���̬��̻l�l���Ƽ�l��̶̻��l�������k���������������������l�������l�f���f�k�f�ʦf�fff�fff�j�fflfffff�flffk�ffl\fff�ffhfffjffff�ff�ffffffflfffffj�ffǈff��jlx�kfl��fk�k�f�lzf�f�fl��fl���ƗY���x�f�lll����ll�l������l�������������llll����ll�f����llll����l�ll���Ʃ�ff���lʈ��j���k���ƨ��l����y��ffff�fff��fl���h���f��������x���ffffffff�fff�ffffl�ff���jk�kj���ƹ�ffffffffkfffilff��l˛��˚�fj�l���l���j������̼��̜�����������l��������lll��������������������ș������������̙l���ƙ��̘��ƶf���������������������������������kɛ�k���f���ƺ�f�kyf�kYl��{ƻ�y��fkɦff�ffl�f�̻ffl�fff�fff��f̻�������̬l�k���̩k�̪��̙��̩�̼���̼���������������������������lȩ�Ʃ��lʚ��ʈ�lh���˫��k�����̺��������������̻�˼̼��̻�ʪ���̗��̗���x���y�������������������l�Ƭf����k������uff��ffxfff�fff˫��l��ll��l̨�f�̺�ffffffff�fff���������l�l�����lll��̼�lll�����l�l���������������l�����������̺���Ǌ��ǈ�yɈ��kw���Ɉ��lɘ�̉����X�������f��|f���f�[fƇ�lfyfffflffffffflfff�fffffffff�ffffffffffffffffflffffflffffffffffffffff$�I    C   #   -   � ��                       B     �   ����������      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��     �� p���� ���� p����5� ��         �f ��     �f �$ ^$ �@      ����� ��   �����   F���� ��  F���� �$ ^$   �  F  ��               1   �������� 
� `� �d �� `� �d �$  �5  �� � 5      �  ��   �������2���� g���  �     f ^�         �� ��            ��Av���2�������J�����      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         7v` weV "fff"O�p"��p"��p"�p3�}p-��p=��p|� }�  }�  ��  ��  ��  ��  �  �  �  �  �  "              `  eV  fff O�  ��  ��  �  �} �� �� ��  |�  }�  ��    =   }   =   =              �������}�}�}�ww~r�� ∈�������������������}�� }�� ��� ��� ����   �   �   �   �   �   �   �   C""42""#2""#2""#2""#s3342"""3333    p   p   p   p   p   p   p    ��������� ��� }�� ��  ��  ����  ��  ��  ��  ��  ��  ��  ��                          � �� ��    "               wvf wfU 7Of`w��f"�� "�p-�}p���� ��� ����x��	�� �� �� "�        f  U` f` f` �p w���� `  eV  ff  O�  ��  �� ����}�                �  �  ��  �            �  �  �   �  ��  �                     �  �  �   � `  eV  ff  O�  ��  ��  ����}���������������p	���         `  eV  ff  O�  ��  ��  ���}�     �  �  �   �  ��  �   �            ��  ��  �   ��  �   ���������������p	���                    3333UUUU                        wwww                    333333333333333333333   w  G� ws@ ws� ws$7w@wwww"                               ����������� ��� �� ��  �    `  eV  ff  O�  ��  ��  � ��}�            """"                 �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "" "  """""" "!   " ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """""" "!   " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                        "! ""! " ""  !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        �w
���̩ۚ,���+��   �   �   �   �  �  9  D3  D2 T2 DB DB �@ ��  ��  ��  �  "" ""�"!��" ��       �                w�  ��� ��� ��� ˼����ɀ�؊�˽ـ��˰��̰�̻@"���"+H�"$X�"$�@"E� U� E� D� ,˸  ��  ��  ,� "" �"" """�"!���� � �              �         �           �       �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                    �     �                                                                                                                                                                                   �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                              �  �  �          ����  �   �             ����                         � "            � "�",�"+� ",                       "  .���"    �     �                         � ���� ��   � � �                                                                                                                                   �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��           
 "� ""� ""� "                       �                             ���                         �  ��                    �����                         �     �                                       �   ���                            �   �                                                                                                                   � ̻ �ۼͺ�	ۚ����C�˽T;��UJ��ET�35J�D3T�  ̰ ̻	�̻���w������wv��wpʨ� ��� ��� ��  "�� .� "�� ��0 "          �  �  ��  �   �         �  �� ʝ ,��+� "" "��CEJ�D5J� J�  �� 
�� �  �� �+� �"" """����    �         ""�"" �  ��                /���"/�  ��                    �                                                                            �               �  �  ��  �   �   �        ��  �  �  �   �                                                                                                                                                                             ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .      �����                                        � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                           �� �����ݼڜ��ک��ک��z�	��� 
�� 
�� 	�� ̘ ɪ  ��  �  �� �� ������������ ���  � � � �� �� ������ ��                      �   ��  ��  �̰ ��� ��˰�̻��̻���������ˉ�U��EP�ET �I� ٕ  �D� �L� ��� ��" ����/�"�"�""�����                                                  �     �     �   �   �   �   �   �                           �   �                    �          �         �   �  �  �   �                                                                                                                                                                                                     �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �              "      �           �  �   �   ��  �                                        ��  "   "   "  �� ��                   ����������                                ��  ��  ���                 ��               �   ��  ���  � �    �                                                                                                                                                     �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �      �   �                                           �   � "��"!��"�"!��!� ���   �       �    �EU �E  
�   �               �"�!/"�  �                                                                                                                                                                                  �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��        �    �  �   �����������     "�"�����   �� �          ����   �       �                                   �    ���  ��                    ��  ��  ���     ��   �  ��  �  �  �         � �������������  �                                                                                                                                        �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��     ʠ "� "  ""� "� ��  ��                  �   �             ʘ ̠ "  " �"" �""  �"                      �    ���� �              �  �� ��  �    � ���                                                                                                                                                                                             	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                            �� ̽��  ��  �   �                        �  ��� ̻� ��� rbp wgz�       ����������                                                                                                                                                                                                                                                   �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �   �                                        ��  ��   �   �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwwDwwAwwA""""wwwwwwqADDGG""""wwwwwwqAqwAwG""""wwwwDDtwwwww""""wwwwwqGDADGqGGqw""""wwwwwwDqGqG""""wwwwwwwwwwwwqwwqww""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUEUUEUUUUUUTDUUUU3333DDDDAEQQDUDEUTUUUU3333DDDDUETQEUADQDEUDUUUU3333DDDDUQUUDUDEUTUUUU3333DDDDEQUEQUEUEUQEUUDUUUU3333DDDDQEEDEEEDUTEUUUU3333DDDDQUUQUUQUUQUUUDUUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(����������������� � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(����������������� 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5���������������� x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x���������������� w w x y�������H���������������������������������H������yxww����������������  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(���������������� , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,���������������� +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+���������������� 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5���������������� =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=����������������     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( ���������������� � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � ����������������� � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � ����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqG � �F � �4J� �I J� �kj �5kr ���"	k~ �. 
k� � CB �CC � �C. � �C4 � �C8 � �K � � K � �B� � �B� � � B� � � B� � �B� � �C � � C � �C � � C! � �cV �c�P � c�X �c� � c� �V "� �V !"� �F"� �F#
� �V$"� �V %"� �F&"� �F'*� �8("� �8 )"� �(*� �(+
� � � ,"& s  -"D { ."R {  /" s@  "H �P 1"R �X  "K �8 3"L �P 4"R �X  "K �X  "H �X  "K �X  "K �X  "G �X  "K �X  "K �X  "K �X  "G �X  "K �X  "G �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������#��-�G�S��8�K�K�R�_� � � � � � � � � � � �,��<�������������������������������������������C�G�X�R�K�_��C�G�R�G�V�Y�Q�O� � � � � �2�0�.�����������������������������������������!��+�J�G�S��,�[�X�Z� � � � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,��<� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� �� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�A�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                