GST@�                                                            \     �                                               c���                       �������� 
 J���������������z���        �h      #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    "�j��,  " ��
  �                                                                               ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������o  b  o   1  +    '           �                  	  7  V  	                  �  )          := �����������������������������������������������������������������������������                                �[  [   J  {�   @  #   �   �                                                                                '       )n)n1n  )�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    L�xE�L|� 	=�O��>|,���@�VM{� n�E_PI3��T0 k� �xE�|E%�0d  $RH�3!   ��     � �}L�|E�L|� 	=�O��?|,���@�VM� n�F_LI3��T0 k� �|E��E%�0d  $RH�3!   ��     � �}L�|F�L|� 	M�P��?|,���@�WM� n�F_LI3��T0 k� �|F��F%�0d  $RH�3!   ��     � �}L��F�L|� 	M�Q��?|,���@�WM� n�G_LI3��T0 k� ��F��F%�0d  $RH�3!   ��     � �}L��G�L|� 	M�R��@|,���@�WM� n�H_HI3��T0 k� ��F��F%�0d  $RH�3!   ��     � �}L~�G�L|� 	M�S��A|,���@�WM�� o I_HI3��T0 k� ��G��G%�0d  $RH�3!   ��     � �}L~�G� D�� 	M�S��B|,���@�XM�� oI_HI3��T0 k� ��G��G%�0d  $RH�3!   ��     � �}L~�HO$D�� 	=�T��C|,���@�XM�� oJ_HI3��T0 k� ��H��H%�0d  $RH�3!   ��     � �}L~�HO$D�� 	=�U� E|,���@�XM�� oJ_HI3��T0 k� ��H��H%�0d  $RH�3!   ��     � �}L~�IO(D�� 	=�U� E!�,���@�XM�� oK_HI3��T0 k� ��I��I%�0d  $RH�3!   ��     � �}L~�IO,	D�� 	=�V�F!�,���@�YM�� oK_HI3��T0 k� ��I��I%�0d  $RH�3!   ��     � �}BN�IO0	D�� 	=�W�G!�,���@�YM�� oL_HI3��T0 k� ��L��L%�0d  $RH�3!   ��     � �}BN�J�0
D�� 	M�W�G!�,���@�YM�� oM_LI3��T0 k� ��O��O%�0d  $RH�3!   ��     � �}BN�J�4D�� 	M�X�H!�,���@�YM�� oM_LI3��T0 k� ��Q��Q%�0d  $RH�3!   ��     � �}BN�K�8D�� 	M�X�I!�,���@�YM�� oN_LI3��T0 k� ��S��S%�0d  $RH�3!   ��     � �}BN�K�8D��!	M�Y�I!�,���@�ZM�� oN_LI3��T0 k� ��U��U%�0d  $RH�3!   ��     � �}BN�K�<D��!	M�Y�I!�,���@�ZM�� oO_LI3��T0 k� ��V��V%�0d  $RH�3!   ��     � �}BN�L�<D��!��Z�J!�,���@�ZM�� oP_LI3��T0 k� ��W��W%�0d  $RH�3!   ��     � �}BN�L�@D��"��Z� K!�,���@�ZM�� oP_LI3��T0 k� ��W��W%�0d  $RH�3!   ��     � �}BN�L�DD��"��[�$L!�,���@�ZM�� oQ_PI3��T0 k� ��W��W%�0d  $RH�3!   ��    � �}BN�M�DD��#��[�$M|,���@�[M�� oQ_PI3��T0 k� ��X��X%�0d  $RH�3!   ��     � �}BN�M�DD��#��\�(N|,���@�[M�� oR_PI3��T0 k� ��X��X%�0d  $RH�3!   ��     � �}BN�M�HD� #��\�,O|,���@�[M�� oS_PI3��T0 k� ��X��X%�0d  $RH�3!   ��     � �}BN�N�HD� $��]�,O|,���@�[M�� oS_PI3��T0 k� ��Y��Y%�0d  $RH�3!   ��     � �}BN�N�HD�%��]�0P|,���@�[M�� oT_PI3��T0 k� ��Y��Y%�0d  $RH�3!   ��     � �}BN�N�LD�%��]�4Q|,���@�[M�� oT_PI3��T0 k� ��Y��Y%�0d  $RH�3!   ��     � �}BN�N�LD�&��^�8R|,���@�\M�� oU_PI3��T0 k� ��Y��Y%�0d  $RH�3!   ��     � �}BN�O�LD�&��^�8R|,���@�\M�� oU_TI3��T0 k� ��Z��Z%�0d  $RH�3!   ��     � �}BN�O�LD�'��_�<S|,���@�\M�� oV_TH3��T0 k� ��Z��Z%�0d  $RH�3!   ��     � �}BN�O�LD�(��_@T|,���@�\M�� oV_TH3��T0 k� ��Z��Z%�0d  $RH�3!   ��     � �}BN�O�LD�(��`@U|,���@�\M�� oW_TH3��T0 k� ��[��[%�0d  $RH�3!   ��     � �}BN�P�LD�)��`DU|,���@�]M�� oW_TH3��T0 k� ��[��[%�0d  $RH�3!   ��     � �}BN�P�L!D�*��`HV|,���@�]M�� oX_TH3��T0 k� ��[��[%�0d  $RH�3!   ��     � �}BN�P�L"D� +��aHW|,���@�]M�� o X_TH3��T0 k� ��[��[%�0d  $RH�3!   ��     � �}BN�P�L$L}$+��aLX|,���@�]M�� o Y_TH3��T0 k� ��[��[%�0d  $RH�3!   ��     � �}BN�Q�H%L}$,��aLX|,���@�]M�� o Y_XH3��T0 k� ��\��\%�0d  $RH�3!   ��     � �}BN�Q�H&L}(-��bPY|,���@�^M�� o Z_XH3��T0 k� ��\��\%�0d  $RH�3!   ��    � �}BN�Q�H(L},.��bTY|,���@�^M�� o Z_XH3��T0 k� ��\��\%�0d  $RH�3!   ��     � �}BN�Q�D)L}0.��cTZ|,���@�^M�� o Z_XH3��T0 k� ��\��\%�0d  $RH�3!   ��     � �}BN�R�D+L}4/��cX[|,���@�^M�� o$[_XH3��T0 k� ��]��]%�0d  $RH�3!   ��     � �}BN�R�D,L}40��cX[|,���@�^M�� o$[_XH3��T0 k� ��]��]%�0d  $RH�3!   ��     � �}BN�R�@.L}80��d\\|,���@�^M�� o$\_XH3��T0 k� ��]��]%�0d  $RH�3!   ��     � �}BN�R�@0L}<1��d\]|,���@�_M�� o$\_XH3��T0 k� ��]��]%�0d  $RH�3!   ��     � �}BN�R�<1L}@2��d`]|,���@�_M�� o$]_XH3��T0 k� ��]��]%�0d  $RH�3!   ��     � �}BN�S�<3L}@2��e`^|,���@�_M�� o$]_\H3��T0 k� ��^��^%�0d  $RH�3!   ��     � �}BN�S�84L}D3��ed^|,���@�_M�� o(]_\H3��T0 k� ��^��^%�0d  $RH�3!   ��     � �}BN�S�46L}H4��ed_|,���@�_M�� o(^_\H3��T0 k� ��^��^%�0d  $RH�3!   ��     � �}BN�S�47L�H4��fh_|,���@�_M�� o(^_\H3��T0 k� ��^��^%�0d  $RH�3!   ��     � �}BN�S�09L�L5��fh`|,���@�`M�� o(__\H3��T0 k� ��^��^%�0d  $RH�3!   ��     � �}BN�T�,:L�P5��fla|,���@�`M�� o(__\H3��T0 k� ��_��_%�0d  $RH�3!   ��     � �}BN�T�(<L�P6��fla|,���@�`M�� o(__\H3��T0 k� ��_��_%�0d  $RH�3!   ��     � �}BN�T�(=L�T7��gpb|,���@�`M�� o(`_\H3��T0 k� ��_��_%�0d  $RH�3!   ��     � �}BN�T�$?L�T7��gpb|,���@�`M�� o,`_\H3��T0 k� ��_��_%�0d  $RH�3!   ��     � �}BN�T� @L�X8��gtc|,���@�`M�� o,`_\H3��T0 k� ��_��_%�0d  $RH�3!   ��     � �}BN�T�BL�\8��htc|,���@�`M�� o,a_\H3��T0 k� ��`��`%�0d  $RH�3!   ��     � �}BN�T�CL�\9��hxd|,���@�aM�� o,a_\H3��T0 k� ��`��`%�0d  $RH�3!   ��     � �}BN�T�DL�`9��hxd|,���@�aM�� o,a_`H3��T0 k� ��`��`%�0d  $RH�3!   ��     � �}BN�T�FL�`:��hxe|,���@�aM�� o,b_`H3��T0 k� ��`��`%�0d  $RH�3!   ��     � �}BN�T�GL�d:��i|e|,���@�aM�� o0b_`H3��T0 k� ��`��`%�0d  $RH�3!   ��     � �}BN�T�HL�h;��i|f|,���@�aM�� o0b_`H3��T0 k� ��`��`%�0d  $RH�3!   ��     � �}BN�T IL�h;��i�f|,���@�aM�� o0c_`H3��T0 k� ��`��`%�0d  $RH�3!   ��     � �}BN�T�KL�l<��i�f|,���@�aM�� o0c_`H3��T0 k� ��a��a%�0d  $RH�3!   ��     � �}BN�U�LL�l<��j�g|,���@�bM�� o0c_`H3��T0 k� ��a��a%�0d  $RH�3!   ��     � �}BN�U�LL�p=��j�g|,���@�bM�� o0d_`H3��T0 k� ��a��a%�0d  $RH�3!   ��     � �}BN�U�ML�p=��j�h|,���@�bM�� o4d_`H3��T0 k� ��a��a%�0d  $RH�3!   ��     � �}BN�V�ML�t>��j�h|,���@�bM�� o4d_`H3��T0 k� ��b��b%�0d  $RH�3!   ��     � �}BN�V�NL�t>��k�i|,���@�bM�� o4d_`G3��T0 k� ��b��b%�0d  $RH�3!   ��     � �}BN�W�OL�x?��k�i|,���@�bM�� o4e_`G3��T0 k� ��c��c%�0d  $RH�3!   ��     � �}BN�W�OL�x?��k�i|,���@�bM�� o4e_`G3��T0 k� ��c��c%�0d  $RH�3!   ��     � �}BN�X�PL�|@��k�j|,���@�bM�� o4e_dG3��T0 k� ��d��d%�0d  $RH�3!   ��     � �}BN�X�QL�|@��l��j|,���@�bM�� o8f_dG3��T0 k� ��d��d%�0d  $RH�3!   ��     � �}BN�Y�RL��A��l��k|,���@�cM�� o8f_dG3��T0 k� ��e��e%�0d  $RH�3!   ��     � �}BN�Z.�SL��A��l��k|,���@�cM�� o8f_dG3��T0 k� ��f��f%�0d  $RH�3!   ��     � �}BN�Z.�SL��B��l��l|,���@�cM�� o8g_dG3��T0 k� ��f��f%�0d  $RH�3!   ��     � �}BN�[.�SL��B��m��l|,���@�cM�� o8g_dG3��T0 k� ��g��g%�0d  $RH�3!   ��     � �}BN�[.�SL��B��mΔm|,���@�cM�� o8g_dG3��T0 k� ��g��g%�0d  $RH�3!   ��     � �}BN�[.�SL��C��mΘm|,���@�dM�� o8g_dG3��T0 k� ��h��h%�0d  $RH�3!   ��     � �}BN�\.�TL��C��mΘm|,���@�dM�� o<h_dG3��T0 k� ��h��h%�0d  $RH�3!   ��     � �}BN�\.�TL��D��mΘn|,���@�dM�� o<h_dG3��T0 k� ��i��i%�0d  $RH�3!   ��     � �}BN�].�UL��D��mΘn|,���@�eM�� o<h_dG3��T0 k� ��i��i%�0d  $RH�3!   ��     � �}BN�].�UL��D��nޘo|,���@�eM�� o<h_dG3��T0 k� ��i��i%�0d  $RH�3!   ��     � �}BN�^.�UL��E��nޘo|,���@�eM�� o<h_dG3��T0 k� ��j��j%�0d  $RH�3!   ��     � �}BN�^.�VL��E��nޘo|,���@�eM�� o<i_dG3��T0 k� ��j��j%�0d  $RH�3!   ��     � �}BN�^.�VL��E �nޘp|,���@�fM�� o<i_dG3��T0 k� ��k��k%�0d  $RH�3!   ��     � �}BN�_.�VL��F �nޔp|,���@�fM�� o<i_hG3��T0 k� ��k��k%�0d  $RH�3!   ��     � �}BN�_.�WL��F �nޔq|,���@�fM�� o@i_hG3��T0 k� ��k��k%�0d  $RH�3!   ��     � �}BN�_.�WL��F �nޔq|,���@�fM�� o@j_hG3��T0 k� ��l��l%�0d  $RH�3!   ��     � �}BN�`.�WL}�G �n�q|,���@�fM�� o@j_hG3��T0 k� ��l��l%�0d  $RH�3!   ��     � �}BN�`.�WL}�GM�n�r|,���@�gM�� o@j_hG3��T0 k� ��l��l%�0d  $RH�3!   ��     � �}BN�a.�XL}�GM�n�r|,���@�gM�� o@j_hG3��T0 k� ��m��m%�0d  $RH�3!   ��     � �}BN�a.�XL}�HM�n�r|,���@�gM�� o@j_hG3��T0 k� ��m��m%�0d  $RH�3!   ��     � �}BN�a.�XL}�HM�n�r|,���@�gM�� o@k_hG3��T0 k� ��n��n%�0d  $RH�3!   ��     � �}BN�b.�YL}�HM�n�r|,���@�hM�� o@k_hG3��T0 k� ��n��n%�0d  $RH�3!   ��     � �}BN�b.�YDݤI��n�r|,���@�hM�� o@k_hG3��T0 k� ��n��n%�0d  $RH�3!   ��     � �}BN�b.�YDݤI��n�r|,���@ hM�� oDk_hG3��T0 k� ��o��o%�0d  $RH�3!   ��     � �}BN�b.�YDݤI��m>�r|,���@ hM�� oDk_hG3��T0 k� ��o��o%�0d  $RH�3!   ��     � �}BN�b.�ZDݨJ��m>�s|,���@ hM�� oDl_hG3��T0 k� ��o��o%�0d  $RH�3!   ��     � �}BN�b.�ZDݨJ��m>|s|,���@ iM�� oDl_hG3��T0 k� ��o��o%�0d  $RH�3!   ��     � �}BN�b.�ZDݬK��m>xs|,���@ iM�� oDl_hG3��T0 k� ��o��o%�0d  $RH�3!   ��     � �}BN�b.�[DݬK��l>xr|,���@ iM�� oDl_hG3��T0 k� ��o��o%�0d  $RH�3!   ��     � �}BN�b.�[DݰL��l>tr|,���@ iM�� oDl_hG3��T0 k� ��p��p%�0d  $RH�3!   ��     � �}BN�b.�[DݴL��l>pr|,���@ iM�� oDl_hG3��T0 k� ��p��p%�0d  $RH�3!   ��     � �}BN�b.�[DݴM��k>lr|,���@ iM�� oDm_hG3��T0 k� ��p��p%�0d  $RH�3!   ��     � �}BN�b.�\DݸN��k>hr|,���@jM�� oDm_hG3��T0 k� ��p��p%�0d  $RH�3!   ��     � �}BN�b.�\DݼN��j>hr|,���@jM�� oDm_lG3��T0 k� ��p��p%�0d  $RH�3!   ��     � �}BN�b.�\D�O��i>dr|,���@jM�� oHm_lG3��T0 k� ��p��p%�0d  $RH�3!   ��     � �}BN�b.�\D��P��i>`q|,���@jM�� oHm_lG3��T0 k� ��p��p%�0d  $RH�3!   ��     � �}BN�b.�\D��Q��hN\q|,���@jM�� oHm_lG3��T0 k� ��p��p%�0d  $RH�3!   ��     � �}BN�b.�]D��Q��gNXq|,���@jM�� oHm_lG3��T0 k� ��p��p%�0d  $RH�3!   ��     � �}L~|b.�]D��R��gNTp|,���@kM�� oHn_lG3��T0 k� ��l��l%�0d  $RH�3!   ��     � �}L~|b.�]D��R��fNPp|,���@kM�� oHn_lG"���T0 k� ��i��i%�0d  $RH�3!   ��     � �}L~|b.�]D��S��fNLo|,���@kM�� oHn_lG"���T0 k� ��g��g%�0d  $RH�3!   ��     � �}L~|b.�^D��S��fNHo|,���@kM�� oHn_lG"���T0 k� ��f��f%�0d  $RH�3!   ��     � �}L~|b�^D��T��eN@n|,���@kM�� oHn_lG"���T0 k� �|e��e%�0d  $RH�3!   ��     � �}L~xb�^D��T��eN<n|,���@kM�� oHn_lG"���T0 k� �xd�|d%�0d  $RH�3!   ��     � �}L~xb�^D��T��eN8m|,���@lM�� oHn_lG"���T0 k� �xc�|c%�0d  $RH�3!   ��     � �}L~xb�^D��U��dN4m|,���@lM�� oHo_lG"���T0 k� �xb�|b%�0d  $RH�3!   ��     � �}L~xc�_D��U��dN0l|,���@lM�� oLo_lG"���T0 k� �xb�|b%�0d  $RH�3!   ��     � �}L~tc�_D��U��d	�0l|,���@lM�� oLo_lG"���T0 k� �tb�xb%�0d  $RH�3!   ��     � �}L~tc��_D��U��d	�0l|,���@lM�� oLo_lG"���T0 k� �tb�xb%�0d  $RH�3!   ��     � �}L~tc��_D��U��d	�0l|,���@lM�� oLo_lG"���T0 k� �tb�xb%�0d  $RH�3!   ��     � �}L~tc��_D��U��d	�0l|,���@lM�� oLo_lG3��T0 k� �tb�xb%�0d  $RH�3!   ��     � �}L~tc��_D��U��d	�0l|,���@mM�� oLo_lG3��T0 k� �tb�xb%�0d  $RH�3!   ��     � �}L�tc�`D��U��d	�0l|,���@mM�� oLp_lG3��T0 k� �tb�xb%�0d  $RH�3!   ��     � �}L�pc�`D��U��d	�,l|,���@mM�� oLp_lG3��T0 k� �pb�tb%�0d  $RH�3!   ��     � �}L�pc�`D��U��d	�,l|,���@mM�� oLp_lG3��T0 k� �pb�tb%�0d  $RH�3!   ��     � �}L�pc�`D��U��d	�,l|,���@mM�� oLp_lG3��T0 k� �pb�tb%�0d  $RH�3!   ��     � �}L�pc�`BM�U��d	�,l|,���@mM�� oLp_lG3��T0 k� �pb�tb%�0d  $RH�3!   ��     � �}L�pc�aBM�U��d	�,l|,���@mM�� oLp_lG3��T0 k� �pb�tb%�0d  $RH�3!   ��     � �}L�lc�aBM�U��d	�,l|,���@mM�� oLp_lG3��T0 k� �lb�pb%�0d  $RH�3!   ��     � �}L�lc�aBM�U��d	�,l|,���@nM�� oLp_lG3��T0 k� �lc�pc%�0d  $RH�3!   ��     � �}L�lc��aBM�U��d	�,l|,���@nM�� oLp_pG3��T0 k� �lc�pc%�0d  $RH�3!   ��    � �}L�lc��a@�U��d	�,l|,���@nM�� oLq_pG"s��T0 k� �lc�pc%�0d  $RH�3!   ��     � �}L�hc��a@�UM�d	�,l|,���@nM�� oPq_pG"s��T0 k� �hc�lc%�0d  $RH�3!   ��     � �}L�hd��a@�UM�d>,l|,���@nM�� oPq_pG"s��T0 k� �hc�lc%�0d  $RH�3!   ��    � �}L�dd��a@�UM�d>,l|,���@nM�� oPq_pG"s��T0 k� �dc�hc%�0d  $RH�3!   ��     � �}L�dd��a@�UM�d>,l|,���@nM�� oPq_pG"s��T0 k� �dc�hc%�0d  $RH�3!   ��     � �}L�dd��a@�UM�d>,l|,���@nM�� oPq_pG"s��T0 k� �`c�dc%�0d  $RH�3!   ��     � �}L�dd��a@�UM�d>(l|,���@nM�� oPq_pG"s��T0 k� �`c�dc%�0d  $RH�3!   ��     � �}L�`d��a@�UM�d>(l|,���@oM�� oPq_pG"s��T0 k� �\c�`c%�0d  $RH�3!   ��     � �}L�`d��a@�UM�d>(l|,���@oM�� oPq_pG"s��T0 k� �\c�`c%�0d  $RH�3!   ��     � �}L�`d��a@�UM�d>(l|,���@oM�� oPq_pG"s��T0 k� �Xc�\c%�0d  $RH�3!   ��     � �}L�`d�a@�UM�d�(l|,���@oM�� oPr_pG"s��T0 k� �Xc�\c%�0d  $RH�3!   ��     � �}L�`d�a@�UM�d�(l|,���@oM�� oPr_pG3��T0 k� �Tc�Xc%�0d  $RH�3!   ��     � �}L�`d�aK��UM�d�(l|,���@oM�� oPr_pG3��T0 k� �Tc�Xc%�0d  $RH�3!   ��     � �}L�`d�aK��UM�d�(l|,���@oM�� oPr_pG3��T0 k� �Tc�Xc%�0d  $RH�3!   ��     � �}L�`d�aK��UM�d�(l|,���@oM�� oPr_pG3��T0 k� �Tc�Xc%�0d  $RH�3!   ��     � �}L�`d�aK��UM�d�(l|,���@oM�� oPr_pG3��T0 k� �Tc�Xc%�0d  $RH�3!   ��     � �}L�`d�aK��UM�d�(l|,���@oM�� oPr_pG3��T0 k� �Tb�Xb%�0d  $RH�3!   ��     � �}L�`d�aK��UM�d�(l|,���@pM�� oPr_pG3��T0 k� �Tb�Xb%�0d  $RH�3!   ��     � �}L�`d�aK��UM�d�(l|,���@pM�� oPr_pG3��T0 k� �Tb�Xb%�0d  $RH�3!   ��     � �}L�`d�aK��TM�d�(l|,���@pM�� oPr_pG3��T0 k� �Tb�Xb%�0d  $RH�3!   ��     � �}L�`d�aK��TM�d�(l|,���@pM�� oTr_pG3��T0 k� �Tb�Xb%�0d  $RH�3!   ��     � �}L�`d�aK��TM�d�(l|,���@pM�� oTr_pG3��T0 k� �Tb�Xb%�0d  $RH�3!   ��     � �}L�`d�aK��TM�d�(l|,���@pM�� oTs_pG3��T0 k� �Ta�Xa%�0d  $RH�3!   ��     � �}L�`d�aK��TM�d�(l|,���@pM�� oTs_pG3��T0 k� �Ta�Xa%�0d  $RH�3!   ��     � �}L�`d�aK��TM�d�$l|,���@pM�� oTs_pG3��T0 k� �Ta�Xa%�0d  $RH�3!   ��     � �}L�`d�`K��TM�d>$l|,���@pM�� oTs_pG3��T0 k� �Ta�Xa%�0d  $RH�3!   ��     � �}L�\c�`K��TM�d>$l|,���@pM�� oTs_pG3��T0 k� �Pa�Ta%�0d  $RH�3!   ��     � �}L�\c�`K��TM�d>$l|,���@pM�� oTs_pG3��T0 k� �Pa�Ta%�0d  $RH�3!   ��     � �}L�\c�`K��TM�d>$l|,���@pM�� oTs_pG3��T0 k� �P`�T`%�0d  $RH�3!   ��     � �}L�\c�`K��TM�d>$l|,���@qM�� oTs_pG3��T0 k� �P`�T`%�0d  $RH�3!   ��     � �}L�\c�`K��TM�d> l|,���@qM�� oTs_pG3��T0 k� �P`�T`%�0d  $RH�3!   ��     � �}L�\b�`K��TM�d> l|,���@qM�� oTs_pG3��T0 k� �P`�T`%�0d  $RH�3!   ��     � �}L~Xb�`K��TM�d> l|,���@qM�� oTs_pG3��T0 k� �L`�P`%�0d  $RH�3!   ��     � �}L~Xb�`K��TM�d> l|,���@qM�� oTs_pG3��T0 k� �L_�P_%�0d  $RH�3!   ��     � �}L~Tb�`K��T}�d� l|,���@qM�� oTs_pG3��T0 k� �L_�P_%�0d  $RH�3!   ��     � �}L~Tb�_K��T}�d� l|,���@qM�� oTs_pG3��T0 k� �H_�L_%�0d  $RH�3!   ��     � �}L~Tb�_K��T}�d�l|,���@qM�� oTt_tG3��T0 k� �H_�L_%�0d  $RH�3!   ��     � �}L~Pa�_K��T}�d�l|,���@qM�� oTt_tG3��T0 k� �D_�H_%�0d  $RH�3!   ��     � �}BNPa�_K��S}�d�l|,���@qM�� oTt_tG3��T0 k� �Lb�Pb%�0d  $RH�3!   ��     � �}BNLa�^K��S}�d�l|,���@qM�� oTt_tG3��T0 k� �Pe�Te%�0d  $RH�3!   ��     � �}BNLa�^K��S}�d�l|,���@qM�� oTt_tG3��T0 k� �Tg�Xg%�0d  $RH�3!   ��     � �}BNH`�^K��S}�d�l|,���@qM�� oTt_tG3��T0 k� �Xh�\h%�0d  $RH�3!   ��    � �}BNH`�^K��S}�d�l|,���@qM�� oXt_tG3��T0 k� �Xh�\h%�0d  $RH�3!   ��     � �}BND`�^K��S}�d�l|,���@qM�� oXt_tG3��T0 k� �Xi�\i%�0d  $RH�3!   ��     � �}BND_��]K��S}�d�l|,���@rM�� oXt_tG3��T0 k� �Xj�\j%�0d  $RH�3!   ��     � �}BN@_��]K��S}�d�l|,���@rM�� oXt_tG3��T0 k� �Xj�\j%�0d  $RH�3!   ��     � �}BN@_��]K��S}�d�k|,���@rM�� oXt_tG3��T0 k� �Tj�Xj%�0d  $RH�3!   ��     � �}BN<^��]K��S}�c^k|,���@rM�� oXt_tG3��T0 k� �Tj�Xj%�0d  $RH�3!   ��     � �}BN8^�|\K��S��c^k|,���@rM�� oXt_tG3��T0 k� �Pi�Ti%�0d  $RH�3!   ��     � �}BN8^�x\K��S��c^k|,���@rM�� oXt_tG3��T0 k� �Li�Pi%�0d  $RH�3!   ��     � �}BN4]�t\K��R��c^k|,���@rM�� oXt_tG3��T0 k� �Lh�Ph%�0d  $RH�3!   ��     � �}BN4]�t\K��R��c^k|,���@rM�� oXt_tG3��T0 k� �Hh�Lh%�0d  $RH�3!   ��     � �}BN0]�p[K��R��c^k|,���@rM�� oXt_tG3��T0 k� �Hh�Lh%�0d  $RH�3!   ��     � �}BN,\�l[K��R��c^k|,���@rM�� oXt_tG3��T0 k� �Dg�Hg%�0d  $RH�3!   ��     � �}BN,\�l[K��R��c^k|,���@rM�� oXu_tG3��T0 k� �@g�Dg%�0d  $RH�3!   ��     � �}BN(\h[K��R��c^k|,���@rM�� oXu_tG3��T0 k� �@g�Dg%�0d  $RH�3!   ��     � �}BN$[dZK��R��c^k|,���@rM�� oXu_tG3��T0 k� �<f�@f%�0d  $RH�3!   ��     � �}BN$[dZK��R��b^k|,���@rM�� oXu_tG3��T0 k� �8f�<f%�0d  $RH�3!   ��     � �}BN [`ZK��R��b^j|,���@rM�� oXu_tG3��T0 k� �4f�8f%�0d  $RH�3!   ��     � �}BNZ`ZK��R��b^j|,���@rM�� oXu_tG3��T0 k� �4e�8e%�0d  $RH�3!   ��     � �}BNZ\YK��R��b^j|,���@rM�� oXu_tG3��T0 k� �0e�4e%�0d  $RH�3!   ��     � �}BNZ\YK��R��bnj|,���@rM�� oXu_tG3��T0 k� �,e�0e%�0d  $RH�3!   ��     � �}BNYXYK��Q��bnj|,���@sM�� oXu_tG3��T0 k� �,e�0e%�0d  $RH�3!   ��     � �}BNYTYK��Q��bnj|,���@sM�� oXu_tG3��T0 k� �(d�,d%�0d  $RH�3!   ��     � �}BNYTXK��Q��bni|,���@sM�� oXu_tG3��T0 k� �$d�(d%�0d  $RH�3!   ��     � �}BNYPXK��Q��bni|,���@sM�� oXu_tG3��T0 k� �$d�(d%�0d  $RH�3!   ��     � �}BNYLXK��Q��bni|,���@sM�� oXu_tG3��T0 k� � d�$d%�0d  $RH�3!   ��     � �}BNYLXK��Q��bni|,���@sM�� oXu_tG3��T0 k� � d�$d%�0d  $RH�3!   ��     � �}BNYLXK��Q��ani|,���@sM�� oXu_tG3��T0 k� � d�$d%�0d  $RH�3!   ��     � �}BNYHWK��Q��ani|,���@sM�� oXu_tG3��T0 k� � d�$d%�0d  $RH�3!   ��     � �}BNYHWK��P��ani|,���@sM�� oXu_tG3��T0 k� �d� d%�0d  $RH�3!   ��     � �}C��`A��C�l.���|/�@��E�O����&�lE3��T0 k� ���%�0d  $RH�3!   ��6    �����C��a���C�d.���|/�@��E�G���� '�lF3��T0 k� �	��	%�0d  $RH�3!   ��6    �����C��a���C�\.�����|/�@��E�?�����'lF3��T0 k� ���%�0d  $RH�3!   ��6    �����EB�b��C�T.����|/�@��E�3������(lF3��T0 k� ����%�0d  $RH�3!   ��6    �����EB�b�s�DH.����|/�@� C�+������)lF3��T0 k� ����%�0d  $RH�3!   ��6    �����EB�c�k�D@.����|/�М C�#�����*lG3��T0 k� �|	��	%�0d  $RH�3!   ��6    �����EB�c�c�D8/��� |/�Д C������*lG3��T0 k� �t�x%�0d  $RH�3!   ��6    �����EB�c�[�D0/���|/�Ќ C������+lG3��T0 k� �h�l%�0d  $RH�3!   ��6    �����EB�c�S�D$/���|/�Є C������,lG3��T0 k� �`�d%�0d  $RH�3!   ��6    �����EB�c�K�D/���|/��x E@������-lG3��T0 k� �X�\%�0d  $RH�3!   ��6    �����C��c�?�D/���|/�@p E@������-lH3��T0 k� �P�T%�0d  $RH�3!   ��6    �����C�xd�7�D/���|/�@h E@�����.�lH3��T0 k� �H�L%�0d  $RH�3!   ��6    �����C�pd�/�D/��|/�@` E@��1���/�lH3��T0 k� �@�D%�0d  $RH�3!   ��6    �����C�hd�'�D�/�|	|/�@XE@��1{��0�lH3��T0 k� �4�8%�0d  $RH�3!   ��6    �����C�`d��D�/?�x|/�@PE@��1s�@�0�lH3��T0 k� �,�0%�0d  $RH�3!   ��6    �����C�Xd��D�/?�p|/�@HE0��1g�@�1�lI3��T0 k� �$�(%�0d  $RH�3!   ��6    �����C�Pd��D�/?�h|/�<E0��1_�@�2�lI3��T0 k� ��%�0d  $RH�3!   ��6    �����C�Hc��D�/?�d|/�4E0��1W�@�3�lI3��T0 k� ��%�0d  $RH�3!   ��6    �����C�@c���D�0?�\|/�,E0��1O�@�3�lI3��T0 k� ��� %�0d  $RH�3!   ��6    �����C�8c���D�0?�T|/�$E0��1G�@�4�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C�0c���D�0o�
P|/�E0��1?�@x5�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C�(c���D�0o�
H|/�E0��17�@p6�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C�b���D�0o�
8|/�E0��1#�@`7�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C�b0��D�0o�
4|/��E0{�A��\8�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C�b0��D�0o�,|/��E0s�A��T9�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C� a0��C�0o�$|/��E0k�A��L:�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C��a0��C�|0o�|/��E c�A��D;�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C��a0��C�t0_�|/���E [�@���<;�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C��`0��C�l0_�|/���E S�@���4<�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C��`0��C�d0_�|/���E K�@���0=�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C��`0��C�\0_� |/���E G�@���(>�lI3��T0 k� ��	��	%�0d  $RH�3!   ��6    �����C��_0�C�P1_�� |/���E�?�@��� >�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C��_0w�C�H1�|�!|/���E�7�@���?�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C��^0k�C�@1�x.�"|/�߼E�3�@���@�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C��^0c�C�81�p.�#|/�ߴE�+�P���@�lI3��T0 k� ����%�0d  $RH�3!   ��6    �����C��]@S�C�$1�`.�%|/�ߨ	E��P����B�lI3��T0 k� ����%�0d  $RH�3!   $�6    �����C��\@K�C�1�\.�&|/�ߠ	E��P����B�lI3��T0 k� ���%�0d  $RH�3!   ��6    �����C��\@?�C�1T.�&|/�ߘ
E��P����C�lI3��T0 k� �x�|%�0d  $RH�3!   ��6    �����C��[@7�C�1L.�'|/�_�
E��P��O�D�lI3��T0 k� �p
�t
%�0d  $RH�3!   ��6    �����C��Z@/�C�1D.�(|/�_�
E��P��O�D�lI3��T0 k� �h�l%�0d  $RH�3!   ��6    �����C��Z@'�C��1<.�(|/�_�E���P��O�E�lI3��T0 k� �d�h%�0d  $RH�3!   ��6    �����C�xY@�C��14.�)|/�_xE���P�O�F�lI3��T0 k� �\�`%�0d  $RH�3!   ��6    �����C�pY@�C��1o,
N�)|/�_tE���Pw�O�G�lI3��T0 k� �T�X%�0d  $RH�3!   ��6    �����C�hX@�C��1o(
N�*|/�_lE���Po�O�G�lI3��T0 k� �L�P%�0d  $RH�3!   ��6    �����C�`W@�C��1o 
N�*|/�_dE���`g�O�H�lI3��T0 k� �D�H%�0d  $RH�3!   ��6    �����C�PV_�C��1o
Nx+|/�_PE���`W�O�J�lI3��T0 k� �0�4%�0d  $RH�3!   ��6    �����C�HU_�D �2o
Np+|/�OHE���`O�	�K�lI3��T0 k� �(�,%�0d  $RH�3!   ��6    �����C�@U_�D �2_ 
Nh+|/�O@E���`G�	�K�lI3��T0 k� � �$%�0d  $RH�3!   ��6    �����C�8T_۷D �2^�
N`+|/�O8E���`?�	�L�lI3��T0 k� ��%�0d  $RH�3!   ��6    �����C�0S_ӶD �2^�
NX+|/�O0E߻�`7�	�L�lI3��T0 k� ��%�0d  $RH�3!   ��6    �����C�,R_˵D �2^�
NL+|/�O(E߷�`/�	�M�lI3��T0 k� ��%�0d  $RH�3!   ��6    ����C�$R_��D �2^�
ND,|/� E߯�`'�	�N�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����}C�Q_��D �2^�
N<,|/�Eߧ�`�	�|N�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����{C�P_��D |2^�
^4+!�/�Eߟ�`�	�xN�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����yC�O_��D t2^�
^,+!�, Eߗ�0�	�pO�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����wC��No��D d2^�
^+!�, ��E߇�?��	�hO�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����uE��Mo��DX2^� 
^+!�, ��E��?��	dP�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����sE��Lo��DP2^� 
^+!�, ��E�w�?��	`P�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����pE��Ko�DH2^� 
^ +!�, ��E�o�?��	\P�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����nE��Jow�D@2^��
]�*!�,��E�g�?��	XP�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����kE��J_o�D82^��
]�*!�,��E�_�?��	TP�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����iE��I_g�D,2^��
]�*!�,��E�W�?��	�PP�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����fE��H__�D$2^��
]�*!�,޼E�O�?��	�LP�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����dE��G_W�D2^��
M�)|,޴E�G�?��	�HP�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����bEиG_O�D2^�
M�)|,ެE�?�?��	�HP�lI3��T0 k� ����%�0d  $RH�3!   ��6    ����`EШE_;�D 3^o�
M�(|,ޜE�/�O��	�@PSlI3��T0 k� �t�x%�0d  $RH�3!   ��6    ����]C�E_3�C��3^k�
M�(|,�E�'�O��	@PSlI3��T0 k� �p�t%�0d  $RH�3!   ��6    ����[C��D_+�C��3^c��'|,�E��O��	<PSlI3��T0 k� �h�l%�0d  $RH�3!   ��6    ����YC��C_#�C��3^[��'|,�E��O��	8PSlI3��T0 k� �`
�d
%�0d  $RH�3!   ��6    ����VC��C��C��3^S��'|,�xE��O��	8PShI3��T0 k� �X�\%�0d  $RH�3!   ��6    ����TC��B��C��3^K��&|,�pE����	4P�hI3��T0 k� �L�P%�0d  $RH�3!   ��6    ����RC�|A��E_�3^C��&|,�hE������0P�hI3��T0 k� �@�D%�0d  $RH�3!   �6    ����RC�tA��E_�3^;��&|,�`E���w��0P�dI3��T0 k� .@�D%�0d  $RH�3!   ��?    ����RC�d?��E_�3N+��%!�,�PE���g��(P�`I3��T0 k� .@
�D
%�0d  $RH�3!   ��?    ����RC�\?��E_�3N#�|%!�,�HE�۳�c��$P�`I3��T0 k� .@�D%�0d  $RH�3!   ��?    ����RC�T>��E_�3N�x$!�,><Enϳ�[�� P�\I3��T0 k� .@�D%�0d  $RH�3!  ��?    ����RC�L>�ןE_�3N��t$!�,>4Enǳ�S��P�XI3��T0 k� .@�D%�0d  $RH�3!  ��?    ����RC�D=�ϟE_�3N��l#!�,>,En���K��P�XI3��T0 k� �@�D%�0d  $RH�3!  ��?    ����RC�<=�ǞE_�3N��h#!�,>$En���C��P�TI3��T0 k� �@�D%�0d  $RH�3!  ��?    ����RC�4<EO|3M���h#!�,>En���?��P�PI3��T0 k� �@�D%�0d  $RH�3!  ��?    ����RC�,;���EOt3M���d"!�,>En���7��P�LI3��T0 k� �@�D%�0d  $RH�3!  ��?    ����RC�$;���EOh3M���`"!�,>D>���/��P�HI3��T0 k� �@�D%�0d  $RH�3!  ��?    ����RC�:���EO`3M���\"!�,> D>���'�� P�DI3��T0 k� >@�D%�0d  $RH�3!  ��?    ����RC�9���EOP3=���X!|,=�D>�o���P�<I3��T0 k� >@�D%�0d  $RH�3!  ��?    ����RC�9���EOD2=���T!|,M�D>w�o���O�8I3��T0 k� >@�D%�0d  $RH�3!  ��?    ����RC��8���EO<2=���T |,M�D>k�o���O�4I3��T0 k� >@�D%�0d  $RH�3!  ��?    ����RC��8�{�EO42=���T |,M�D>c�o���O�0I3��T0 k� �@�D%�0d  $RH�3!  ��?    ����RD�7�s�C�,2=���P |,M�D>[�n����N,I3��T0 k� �@�D%�0d  $RH�3!  ��?    ����RD�7�k�C�$1=���P|,M�D>O�n����N(I3��T0 k� �<�@%�0d  $RH�3!  ��?    ����RD�6�c�C�1=���P|,M�D>G�n���N I3��T0 k� �<�@%�0d  $RH�3!   ��?    ����RD�6W�C�1M���P|,M�D>?�^���MI3��T0 k� �<�@%�0d  $RH�3!   ��?    ����RD�5O�C�0M���L|,M�D>3�^ߧ��LI3��T0 k� .<�@%�0d  $RH�3!   ��?    ����RD�4?�C��0M���L|,M�DN#�^ӥ��KI3��T0 k� .<�@%�0d  $RH�3!   /�?    ����RD�47�C��/M���L|,M�DN�^ˤ��KI3��T0 k� .<�@%�0d  $RH�3!   ��?    ����RD�4^/�E��/=x ML|,]�DN�^ã��J I3��T0 k� .<�@%�0d  $RH�3!   ��?    ����RD�3^'�E��/=pML|,]�DN�^����I�I3��T0 k� �<�@%�0d  $RH�3!   �?    ����RD�3^�E��.=lML|,]�DM��^����H�I3��T0 k� �<�@%�0d  $RH�3!   ��?    ����RD�2^�E��-=`ML|,]�E��^����F�I3��T0 k� �< �@ %�0d  $RH�3!   ��?    ����RD�1^�E޸-=X�L|,]�E����E�I3��T0 k� �<!�@!%�0d  $RH�3!   ��?    ����RD�1]��Eް-=P�L|,]�E�߼��D�I3��T0 k� �<"�@"%�0d  $RH�3!   ��?    ����RDt1]�Eި,=H�L|,]�E�ӽ�C�I3��T0 k� �<"�@"%�0d  $RH�3!   ��?    ����RDl0]�Eޠ,=D�L|,]�E�˾�B�I3��T0 k� �<#�@#%�0d  $RH�3!   ��?    ����RDd0MߐEޘ,=<�L|,]�D�ǿ���A�I3��T0 k� �<$�@$%�0d  $RH�3!   ��?    ����RD\/M׏I��,=4	�L|,m�D����{��@�I3��T0 k� �<%�@%%�0d  $RH�3!   ��?    ����RDL/MǏI�|+-4	�L|,m|D����k��>�I3��T0 k� �<&�@&%�0d  $RH�3!   ��?    ����PDD.M��I�t+-,
�L|,m|D����c��=�I3��T0 k� �@)�D)%�0d  $RH�3!   ��"    ����NC�<.M��I�l+-$�L|,mx
D����[��;�I3��T0 k� �<+�@+%�0d  $RH�3!   ��"    �  �LC�4.M��E�d*- �L|,mx
D����S��|:�I3��T0 k� �8+�<+%�0d  $RH�3!   ��"    � �KC�$-M��E�T*��L|,mxD����C��x8�I3��T0 k� �,*�0*%�0d  $RH�3!   ��"    � �JC� -M��E�L*��L|,}tD����;��x6�I"s��T0 k� �$*�(*%�0d  $RH�3!   ��"    � �IC�,M��E�D*��L|,}tE�{��3��t5�xI"s��T0 k� �*� *%�0d  $RH�3!   ��"    � �HC�,M�E�<*� �L|,}tE�s��+��t4�pI"s��T0 k� �/�/%�0d  $RH�3!   ��"    � �GC��+Mo�E�,*���L|,}pE�g����p1�`I"s��T0 k� �3�3%�0d  $RH�3!   ��"    � �FC��+Mc�E�$*���L|,}pE�_�^�~p0�XI"s��T0 k� � 6�6%�0d  $RH�3!   ��"    � �EE��+=[�E�*L��H|,}lE�[�^�~l.�PI"s��T0 k� �5�5%�0d  $RH�3!   �"    � �PE��*=S�E�*L��H|,}lE�S�^�~l-�HI"s��T0 k� �,3�03%�0d  $RH�3!   ��/    � �[E��*=C�H.+L��H|,}lE�G�]�~h)�8I"s��T0 k� �T0�X0%�0d  $RH�3!   ��/    � �fE��)=;�H-�+L�MH|,}hE�C�]�~h(�0I"s��T0 k� �l/�p/%�0d  $RH�3!   ��/    � �qI��)=3�H-�+L�ML|,}h E�;�]�~h&�(I3��T0 k� ��-��-%�0d  $RH�3!   �/    � �rI��)=+�H-�+L�ML|,}h F7�]ۇ~d$� I3��T0 k� >�-��-%�0d  $RH�3!   ��/    � �sI��)=#�H-�+L� ML|,}k�F/�]ӆ~d#�I3��T0 k� >|,��,%�0d  $RH�3!   ��/    � �sI��)=�H=�+L�!ML|,}g�F+�]˅~d!�I3��T0 k� >|,��,%�0d  $RH�3!   ��/    � �sCޤ)=�H=�+L�$}L|,}g�F�M��~\��I3��T0 k� >x+�|+%�0d  $RH�3!  ��/    � �sCޜ)=�H=�,L�&}L|,}g�F�M��~\��I3��T0 k� �x+�|+%�0d  $RH�3!  ��/    � �sCޘ(<��H=�,\�(}L|,}c�F�M��nX��I3��T0 k� �x*�|*%�0d  $RH�3!  ��/    � �sCސ(,��HM�,\�)}P|,}c�F�M��nT�I3��T0 k� �t*�x*%�0d  $RH�3!  ��/    � �sCވ',�HM�,\�+}P|,}c�F�M��nT�I3��T0 k� �t)�x)%�0d  $RH�3!  ��/    � �sO^�',�HM�,\�,mP|,}c�F�M��nP�I3��T0 k� �t)�x)%�0d  $RH�3!  ��/    � �rO^x%,ߖHM�,,�0mP|,}_�F�M��nL�I"���T0 k� .d%�h%%�0d  $RH�3!  ��     � �qO^p%,חHM�,,�2mP
|,}_�F��M{�nH�I"���T0 k� .T"�X"%�0d  $RH�3!  ��     � �pO^l$,ӘHM�,,�3mL	|,}_�F��Mo�nD�I"���T0 k� .L �P %�0d  $RH�3!  ��     � �oO^d$,ϙHM�,,�5%�L|,}_�E���Mg�nD
�I"���T0 k� .@�D%�0d  $RH�3!  ��     � �nO^`#,ǚHM�-,�7%�L|,}[�E���M_�n@�I"���T0 k� .8�<%�0d  $RH�3!  ��     � �mO^\#,ÛHM|-,�9%�L|,}[�E���=W�n<�I"���T0 k� N0�4%�0d  $RH�3!  ��     � �mO^P",��HMp-,|<%�L|,}[�E���=G�n8�I"���T0 k� N$�(%�0d  $RH�3!  ��     � �mO^H!��HMl-,x>%�H|,}[�B��=?�^4 �I"���T0 k� N� %�0d  $RH�3!  ��     � �mO^D!��HMd-,x@%�H|,}[�B��=7�^3�|I"���T0 k� N�%�0d  $RH�3!  ��     � �mO^@ ��HM`-tB%�H|,}W�B��=/�^/�tI3��T0 k� ��%�0d  $RH�3!  ��     � �mO^8 ��HMX-tC%�H|,}W�B��='�^+�lI3��T0 k� ��%�0d  $RH�3!  ��     � �mO^4��HMT-tE%�H|,}W�B��=�^'�dI3��T0 k� ��%�0d  $RH�3!  ��     � �mO^0��HMP-pG%�D|,}W�B��
=�^#�\I3��T0 k� ��%�0d  $RH�3!   ��     � �mO^,��HMH-pI%�D|,}W�B��=�^�TI3��T0 k� ��� %�0d  $RH�3!   ��     � �mO^ ��HM<.pL%�D|,}W�B��=�^�@I3��T0 k� ����%�0d  $RH�3!   /�     � �mO^��HM8.pN%�D |,}S�B��,��^�8I3��T0 k� ����%�0d  $RH�3!   ��     � �mO^���I�4.pO%�D |,}S�B��,�^�0I3��T0 k� ����%�0d  $RH�3!   ��     � �mO^���I�0.pQ%�C�|,}S�B��,�N��(I3��T0 k� ����%�0d  $RH�3!   ��     � �mI����I�,.pS%�C�|,}S�B��,�N�� I3��T0 k� ����%�0d  $RH�3!   ��     � �nI����I�$.�pT%�C�|,}S�B��,�M���I3��T0 k� ����%�0d  $RH�3!   ��     � �oI� ���I�.�pW%�C�|,}S�B��,׏M���I3��T0 k� ����%�0d  $RH�3!   ��     � �pI�����I�.�tX%�C�|,}S�B��,ӐM��� I3��T0 k� ����%�0d  $RH�3!   ��     � �pE�����I�.�tZ%�?�|,}O�B��,ϑM����I3��T0 k� ����%�0d  $RH�3!   ��     � �pE�����I�.�t[%�?�|,}O�B��,ǒM����I3��T0 k� ����%�0d  $RH�3!   ��     � �pE�����I�.�x\%�?�|,}O�B��,ÔM����I3��T0 k� ����%�0d  $RH�3!   ��     � �pE�����I�.�x]%�?�|,}O�B��,��M����I3��T0 k� ����%�0d  $RH�3!   ��     � �pE�����I�0�|_%�?�|,}O�B� ��M����I3��T0 k� ����%�0d  $RH�3!   ��     � �pE�����I�0��`%�?�|,}O�B���M����I3��T0 k� ����%�0d  $RH�3!   ��     � �pE�����I�1��a%�;�|,}O�B� ��=����I3��T0 k� ��"��"%�0d  $RH�3!   ��     � �pE�����I�1|�b%�;�|,}O�B� ��=���I3��T0 k� ��%��%%�0d  $RH�3!   ��     � �pE�����I�2|�c%�;�|,}O�B�!��=���I3��T0 k� ��'��'%�0d  $RH�3!   ��     � �pE�����E} 2|�c];�|,}K�B�!���=���I3��T0 k� ��)��)%�0d  $RH�3!   ��     � �pE����E|�3|�e]7�|,}K�B�"���M���I3��T0 k� ��*��*%�0d  $RH�3!   ��     � �pE����E|�3��e]7�|,}K�B�"���M���I3��T0 k� ��+��+%�0d  $RH�3!   ��     � �pE����E|�3��e]7�|,}K�B�"���M����I3��T0 k� ��,��,%�0d  $RH�3!   ��     � �pE��ùE��3��f]3�|,}K�B� #���M����I3��T0 k� ��-��-%�0d  $RH�3!   ��     � �pE��ǹE��3��f]3�|,}K�B�$#���M���xI3��T0 k� �|-��-%�0d  $RH�3!   ��     � �pE��ϻE��3��g]/�|,}K�B�,$���=�� hI3��T0 k� �p-�t-%�0d  $RH�3!   ��     � �pE���ӻE��3��gM+�|,}G�B�0$���=�� `I3��T0 k� �x.�|.%�0d  $RH�3!   ��     � �pE���׼E��3��gM'�|,}C�B�4%���=�� XI3��T0 k� �|.��.%�0d  $RH�3!   ��     � �pE���۽E��2��gM'�|,}C�B�<%���=�� PI3��T0 k� ��/��/%�0d  $RH�3!   ��     � �pE�x��E�2��gM�|,}?�B�D&���={�	�@I3��T0 k� �x0�|0%�0d  $RH�3!   ��     � �oE�x��E�2��gM�|,};�B�H'���-{�	�<I3��T0 k� �x0�|0%�0d  $RH�3!   �     � �pE�x��E�2��fM�|,};�B�L(���-w�	�4I3��T0 k� �|0��0%�0d  $RH�3!   ��     � �qA�x���E�2��fM�|,}7�B�P(���-w�	�0I3��T0 k� �x.�|.%�0d  $RH�3!   ��     � �rA�x���E�2��f=�|,}7�B�P)���-{�	�(I3��T0 k� �t,�x,%�0d  $RH�3!   ��     � �sA�x��J�1��e=�|,}3�B�T*���-{�	�$I3��T0 k� �p+�t+%�0d  $RH�3!   ��     � �tA�x��J�1��e=�|,}/�B�\,�����	�I3��T0 k� �l*�p*%�0d  $RH�3!   ��     � �uBMx��J�1��d=�|,}/�B�`-����	�I3��T0 k� �t*�x*%�0d  $RH�3!   ��     � �vBMx��J�1|�c=�|,}+�B�d.����	�I3��T0 k� �|*��*%�0d  $RH�3!   ��     � �wBMx�#�E��1|�c<��|,}+�B�l.����	�I3��T0 k� ��*��*%�0d  $RH�3!   ��     � �xBMx�+�E��1|�b,��|,}'�B�p/����	�I3��T0 k� ��*��*%�0d  $RH�3!   ��     � �yBMx�3�E��0|�a,��|,}'�B�t0����	� I3��T0 k� ��*��*%�0d  $RH�3!   ��     � �zBM|�C�E��0|�`,��|,}#�B��2����	��I3��T0 k� ��*��*%�0d  $RH�3!   ��     � �{F|�G�E��0|�_,��|,}�B��2õ��	��I3��T0 k� ��+��+%�0d  $RH�3!   ��     � �|F|�O�E��/l�^,��|,}�B��3�Ƕ��	��I3��T0 k� ��+��+%�0d  $RH�3!   ��     � �}F��W�E��/l�],��|,}�B��4�˶��	��I3��T0 k� ��+��+%�0d  $RH�3!   �     � �}F��g�E��.l�[���|,}�B��5�Ӹ��	��I3��T0 k� ��,��,%�0d  $RH�3!   �     � �}E���o�E�.l�Z���|,}�B��6�׸��_�I3��T0 k� ��)��)%�0d  $RH�3!   ��     � �}E�� �{�E�.��Y���|,}�B��7L۹��_�I3��T0 k� ��&��&%�0d  $RH�3!   ��     � �}E�� ���E�-��X���|,}�@�7Lߺ��_�I3��T0 k� ��$��$%�0d  $RH�3!   ��     � �}E��!���E�-��U���|,}�@�9L���_�I3��T0 k� ��#��#%�0d  $RH�3!   ��     � �}@-�!���E��-��T���|,}�@�:L���_�I3��T0 k� ��"��"%�0d  $RH�3!   ��     � �}@-�!���E��,��S���|,}�@�:L���_�I3��T0 k� ��"��"%�0d  $RH�3!   ��     � �}@-�"���E��,��Q���|,}�@�;L���_�I3��T0 k� ��"��"%�0d  $RH�3!   ��     � �}@-�"���E��,��P���|,}�@�;L���_�I3��T0 k� ��"��"%�0d  $RH�3!   ��     � �}@-�"���E��,��O���|,}�@�<L����_�I3��T0 k� ��#��#%�0d  $RH�3!   ��     � �}@-�#���D��,�M�� |,��@�=L�����_�I3��T0 k� ��#��#%�0d  $RH�3!   ��     � �}@-�#���D��,�L�|,��@�=L�����_�I3��T0 k� ��#� #%�0d  $RH�3!   ��     � �}@-�$���D��,�I�|,��@�?M����_�I3��T0 k� �$�$%�0d  $RH�3!   ��     � �}@-�$���D��,�G�|,��@�?M����_�I3��T0 k� �$�$%�0d  $RH�3!   ��     � �}E��$���D��,�F�|,��@�@M�-��_�I3��T0 k� ��*� *%�0d  $RH�3!   ��     � �}E��%���D��-�D�|,���@�@M�-��_�I3��T0 k� ��.��.%�0d  $RH�3!   ��     � �}E��%���L|�-�B�|,���@�AM�-��_�I3��T0 k� ��2��2%�0d  $RH�3!   ��     � �}E��&��L|�-�A�	|,���@�AM�-��_�I3��T0 k� ��4��4%�0d  $RH�3!   ��     � �}E��&��L|�-�?�
|,l��@ BM�-��_�I3��T0 k� ��6��6%�0d  $RH�3!   ��     � �}E��'��L|�-�?�|,l��@CM���_�I3��T0 k� ��8��8%�0d  $RH�3!   ��     � �}L}�(��L|�-��>�|,l��@DM���_�I3��T0 k� ��4��4%�0d  $RH�3!   ��     � �}L}�(�'�L|�,��>�|,l��@DM���_�I3��T0 k� ��1��1%�0d  $RH�3!   ��     � �}L}�)�+�L|�,��=�|,l��@EM#���_�I3��T0 k� ��/��/%�0d  $RH�3!   ��     � �}L}�)�3�L|�+��< |,l��@EM#���_�I3��T0 k� ��.��.%�0d  $RH�3!   ��     � �}L}�*�;�L|�+��<|,l��@FM'���_�I3��T0 k� ��-��-%�0d  $RH�3!   ��     � �}L}�*�?�L|�*��;|,l��@ FM+��_�I3��T0 k� ��-��-%�0d  $RH�3!   ��     � �}L}�+�G�L|�)��:|,���@$GM+��_�I3��T0 k� ��-��-%�0d  $RH�3!   ��     � �}L~ ,�K�L|�)��:|,���@(GM/��_�I3��T0 k� ��,� ,%�0d  $RH�3!   ��     � �}L~,�S�L|�(� 9|,���@,HM/��_�I3��T0 k� � ,�,%�0d  $RH�3!   ��     � �}L~-�[�L��(�9|,���@0HM3�� _�I3��T0 k� �,�,%�0d  $RH�3!   ��     � �}L~-�_�L��'�8|,���@4IM7��$_�I3��T0 k� �-�-%�0d  $RH�3!   ��     � �}L~.�g�L��'�8-|,���@8IM7��,_�I3��T0 k� �-�-%�0d  $RH�3!   ��     � �}L~.�k�L��'�8-|,���@<JM;��0_�I3��T0 k� �.�.%�0d  $RH�3!   ��     � �}L~/�o�L��&�7-|,���@@JM;��8_�I3��T0 k� �.�.%�0d  $RH�3!   ��     � �}L�/�w�L��&�7- |,���@@JM?��< _�I3��T0 k� �/� /%�0d  $RH�3!   ��     � �}L� /�{�L��&� 7-(|,���@DKMC��< _�I3��T0 k� � /�$/%�0d  $RH�3!   ��     � �}L�$0��L��&�(6-,!|,���@HKMC��@!_�I3��T0 k� �$0�(0%�0d  $RH�3!   ��     � �}L�(1��L��&�,6-0"|,���@LLMG��H"_�I3��T0 k� �(1�,1%�0d  $RH�3!   ��     � �}L�,2��L��%�06-4#|,���@PLMG��P$_|I3��T0 k� �(1�,1%�0d  $RH�3!   ��     � �}L�03��L��%�86-<$|,���@PLMK��T%_|I3��T0 k� �,2�02%�0d  $RH�3!   ��     � �}L�03��L��%�<6-@&|,���@TMMK��\&_xI3��T0 k� �03�43%�0d  $RH�3!   ��     � �}L�44��L��%�D6-@&|,���@XMMO��`'_xI3��T0 k� �44�84%�0d  $RH�3!   ��     � �}L�85��L��%�H7�H'|,���@\NMO��h)_tI3��T0 k� �84�<4%�0d  $RH�3!   ��    � �}L�85��L��$�P7�L'|,���@\NMS��l*_tI3��T0 k� �85�<5%�0d  $RH�3!   ��     � �}L�<6��L��$�T8�P(|,���@`NMS��t+_pI3��T0 k� �<6�@6%�0d  $RH�3!   ��     � �}L�@7��L��$�\9�X)|,���@dOMW��x,_pI3��T0 k� �@6�D6%�0d  $RH�3!   ��     � �}L�D7��L��$�`:�\*|,���@hOMW���-_pI3��T0 k� �@7�D7%�0d  $RH�3!   ��     � �}L�D8��L��$�h:�d*|,���@hOMW���/_lI3��T0 k� �D8�H8%�0d  $RH�3!   ��     � �}L�H9��L��#�l;�h+|,���@lPM[���0_lI3��T0 k� �H8�L8%�0d  $RH�3!   ��     � �}L�L9���L��#t<�p,|,���@pPM[���1_hI3��T0 k� �H9�L9%�0d  $RH�3!   ��     � �}L�L:���L��#x=�t-|,���@pPM_���2_hI3��T0 k� �L:�P:%�0d  $RH�3!   ��     � �}L�P;���L��#�>�|.|,���@tQM_���3_hI3��T0 k� �P:�T:%�0d  $RH�3!   ��     � �}L�T;���L��#�?��/|,���@xQMc���4_dI3��T0 k� �P;�T;%�0d  $RH�3!   ��    � �}L�T<���L��#�@��0|,���@xQMc���5_dI3��T0 k� �T<�X<%�0d  $RH�3!   ��     � �}L�X<���L��#�A�1|,���@|RMc���6_dI3��T0 k� �X<�\<%�0d  $RH�3!   ��     � �}L�X=���L��"�B�2|,���@�RMg���7_`I3��T0 k� �X=�\=%�0d  $RH�3!   ��     � �}L�\>���L��"	=�C�3|,���@�RMg���8_`I3��T0 k� �\=�`=%�0d  $RH�3!   ��     � �}L�`>���L��"	=�D�4!�,���@�SMk���9_`I3��T0 k� �\>�`>%�0d  $RH�3!   ��     � �}L�`?���L��"	=�E�5!�,���@�SMk���:_\I3��T0 k� �`?�d?%�0d  $RH�3!   ��     � �}L�d?���L��"	=�E��5!�,���@�SMk���;_\I3��T0 k� �d?�h?%�0d  $RH�3!   ��     � �}L�d@���L��"	=�F��6!�,���@�TMo���<_\I3��T0 k� �d@�h@%�0d  $RH�3!   ��     � �}L�h@���L��!	=�G��7!�,���@�TMo���=_XI3��T0 k� �h@�l@%�0d  $RH�3!   ��     � �}L�hA���L��!	M�H��8!�,���@�TMs� n�>_XI3��T0 k� �hA�lA%�0d  $RH�3!   ��     � �}L�lA���L��!	M�I��8!�,���@�TMs� n�?_XI3��T0 k� �lA�pA%�0d  $RH�3!   ��     � �}L�lB�� L��!	M�J��9!�,���@�UMs� n�@_TI3��T0 k� �lB�pB%�0d  $RH�3!   ��     � �}L�pB��L��!	M�K��:!�,���@�UMw� n�A_TI3��T0 k� �pB�tB%�0d  $RH�3!   ��     � �}L�pC� L��!	M�K��;!�,���@�UMw� n�B_TI3��T0 k� �pC�tC%�0d  $RH�3!   ��     � �}L�tC�L��!	=�L��<!�,���@�UMw� n�B_PI3��T0 k� �tC�xC%�0d  $RH�3!   ��     � �}L�tD�L��!	=�M��<|,���@�VM{� n�C_PI3��T0 k� �tD�xD%�0d  $RH�3!   ��     � �}L�xD�L�� 	=�N��=|,���@�VM{� n�D_PI3��T0 k� �xD�|D%�0d  $RH�3!   ��     � �}                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��MT ]�)�)� p �� Y^
  $ $     ���yR     Yu�����    ���             /  Z�}          ��     ���  0	%           W��   � �  	   �����     Wۚ���a    ���q                Z�}          	��  (  ���   0	           P�  � �
     �t�     Q��tJ�    �>�j             ;	 Z�}           ��    ���  8	           a¼   � �
	   �qM     aק�qMB    ���[                	 Z�}         ���    ���   8          i�)   � �	    .��#�     i���X�    �=�z              (	 Z�}          ��    ���   P
	
          ��  ��	      B��     ����                             ���z              8  ���    P             ��=C        V�+�     ��=C�+�                          �         �     ��B   H	$
          sc�          j���     sXH����     � n              � �          �      ��@   8�           ��=  $ $       ~�sh�    ��c�sc     : U                 C �         �@     ��@   (
          u�)         ����4     u�x����     � n            
     �        	 ��     ��J   0
9          Gtu         ��ݘE     Gtu�ݔ�       2                 A �         
 ��     ��@   H

!         ��� ��     � ���    ��� ���                           ���4              x  ��@                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          d�  ��        ����#     d�N��WM    ��� "              x                j  �        �                          d    ��        ���       d  ��           "                                                �                         �����t�q����+���s���� �������  
               	
  *   RK ��G       �$ ``� �� @a� �d  b  �� f� � 0f� Ф d� &� _ ���< ����J ����X ���� ���� ����  ����. ����< ����J ����X � 
�� V� 
�\ W  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �� �R� � }`���� � 
� W� 
�� W� 
�\ W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����}�� �� �  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    "�j�� , " �
� �  �  
�  Y    ��     ���       Y    ��     ���       u    ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  � %%9      �� � �  ���        �#T ���        �        ��        �        ��        �     ��      �� 1�        ��                         ��  0  ����                                    �                ����             Y�� ���%��   �} 2               85 Petr Klima   sh     0:01                                                                        2  1     �_� �_� �FCB �O CJ �HCK	+cV �C c^ � �CQ � 	C"Y � 
C#I � C$I � C%T � C&O �c~ � � c� � �	K= �KC �KC �C._ �C1` �C3X � C6g �C7V �J�L � J�\ � �[ � �Z �B�E � B�M �kjd c�h � c�x {!c�9 � "c�A �#"�G � $"�Y �%�C �&
�R �'"�G � ("�Y �)"�C �**�R �+"�c � ,"�u �-�_ � 
�n � 
�n � 
�n �1�S � 
�b � 
�` �4�2 � 
�A � 
�8 � 
�* � 8"P � 9"& y.  "* y � ;"P �" <"& z2  "* z:  "J �>  *Go                                                                                                                                                                                                                         �� R         �     @ 
        �     S P E e  ��         	           	 �������������������������������������� ���������	�
��������                                                                                          ��    ��:�� ��������������������������������������������������������   �4, 8� ���@��@��A�����                                                                                                                                                                                                                                                                                                                                            7 ��	@m��5��j�x�                                                                                                                                                                                                                             ]  	  (        D�J    	  �                             ������������������������������������������������������                                                                                                                                          �      �      �                � �          	  
 	 
 	 	 ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ���            .                     
  #    ��  H�J     .�                             �������������������������������������������������������                                                                                                                                      :L 7    �      [        �    B I D   }      
 	  
	 
 	 	 ���������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������            r                                                                                                                                                                                                                                         
                                                                       �             


            ��  }�                       N�           +                                                    ����    ������������   '������������   ����������������    ��������   	����������������  's������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" A C 6               	                  � �Y� �\        |3b�T�q�$Hb2�                                                                                                                                                                                                                                                                   )n)n1n  )�                            d      a            d      m                                                                                                                                                                                                                                                                                                                                                                                                                > �  >�  J�  2�  C#�  EZm�  �N /��f���� Y�˖�����������������������c�                      ��       	 	 �   & AG� �  j   
              �                                                                                                                                                                                                                                                                                                                                        B C   �                        !��                                                                                                                                                                                                                            Y��   �� � ���      �� B 	     ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ������������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    3      +      d                       B         �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$    `d  �@���6 ��  �@���6 �$ ^$ �s@  �@  �s@      p 
�� 	��   ����@ ��   � � �$ ^$      �  ��              � ��� ��  �  � ��� �� � ��� �$ c �  ��c  �      �  ��   \�����������J   g��� 	       f ^�         �� �       \      ��M��������J���J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         7v` weV "fff"O�p"��p"��p"�p3�}p-��p=��p|� }�  }�  ��  ��  ��  ��  �  �  �  �  �  "              `  eV  fff O�  ��  ��  �  �} �� �� ��  |�  }�  ��    =   }   =   =              �������}�}�}�ww~r�� ∈�������������������}�� }�� ��� ��� ����   �   �   �   �   �   �   �   C""42""#2""#2""#2""#s3342"""3333    p   p   p   p   p   p   p    ��������� ��� }�� ��  ��  ����  ��  ��  ��  ��  ��  ��  ��                          � �� ��    "               wvf wfU 7Of`w��f"�� "�p-�}p���� ��� ����x��	�� �� �� "�        f  U` f` f` �p w���� `  eV  ff  O�  ��  �� ����}�                �  �  ��  �            �  �  �   �  ��  �                     �  �  �   � `  eV  ff  O�  ��  ��  ����}���������������p	���         `  eV  ff  O�  ��  ��  ���}�     �  �  �   �  ��  �   �            ��  ��  �   ��  �   ���������������p	���                    3333UUUU                        wwww                    333333333333333333333   w  G� ws@ ws� ws$7w@wwww"                               ����������� ��� �� ��  �    `  eV  ff  O�  ��  ��  � ��}�            """"                  w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "" "  """""" "!   " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """""" "!   " ""  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  " ! " ""  "!  "! " ""            """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                             �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �          
 "� ""� ""� "                       �                             ���                         �  ��                    �����                                        � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                           �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw     �  �  ��  �   �   �         ��                                 � ���� ��   � � �         � � ��      �                                                                                                                                "  "(��ȩ�ܚ��ۊ����� ��  �   �   �   �   �� ��� ̻� ˽� ��� �w� �������������������������� �̻ ���         �   �       �   �   "" �+� Ȼ� ɫ� ɨ� ��                �� �I��3 ��D 
UD 
UD TD  T�  ˸  ��  �� ̰ �+ ��"/ �"/  ����  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �   �   �                .      �����                      �  �  �   �   ��  �                            �   ���                            �   �                                                                                                         �  �  �  �� ݚ� }�Ȫ��˙������˼� ��  ��  ��  ��  ��  I� H� �E X�T X�S T�D �[ ˻  ˸  ��  
� �,"��"" "  �" �  ""� �� ˻ �˻ ��ݪ��کɨ��ˀ�̽ ��� ��  ̽  ̻  ̻  ˉ  ��  �D  DC  C3  #;  ;�� �� ��  �� "�  "  �"/ / ����� ��  �      �   �          �  �  "     "  "  "   "�  �  �   �   
                            �          �   �          �                    ��  ���� ��    �����                                       ���                                                                                                                                                                           ۻ� ۽� ��� H�DH�D�DP�E X�T H�P H�@ Ȥ� ̻� ˘ �� "*� �/�""/""/���                       ��  ۼ� ݻ� w�� b}ذgvz�w������ɨ�ͨ���ڋ��٭���ۻݻ� �   �          �   �   .   ."  ""  ""  ,   �   
            "  "  ""  "�   �           �   ��  �      �                                     �  �  �  ��  �  �  �  ��  �             �   �   �             � � "            � "�",�"+� ",                       "  .���"    �     �                                                                                                                                                                                          �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                    �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��     �   �  �  �  �  �   �                    �� �� �� w� m| ��  �  ��  ��  �   �                     "  ""  """"""
�                               	�    �     �                                                                                                                                                                                     �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �    �   ��  �  ��  �             �  �   �   ��  �            ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    � �� �  �  �      �   �     ���                                                                                                                                                                                                  �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   �   �"  ""  !� �� ��  �               �   ������  ��                      �   �                      �������  ���    �        �  ��  �                            �  �˰ ��� �wp ���      � �������������  �                                                                                                                                                              	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                                   ��                  �                        ���� ��� ����                �  ��  �                            �  �˰ ��� �wp ���                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  ��  ��  �                       �,� �"/�""�"/� "/  �         "  "  ""  "+� �� � ��   �  "   "�  +�  
�� ��� D�D 4ETO3    �   �   �   D   E�  U�  UO                         "  "  "      � �������������  �                                                                                                                                                                �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                �  ��  �               �                                                                                                                                                                                    �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(����������������� � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(����������������� 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5���������������� x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x���������������� w w x y�������H���������������������������������H������yxww����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq_� �_� �FCB �O CJ �HCK	+cV �C c^ � �CQ � 	C"Y � 
C#I � C$I � C%T � C&O �c~ � � c� � �	K> �KD �KD �C._ �C1` �C3X � C6g �C7V �J�L � J�\ � �[ � �Z �B�E � B�M �kjd c�h � c�x {!c�9 � "c�A �#"�G � $"�Y �%�C �&
�R �'"�G � ("�Y �)"�C �**�R �+"�c � ,"�u �-�_ � 
�n � 
�n � 
�n �1�S � 
�b � 
�` �4�2 � 
�A � 
�8 � 
�* � 8"P � 9"& y.  "* y � ;"P �" <"& z2  "* z:  "J �>  *Go3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������;�U�T��=�[�M�T�[�Z�Z� � � � � � � � � �/�.�7�����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.����������������������������������������#� ��9�K�Z�X��5�R�O�S�G� � � � � � � � � � �/�.�7�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������/�.�7� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 