GST@�                                                            \     �                                               � ���      �              ����e $�	 J�������������������        �g      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"��   " `  J  jF��    "�j "����
��
��     �j�� 
   ��
  �                                                                               ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������oo    og     +      '            ��                     	  7  V  	                  �            :8 �����������������������������������������������������������������������������                                ��  �       |�   @  #   �   �                                                                                '       )n)n1n  �    H   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��E�O�C�o���E��ZlC�C�Ӯ������қ��#�3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� J��E�G�C�k����E��ZlC�C�ˮ������җ��#�3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� G��E�C�C�c���E���ZlC�C�������җ���3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� D��E�3�C�c�� E��ZlC�C������җ���3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� @��E�+�C�[�� Er�ZlC�EQ�������җ���3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� <��E�#�C�S��Er�ZlC�EQ�������җ���3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� 9��E��C�K�?�Er�ZlC�EQ�������җ���3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� 6��I��C�G�?�Er�ZlC�EQ������җ���3��T0 k� ������&�1D"3Q2	4#'Q  �'    ��� 0��I��C�?�?�Er�ZlC�EQ���������3��T0 k� �{���&�1D"3Q2	4#'Q  ��/    ��� *��I���C�7�?�Er#�ZlC�EQw�!��������3��T0 k� �o��s�&�1D"3Q2	4#'Q  ��/    ��� $��I���C�/�?�Er'�ZlC�EQk�!��������3��T0 k� �c��g�&�1D"3Q2	4#'Q  ��/    ��� ��I���C����Er3�ZlC�EQ[�!��������3��T0 k� �K��O�&�1D"3Q2	4#'Q  ��/    ��� ��I���C����Er7�ZlC�EQS�!���������3��T0 k� �?��C�&�1D"3Q2	4#'Q  ��/    ��� ��I���C����Er;�ZlC�EQG�1��{������3��T0 k� �3��7�&�1D"3Q2	4#'Q  ��/    ��� ��I���C����Eb?�ZlC�EQ?�1��s�������3��T0 k� �'��+�&�1D"3Q2	4#'Q  ��/    ��� ��I���C����	EbG�ZlC�C�7�1{�k�������3��T0 k� ���#�&�1D"3Q2	4#'Q  ��/    ��� ��I���C���|	EbK�ZlC�C�+�1s�c�������3��T0 k� ����&�1D"3Q2	4#'Q  ��&    ��� ��I���C���x
EbO�ZlC�C�#�1o�[�������3��T0 k� �����&�1D"3Q2	4#'Q  ��&    ��� ��I���C����pEbS�ZlC�C��Ag�W�������3��T0 k� ����&�1D"3Q2	4#'Q  ��&    �������I���C���hEbS�ZlC�C��A_�O�������3��T0 k� �۱�߱&�1D"3Q2	4#'Q  ��&    �������I���C���`EbW�ZlC�EQ�A[�G�������3��T0 k� �ׯ�ۯ&�1D"3Q2	4#'Q  ��&    �������I���C���XEb[�ZlC�EP��AS�?�	�����3��T0 k� �ӭ�׭&�1D"3Q2	4#'Q  ��&    �������Ea��C���PEb_�ZlC�EP��AO�3�	�����3��T0 k� �ˬ�Ϭ&�1D"3Q2	4#'Q  ��&    �������Ea��C���HEb_�ZlC�EP�AG�+�	�����3��T0 k� �ǫ�˫&�1D"3Q2	4#'Q  ��&    �������Ea��C���@Ebc�ZlC�EP�AC�#�	�����3��T0 k� ����ê&�1D"3Q2	4#'Q  ��&    �������Ea��C���8ERc�ZlC�EP۳A;��	�����3��T0 k� ������&�1D"3Q2	4#'Q  ��&    �������Ea��C���0ERg�ZlC�EPϳA7��	�����3��T0 k� ������&�1D"3Q2	4#'Q  ��&    �������Ea��C���(ERg�ZlC�A`ǳA/��
�����3��T0 k� ������&�1D"3Q2	4#'Q  ��&    �������EQ{�E��� ERk�ZlC�A`��A+��
�����3��T0 k� ������&�1D"3Q2	4#'Q  ��&    �������EQs�E���ERk�ZlC�A`��A#���
��B��3��T0 k� �w��{�&�1D"3Q2	4#'Q  ��&    �������EQk�Eѻ�ERk�ZlC�A`��A���
��B��3��T0 k� �g��k�&�1D"3Q2	4#'Q  ��&    �������EQc�Eѷ�ERk�ZlC�A`��A���
��B��3��T0 k� �W��[�&�1D"3Q2	4#'Q  ��&    �������EQ[�Eѯ�C�k�ZlC�EЗ�A���	��B��3��T0 k� �W��[�&�1D"3Q2	4#'Q  ��&    �������EQS�Eѫ��C�k�ZlC�EЏ�A���	��B��3��T0 k� �W��[�&�1D"3Q2	4#'Q  ��&    �������EQS�Eѣ��C�k�ZlC�EЇ�A����	�� ��3��T0 k� �S��W�&�1D"3Q2	4#'Q  ��&    �������EQO�EA���C�k�ZlC�E�{�A����	�� ��3��T0 k� �O��S�&�1D"3Q2	4#'Q  ��&    �������EQG�EA���C�k�ZlC�E�s�@����	�� ��3��T0 k� �K��O�&�1D"3Q2	4#'Q  ��&    �������EQ?�EA���C�k�ZlC�E�k�@����
�� ��3��T0 k� �C��G�&�1D"3Q2	4#'Q  ��&    �������EA;�EA����C�k�ZlC�E�c�@����
�� ��3��T0 k� �?��C�&�1D"3Q2	4#'Q  ��&    �������EA3�EA����C�g�ZlC�E�W�@����
�� ��3��T0 k� �7��;�&�1D"3Q2	4#'Q  ��&    �������EA+�EA���C�g�ZlC�E�O�P����
�� ��3��T0 k� �+��/�&�1D"3Q2	4#'Q  ��&    �������EA#�EAw���C�c�ZlC�E�G�P����
�� ��3��T0 k� �#��'�&�1D"3Q2	4#'Q  ��&    �������EA�EAo���C�c�ZlC�E�;�P����	� ��3��T0 k� ����&�1D"3Q2	4#'Q  ��&    �������EA�EAk���C�_�ZlC�A�3�P����	� ��3��T0 k� ����&�1D"3Q2	4#'Q  ��&    �������EA�C�_���C�_�ZlC�A�+�P���w�	�ø ��3��T0 k� �����&�1D"3Q2	4#'Q  ��&    �������EA�C�S���C�[�ZlC�A��P���o�	�÷ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��&    �������EA�C�G���C�[�ZlC�A��P���g�	�ö ��3��T0 k� ������&�1D"3Q2	4#'Q  ��&    �������EA�C�?�~�C�W�ZlC�A��P���_�
õ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��&    �������C���C�3�~�C�S�Z�C�A��P���W�
Ǵ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��&    �������C���C�'�~�C�O�Z�C�A���P���O�
ǳ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��&    �������C���C��~�C�K�Z�C�A��P���C�
ǲ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��&    �������C���C��~�C�G�Z�C�A��@���;�
Ǳ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    �������C���C��~�C�C�Z�C�E_ߺ@���3�	�ǰ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    �������C���C���~�C�?�Z�C�E_׺@���+�	�˰ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    �������E���C���~�C�;�Z�C�E_ϻ@��#�	�˯ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    �������E���C��~�D7�Z�C�E_ǻ@w���	�ˮ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    �������Eп�C��~�D3�Z�C�E_��@o���	�˭ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    �������Eз�C�ۺn�D/�Z�C�E_��@k��
Ϭ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    �������EЯ�C�Ӹn�D+�Y|C�E_��@c� ��
Ϭ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    �������EЧ�C�Ƿn�D#�Y|C�E_��@[� ��
ϫ ��3��T0 k� �����&�1D"3Q2	4#'Q  ��6    �������EЛ�C���n�D�Y|C�E_��@S� ��
Ϫ ��3��T0 k� �w��{�&�1D"3Q2	4#'Q  ��6    �������EГ�C���n�D�Y|C�E@K� ��
ϩ ��3��T0 k� �o��s�&�1D"3Q2	4#'Q  ��6    �������EГ�C�����D�Y|C�E0C����	�ө ��3��T0 k� �c��g�&�1D"3Q2	4#'Q  ��6    �������EЋ�C�����D�Y|C�E��0;����	�Ө ��3��T0 k� �[��_�&�1D"3Q2	4#'Q  ��6    �������C���C�����D�Y|C�E�s�03����	�ӧ ��3��T0 k� �S��W�&�1D"3Q2	4#'Q  ��6    �������C�{�C�����D�Y|C�E�k�0+����	�Ӧ ��3��T0 k� �K��O�&�1D"3Q2	4#'Q  ��6    ������ C�s�C�����D��Y|C�E�c�0#���	�Ӧ ��3��T0 k� �?��C�&�1D"3Q2	4#'Q  ��6    ������ C�k�C�����D��Y|C�E�W�0���
ӥ ��3��T0 k� �7��;�&�1D"3Q2	4#'Q  ��6    ������ C�c�C����D��Y|C�E�O�0���
פ ��3��T0 k� �/��3�&�1D"3Q2	4#'Q  ��6    ������ C�[�C�w�~�D��Y|C�E�G�0���
פ ��3��T0 k� �#��'�&�1D"3Q2	4#'Q  ��6    ������ C�S�E�o�~�D��Y|C�E�?�@����
ף ��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ������ C�G�E�g�~|D��Y|C�E�7�O�����
ף ��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ����~� C�?�E�_�~xD��Y|C�E�+�O��0��	�ע ��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ����|� C�7�E�W�~xD��Y|C�E�#�O��0�	�ס ��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ����z� C�/�E�O�~tD��Y|C�E��O��0w�	�ۡ ��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ����x� C�'�E�G�~tD��Y|C�E��O��0o�	�۠ ��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ����v� C��E�?�npD��Y|C�E��O��0g�	�۠ ��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ����t� C��E�7�nlC��Y|C�E��O��0_�
۟ ��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ����r� C��E�+�nlC��Y|C�E���O��0W�
۞ ��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ����p� C��E�#�nhC��Y|C�E���O��0O�
۞ ��3��T0 k� �����&�1D"3Q2	4#'Q  ��6    ����n� C���E��ndC��Y|C�E���O��0C�
ߝ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����l� E���E��>`C��Y|C�E���O��0;�
ߝ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����j� E���E��>\
C��Y|C�E���_��03�	�ߜ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����h� E���E���>\C��Y|C�E���_��0+�	�ߜ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����f� E���E���>XC�{�Y|C�F��_��@#�	�ߛ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����d� E���E��>TC�s�Y|C�F��_��@�	�ߛ ��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� E���E���PC�o�Y|C�F��_��@�	�ߚ ��3��T0 k� ������&�1D"3Q2	4#'Q  �6    ����c� E���E�ۘ�LAQg�Y|C�F��ϛ�@�r� b��3��T0 k� ������&�1D"3Q2	4#'Q  �6    ����c� A_��E�Ә�HAQ_�Y|C�F��ϗ�@�r� b��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_��E�˗�HAQW�Y|C�F��Ϗ�O��r� b��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_��A�Ö�G�AQO�Y|C�F��ϋ�O��r� b��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_��A����C�AQG�Y|C�B^��σ�O��r� b��3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_��A����?�AQC�Y|C�B^����O��r� ���3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_��A����;�AQ;�Y|C�B^���w�O��b� ���3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_��A����;�AQ3�Y|C�B^���s�O��b� ���3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_��A����7�AQ/�Y|C�B^���k�_��b� ���3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_{�A����3�AQ'�Y|C�B^���g�_��b� ���3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_s�A���/�AQ�Y|C�B^���_�_��b���3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_k�A���/�AQ�Y|C�E~���[�_��b���3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_g�A�{�+�AQ�Y|C�E~���S�_��b���3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A__�A�s�+�AQ�Y|C�E~��K�_��R���3��T0 k� ������&�1D"3Q2	4#'Q  ��6    ����c� A_W�A�k�'�AQ�a�C�E~{��G�_��Rߎ��3��T0 k� �� �� &�1D"3Q2	4#'Q  ��6    ����c� A_O�A�c��+�AQ�a�C�E~w��?�_��Rߎ��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ����c� A_K�A�_��/�AP��a�C�E~s��7�_��RߍR��3��T0 k� ����&�1D"3Q2	4#'Q  ��6    ����cC� A_C�A�W��/�AP��a�C�E~o��3�_��RیR��3��T0 k� �|��&�1D"3Q2	4#'Q  ��6    ����cC� A_?�A�O��3�AP��a�C�E~o��+�_{�RۋR��3��T0 k� �x	�|	&�1D"3Q2	4#'Q  ��6    ����cC� A_7�A�G��3�AP��a�C�E~k��#�os�R׊R��3��T0 k� �t�x&�1D"3Q2	4#'Q  ��6    ����cC� A_/�A�C��7�AP��a�C�E~g���ok��׉R��3��T0 k� �t�x&�1D"3Q2	4#'Q  ��6    ����cC� A_+�A�;��;�AP��a�C�E~c���oc��ӈ���3��T0 k� �p�t&�1D"3Q2	4#'Q  ��6    ����cC� A_#�A�7��;�AP��a�C�En_�� o[��ӈ���3��T0 k� �\�`&�1D"3Q2	4#'Q  ��6    ����cC� A_�A�/��?�AP��a�C�En_��oS��χ���3��T0 k� �L�P&�1D"3Q2	4#'Q  ��6    ����cC� A_�A�+��?�AP��a�C�EnX ��oK��ˆ���3��T0 k� �@�D&�1D"3Q2	4#'Q  ��6    ����cC� A_�A�#��C�AP��Y|C�EnT��?C��˅���3��T0 k� �4�8&�1D"3Q2	4#'Q  ��6    ����c� A_�A���G�AP��Y|C�EnP��?;��ǅ���3��T0 k� �,�0&�1D"3Q2	4#'Q  ��6    ����c� A_�A���G�AP��Y|C�EnL��?3��Ä���3��T0 k� �(�,&�1D"3Q2	4#'Q  ��6    ����c� A_�A���K�AP��Y|C�EnH	��?/�⿃���3��T0 k� � �$&�1D"3Q2	4#'Q  ��6    ����c� A^��A���K�AP��Y|C�EnD��?'�⻂���3��T0 k� ��&�1D"3Q2	4#'Q  ��6    ����c� A^��A���O�AP��Y|C�En@>�?�ⷂ���3��T0 k� ��&�1D"3Q2	4#'Q  ��6    ����c� A^�A����O�AP��Y|C�En<>�?�ⳁ���3��T0 k� ��&�1D"3Q2	4#'Q  ��6    ����c� A^�A����S�AP��Y|C�M>8>�?�����3��T0 k� � � &�1D"3Q2	4#'Q  ��6    ����c� A^�A����S�AP��Y|C�M>4>�	?�����3��T0 k� �#�#&�1D"3Q2	4#'Q  ��6    ����c� A^�A���W�AP��Y|C�M>0>�	?�����3��T0 k� �%�%&�1D"3Q2	4#'Q  ��6    ����c� A^߼A���W�AP��Y|C�M>,>�
>������3��T0 k� �'�'&�1D"3Q2	4#'Q  ��6    ����c� A^ۼA���[�AP��a�C�M>(�
>������3��T0 k� �)�)&�1D"3Q2	4#'Q  ��6    ����c� A^׼A���[�AP��a�C�M>$�>������3��T0 k� �*�*&�1D"3Q2	4#'Q  ��6    ����c� A^ϼA�ۆ�_�AP��a�C�M> �>������3��T0 k� �,�,&�1D"3Q2	4#'Q  ��6    ����c� A^˼A�ׅ�_�AP��a�C�M> �N������3��T0 k� �.�.&�1D"3Q2	4#'Q  ��6    ����c� A^ǻA�Ӆ�c�AP��a�C�M> �N�����3��T0 k� �0�0&�1D"3Q2	4#'Q  ��6    ����c� A^ûA�υNc�AP��a�C�M>"�|N�����3��T0 k� �2�2&�1D"3Q2	4#'Q  ��6    ����c� A^��A�˄Nc�AP�a�C�MN$�tN�����3��T0 k� �3�3&�1D"3Q2	4#'Q  ��6    ����c� A^��A�ÄNg�AP�a�C�MN&�lN��w���3��T0 k� � 5�5&�1D"3Q2	4#'Q  ��6    ����c� A^��A���Ng�AP{�a�C�MN'�dN��s���3��T0 k� ��6� 6&�1D"3Q2	4#'Q  ��6    ����c� A^��A���Nk�APw�a�C�MN)�\N��o���3��T0 k� ��8��8&�1D"3Q2	4#'Q  ��6    ����c� A^��A���Nk�APs�a�C�MN+�TN��k���3��T0 k� ��:��:&�1D"3Q2	4#'Q  ��6    ����c� A^��A���No�APo�Y|C�MN,�LN��c���3��T0 k� ��;��;&�1D"3Q2	4#'Q  ��6    ����c� A^��A���No�APk�Y|C�MN .�DN��_���3��T0 k� ��=��=&�1D"3Q2	4#'Q  ��6    ����c� A^��A���No�APg�Y|C�MN 0�<N��[���3��T0 k� ��?��?&�1D"3Q2	4#'Q  ��6    ����c� A^��A���Ns�APc�Y|C�MM�1�4N��W���3��T0 k� ��@��@&�1D"3Q2	4#'Q  ��6    ����c� A^��A���Ns�AP_�Y|C�M=�3�0N��S���3��T0 k� ��B��B&�1D"3Q2	4#'Q  ��6    ����c� A^��A���Ns�AP_�Y|C�M=�4�(N��K���3��T0 k� ��C��C&�1D"3Q2	4#'Q  ��6    ����c� A^��A���Nw�AP[�Y|C�M=�6� 
N��G��3��T0 k� ��E��E&�1D"3Q2	4#'Q  ��6    ����c� A^��A���Nw�APW�Y|C�M=�7�
N��C�{�3��T0 k� ��F��F&�1D"3Q2	4#'Q  ��6    ����c� A^��A���N{�APS�Y|C�M=�9�	N��?�s�3��T0 k� ��H��H&�1D"3Q2	4#'Q  ��6   ����c� A^��A���N{�APO�Y|C�M=�:�	N��";�o�3��T0 k� ��I��I&�1D"3Q2	4#'Q  ��6    ����c� A^��A���N{�APO�Y|C�M=�<�N��"7�g�3��T0 k� ��K��K&�1D"3Q2	4#'Q  ��6    ����c� A^��A���N�APK�Y|C�M=�=� N��"3�_�3��T0 k� ��L��L&�1D"3Q2	4#'Q  ��6    ����c� A^�A���N�APG�Y|C�M=�>��N�"/�[�3��T0 k� ��M��M&�1D"3Q2	4#'Q  ��6    ����c� A^{�A���N�APC�Y|C�A��@��N{�"+�S�3��T0 k� ��M��M&�1D"3Q2	4#'Q  ��6    ����c� A^w�A���N��APC�Y|C�A��A��Nw�"'�K�3��T0 k� ��L��L&�1D"3Q2	4#'Q  ��6    ����c� A^s�A��N��AP?�Y|C�A��B��Ns�"#��G�3��T0 k� ��L��L&�1D"3Q2	4#'Q  ��6    ����c� A^o�A�{�N��AP;�Y|C�A��C��No�"��?�3��T0 k� ��M��M&�1D"3Q2	4#'Q  ��6    ����c� A^o�A�w�N��AP;�Y|C�A��E��Nk�"��7�3��T0 k� ��M��M&�1D"3Q2	4#'Q  ��6   ����c� A^k�A�s�N��AP7�Y|C�A��F��Ng�"��/�3��T0 k� ��N��N&�1D"3Q2	4#'Q  ��6    ����c� A^g�A�s�N��AP3�Y|C�A��G��Nc�"��'�3��T0 k� ��O��O&�1D"3Q2	4#'Q  ��6   ����c� A^c�A�o�N��AP3�Y|C�A��H�� N_�"��#�3��T0 k� ��P��P&�1D"3Q2	4#'Q  ��6    ����c� A^c�A�k�N��AP/�Y|C�A��J���N_�"���3��T0 k� ��Q��Q&�1D"3Q2	4#'Q  ��6   ����c� A^_�A�g�N��AP+�Y|C�A��K���N[�"���"s��T0 k� ��R��R&�1D"3Q2	4#'Q  ��6    ����c� A^[�A�c�N��AP+�Y|C�M=�L���NW�"���"s��T0 k� ��U��U&�1D"3Q2	4#'Q  ��6    ����c� A^[�A�_�N��AP'�Y|C�M=�M���NS�"���"s��T0 k� ��X��X&�1D"3Q2	4#'Q  ��6    ����c� A^W�A�_�N��AP'�Y|C�M=�N���NO�!�����"s��T0 k� ��Z��Z&�1D"3Q2	4#'Q  ��6    ����c� A^S�A�[�N��AP#�Y|C�M=�O���NK�!�����"s��T0 k� ��]��]&�1D"3Q2	4#'Q  ��6    ����c� A^S�A�W�N��AP�Y|C�M=�P���NG�!�����"s��T0 k� ��_��_&�1D"3Q2	4#'Q  ��6    ����c� A^O�A�S�N��AP�Y|C�M=�Q���NC�!����"s��T0 k� ��`��`&�1D"3Q2	4#'Q  ��6    ����c� A^K�A�S�N��AP�Y|C�M=�R���NC�!����"s��T0 k� ��a��a&�1D"3Q2	4#'Q  ��6    ����c� A^K�A�O�N��AP�Y|C�M=�S���N?�!����"s��T0 k� ��b��b&�1D"3Q2	4#'Q  ��6    ����c� A^G�A�K�N��AP�Y|C�M=�T���N;�!����"s��T0 k� ��c��c&�1D"3Q2	4#'Q  ��6    ����c� A^C�A�G�N��AP�Y|C�M=�U���N7�!���"s��T0 k� ��d��d&�1D"3Q2	4#'Q  ��6    ����c� A^C�A�G�N��AP�Y|C�MM�V���>3�!���3��T0 k� ��e��e&�1D"3Q2	4#'Q  ��6    ����c� A^?�A�C�N��AP�Y|C�MM�W���>3�!���3��T0 k� ��f��f&�1D"3Q2	4#'Q  ��6    ����c� A^?�A�?�N��AP�Y|C�MM�X���>/�!߉��3��T0 k� ��g��g&�1D"3Q2	4#'Q  ��6    ����c� A^;�A�?�N��AP�Y|C�MM�Y��>+�!߉��3��T0 k� ��h��h&�1D"3Q2	4#'Q  ��6    ����c� A^7�A�;�N��AP�Y|C�MM�Z�{�>'�!ۊ��3��T0 k� ��i��i&�1D"3Q2	4#'Q  ��6    ����c� A^7�A�7�N��AP�Y|C�MM�[�w�>'�!׊��3��T0 k� ��j��j&�1D"3Q2	4#'Q  ��6    ����c� A^3�A�7�N��AP�Y|C�MM�\�s�>#�!ӊ��3��T0 k� ��k��k&�1D"3Q2	4#'Q  ��6    ����c� A^3�A�3�N��AP�Y|C�MM�]�o�>�!ӊ{�3��T0 k� ��k��k&�1D"3Q2	4#'Q  ��6    ����c� A^/�A�/�N��AP�Y|C�MM�^�k�>�!ϊs�3��T0 k� ��l��l&�1D"3Q2	4#'Q  ��6    ����c� A^/�A�/�N��AP�Y|C�M=�_�g�>�!ϊk�3��T0 k� ��n��n&�1D"3Q2	4#'Q  ��6    ����c� A^+�A�+�N��A_��Y|C�M=�_�c�>�!ˊc�3��T0 k� ��o��o&�1D"3Q2	4#'Q  ��6   ����c� A^+�A�+�N��A_��Y|C�M=�`�_�>�!Ǌ[�"���T0 k� ��p��p&�1D"3Q2	4#'Q  ��6    ����c� A^'�A�'�N��A_��Y|C�M=�a�[�>�!ǊS�"���T0 k� ��q��q&�1D"3Q2	4#'Q  ��6    ����c� A^'�A�#�N��A_��Y|C�M=�b�W�>�!ËG�"���T0 k� ��q��q&�1D"3Q2	4#'Q  ��6    ����c� A^#�A�#�N��A_��Y|C�M=�c�S�>�!Ë?�"���T0 k� ��r��r&�1D"3Q2	4#'Q  ��6    ����c� A^#�A��N��A_��Y|C�M=�c�O�>�!��7�"���T0 k� ��s��s&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�M=�d]K�=��!��/�"���T0 k� ��t��t&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�M=�e]G�=����'�"���T0 k� ��u��u&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��f]C�M����#�"���T0 k� ��s��s&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��f]?�M����"���T0 k� ��r��r&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��g]?�M����"���T0 k� ��r��r&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��h];�M����"���T0 k� �|r��r&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��h]7�M����3��T0 k� �|q��q&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��i]3�M�ᯋ��3��T0 k� �|q��q&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��j]/�M۸ᫌ��3��T0 k� �xr�|r&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��k]/�M׸᧌��3��T0 k� �xr�|r&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��k]+�Mӷ᧌ ��3��T0 k� �xs�|s&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��l]'�M˶ᣌ ��3��T0 k� �tt�xt&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��l]#�Mǵ៌ ��3��T0 k� �tt�xt&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��m]#�	�ôᛌ ��3��T0 k� �tu�xu&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��nm�	���ᗌ ��3��T0 k� �pu�tu&�1D"3Q2	4#'Q  ��6    ����c� A^�A��N��A_��Y|C�A��nm�	���ᓌ ��3��T0 k� �pv�tv&�1D"3Q2	4#'Q  ��6    ����c� A^�A���N��A_��Y|C�A��om�	���ᓌ ��3��T0 k� �pw�tw&�1D"3Q2	4#'Q  ��6    ����c� A^�A���N��A_��Y|C�A��om�	���Ꮜ ��3��T0 k� �pw�tw&�1D"3Q2	4#'Q  ��6    ����c� A^�A���N��A_��Y|C�A��pm�	���ዌ ��3��T0 k� �lx�px&�1D"3Q2	4#'Q  ��6    ����c� A^�A���N��A_��Y|C�A��qm�	ͧ�� ��3��T0 k� �lx�px&�1D"3Q2	4#'Q  ��6    ����c� A^�A���N��A_��Y|C�A��qm�	ͣ��� ��3��T0 k� �ly�py&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_��Y|C�A��rm�	͟��{� ��3��T0 k� �lz�pz&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_��Y|C�A��rm�	͛��w� ��3��T0 k� �hz�lz&�1D"3Q2	4#'Q  ��6    ����c� A]��A��N��A_��Y|C�A��sm�	͛��s� ��3��T0 k� �h{�l{&�1D"3Q2	4#'Q  ��6    ����c� A]��A��N��A_��Y|C�A��sm�	����o� ��3��T0 k� �h{�l{&�1D"3Q2	4#'Q  ��6    ����c� A]��A��N��A_��Y|C�A��tm�	����g� ��3��T0 k� �h|�l|&�1D"3Q2	4#'Q  ��6    ����c� A]��A��N��A_��Y|C�A��tl��	����c� ��3��T0 k� �d|�h|&�1D"3Q2	4#'Q  ��6    ����c� A]��A��N��A_��Y|C�A�|ul��	����_� ��3��T0 k� �d}�h}&�1D"3Q2	4#'Q  ��6    ����c� A]��A��N��A_��Y|C�A�|ul��	����W� �3��T0 k� �d}�h}&�1D"3Q2	4#'Q  ��6    ����c� A]��A��N��A_��Y|C�A�|vl��	͋��S� {�3��T0 k� �d~�h~&�1D"3Q2	4#'Q  ��6    ����c� A]��A��N��A_��Y|C�A�|vl��	͋�K� w�3��T0 k� �`~�d~&�1D"3Q2	4#'Q  ��6    ����c� A]�A��N��A_��Y|C�A�xwl��	͇�G� o�3��T0 k� �`�d&�1D"3Q2	4#'Q  ��6    ����c� A]�A��N��A_��Y|C�A�xwl�	͇�?� k�3��T0 k� �`�d&�1D"3Q2	4#'Q  ��6    ����c� A]�A��N��A_��Y|C�A�xxl�	͇�;� g�3��T0 k� �`��d�&�1D"3Q2	4#'Q  ��6    ����c� A]�A��N��A_��Y|C�A�xxl�	���3� c�3��T0 k� �`��d�&�1D"3Q2	4#'Q  ��6    ����c� A]�A��N��A_��Y|C�A�xyl�	���/� _�3��T0 k� �\��`�&�1D"3Q2	4#'Q  ��6    ����c� A]�A��N��A_��Y|C�A�tyl�	���'� [�3��T0 k� �\��`�&�1D"3Q2	4#'Q  ��6    ����c� A]�A��N��A_��Y|C�A�tyl�	���� S�3��T0 k� �\��`�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�߈N��A_��Y|C�A�tzl�	���� O�3��T0 k� �\��`�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�߈N��A_��Y|C�A�tzl�	̓�� K�3��T0 k� �\��`�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�߈N��A_��Y|C�A�t{l�	̓�� G�3��T0 k� �X��\�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�ۈN��A_��Y|C�A�p{l�	̓�� C�3��T0 k� �X��\�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�ۈN��A_��Y|C�A�p|lߘ	̓��� ?�3��T0 k� �X��\�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�ۈN��A_��Y|C�A�p|lߗ	̓��� ;�3��T0 k� �X��\�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�ۈN��A_��Y|C�A�p|lۖ���� 7�3��T0 k� �X��\�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�׈N��A_��Y|C�A�p}lە���� 3�3��T0 k� �X��\�&�1D"3Q2	4#'Q  ��6   ����c� A]�A�׉N��A_��Y|C�A�p}lה���ߎ /�3��T0 k� �T��X�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�׉N��A_��Y|C�A�l}lד���׎ +�3��T0 k� �T��X�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�׉N��A_��Y|C�A�l~lג���ώ '�3��T0 k� �T��X�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�ӉN��A_��Y|C�A�l~lӑ]���� #�3��T0 k� �T��X�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�ӉN��A_��Y|C�A�llϐ]�����3��T0 k� �T��X�&�1D"3Q2	4#'Q  ��6    ����c� A]�A�ӉN��A_��Y|C�A�llϏ]��೎�3��T0 k� �P��T�&�1D"3Q2	4#'Q  ��6    ����c� A]ߨA�ωN��A_��Y|C�A�l~lώ]��૏�3��T0 k� �P��T�&�1D"3Q2	4#'Q  ��6    ����c� A]ߨA�ωN��A_��Y|C�A�h~lˍ]��࣏�3��T0 k� �P��T�&�1D"3Q2	4#'Q  ��6    ����c� A]ߨA�ωN��A_��Y|C�A�h~\ˌ]������3��T0 k� �P��T�&�1D"3Q2	4#'Q  ��6    ����c� A]ߨA�ωN��A_��Y|C�A�h~\ˌ]������3��T0 k� �P��T�&�1D"3Q2	4#'Q  ��6    ����c� A]ߨA�ωN��A_��Y|C�A�h}\ǋ]�������3��T0 k� �P��T�&�1D"3Q2	4#'Q  ��6    ����c� A]ۨA�ˉN��A_��Y|C�A�h}\Ǌ]�������3��T0 k� �P��T�&�1D"3Q2	4#'Q  ��6    ����c� A]ۨA�ˉN��A_��Y|C�A�h}\É]���{���3��T0 k� �L��P�&�1D"3Q2	4#'Q  ��6    ����c� A]ۨA�ˉN��A_��Y|C�A�h}\É]���s����3��T0 k� �L��P�&�1D"3Q2	4#'Q  ��6    ����c� A]ۨA�ˉN��A_��Y|C�A�d|�È���k����3��T0 k� �L��P�&�1D"3Q2	4#'Q  ��6    ����c� A]ۧA�ǉN��A_��Y|C�A�d|������c����3��T0 k� �L��P�&�1D"3Q2	4#'Q  ��6    ����c� A]ۧA�ǉN��A_��Y|C�A�d|������[����3��T0 k� �L��P�&�1D"3Q2	4#'Q  ��6    ����c� A]קA�ǊN��A_��Y|C�A�d|������S����3��T0 k� �L��P�&�1D"3Q2	4#'Q  ��6    ����c� A]קA�ǊN��A_��Y|C�A�d|������K����3��T0 k� �L��P�&�1D"3Q2	4#'Q  ��6    ����c� A]קA�ǊN��A_��Y|C�A�d{�����C����3��T0 k� �L��P�&�1D"3Q2	4#'Q  ��6    ����c� A]קA�ÊN��A_��Y|C�A�d{�����;����3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]קA�ÊN��A_��Y|C�A�d{�����3����3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]קA�ÊN��A_��Y|C�A�`{�����+����3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ӧA�ÊN��A_��Y|C�A�`{�����#����3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ӧA�ÊN��A_��Y|C�A�`zL���������3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ӧA�ÊN��A_��Y|C�A�`zL���������3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ӧA���N��A_��Y|C�A�`zL�� ��������3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ӧA���N��A_��Y|C�A�`zL�� ��������3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ӧA���NÍA_��Y|C�A�`zL�� ��������3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ӧA���NÍA_��Y|C�A�`z �� �������3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]ӧA���NÍA_��Y|C�A�`y �� �������3��T0 k� �D�H&�1D"3Q2	4#'Q  ��6    ����c� A]ϦA���NÍA_��Y|C�A�\y �� �������3��T0 k� �D�H&�1D"3Q2	4#'Q  ��6    ����c� A]ϦA���NÎA_��Y|C�A�\y �� ���ې���3��T0 k� �D�H&�1D"3Q2	4#'Q  ��6    ����c� A]ϦA���NÎA_��Y|C�A�\y �� ���Ӑ��3��T0 k� �D�H&�1D"3Q2	4#'Q  ��6    ����c� A]ϦA���NÎA_��Y|C�A�\y��� ���ː��3��T0 k� �D�H&�1D"3Q2	4#'Q  ��6    ����c� A]ϦA���NÎA_��Y|C�A�\y�Ë ���Ð��3��T0 k� �D�H&�1D"3Q2	4#'Q  ��6    ����c� A]ϦA���NÎA_��Y|C�A�\x�Ë �������3��T0 k� �D~�H~&�1D"3Q2	4#'Q  ��6    ����c� A]ϦA���NÎA_��Y|C�A�\x�ǋ �������3��T0 k� �D~�H~&�1D"3Q2	4#'Q  ��6    ����c� A]ϦA���NÎA_��Y|C�A�\x�ˋ �����ߣ�3��T0 k� �D~�H~&�1D"3Q2	4#'Q  ��6    ����c� A]˦A���NÏA_��Y|C�A�\x�ˋ �����ߟ�3��T0 k� �@~�D~&�1D"3Q2	4#'Q  ��6    ����c� A]˦A���NÏA_��Y|C�A�\x�ϋ݃���ߛ�3��T0 k� �@~�D~&�1D"3Q2	4#'Q  ��6    ����c� A]˦A���NÏA_��Y|C�A�\x�Ӌ݃���ߓ�3��T0 k� �@~�D~&�1D"3Q2	4#'Q  ��6    ����c� A]˦A���NÏA_��Y|C�M=Xx�׋݃���ߏ�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]˦A���NÏA_��Y|C�M=Xw�ۋ݃���߇�3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]˦A���NÏA_��Y|C�M=Xw�ۋ݃��߃�3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]˦A���NÏA_��Y|C�M=Xw�ߌ݃�w��{�3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]˦A���NǐA_��Y|C�M=Xw��݃�o��w�3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6   ����c� A]˦A���NǐA_�Y|C�M=Xv��݃�g��o�3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]˦A���NǐA_�Y|C�M=Xv��݃�_��k�3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ǦA���NǐA_�Y|C�M=Xv��݃�W��c�3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ǦA���NǐA_{�Y|C�M=Xv��݃��O��[�3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ǦA���NǐA_{�Y|C�M=Xu���݃��G�?W�3��T0 k� �H��L�&�1D"3Q2	4#'Q  ��6    ����c� A]ǦA���NǐA_{�Y|C�MMXu���݃��?�?O�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]ǥA���NǑA_w�Y|C�MMXu��݃��7�?K�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]ǥA���NǑA_w�Y|C�MMXu��탫�/�?C�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]ǥA���NǑA_w�Y|C�MMXt��탫�'�?;�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]ǥA���NǑA_s�Y|C�MMTt��탫��?7�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]ǥA���NǑA_s�Y|C�MMTt��탫��?/�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]ǥA���NǑA_s�Y|C�MMTt��탫��?+�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]ǥA���NǑA_o�Y|C�MMTs��탫��?#�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���NǑA_o�Y|C�MMTs#�탫��?�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���NÑA_o�Y|C�M=Ts'�탫��?�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���NÒA_k�Y|C�M=Ts+�탫��?�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A_k�Y|C�M=Ts3�탫��?�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A_k�Y|C�M=Tr7�탫���?�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A_k�Y|C�M=Tr	=;�탫���?�3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A_g�Y|C�M=Tr	=?�탫���>��3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A_g�Y|C�M=Tr	=C�탫��>��3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A_g�Y|C�M=Tr	=G�탫�N��3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A_c�Y|C�M=Tq	=G�탫�N��3��T0 k� �D��H�&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A_c�Y|C�A�Tq	MK�탫�N��3��T0 k� �@�D&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A_c�Y|C�A�Tq	MO�탫�N��3��T0 k� �<}�@}&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A_c�Y|C�A�Tq	MS�탫�N��3��T0 k� �<|�@|&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A__�Y|C�A�Tq	MS�탫�N��3��T0 k� �<z�@z&�1D"3Q2	4#'Q  ��6    ����c� A]åA���N��A__�Y|C�A�Pp	MW�탫�N��3��T0 k� �8y�<y&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A__�Y|C�A�Pp	=W�탫ߐN��3��T0 k� �8x�<x&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A__�Y|C�A�Pp	=[�탫ߐN��3��T0 k� �8x�<x&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A__�Y|C�A�Pp	=[�탫ېN��3��T0 k� �8x�<x&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_[�Y|C�A�Pp	=_�탫אN��3��T0 k� �8x�<x&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_[�Y|C�A�Pp	=_�탫אN��3��T0 k� �8w�<w&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_[�Y|C�A�Po	M_�탫ӐN��3��T0 k� �8w�<w&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_[�Y|C�A�Po	Mc�탫ϐN��3��T0 k� �8w�<w&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_W�Y|C�A�Po	Mc�탫.ϐN��3��T0 k� �8w�<w&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_W�Y|C�A�Po	Mc�탫.ːN��3��T0 k� �8w�<w&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_W�Y|C�A�Po	Mc�탫.ːN��3��T0 k� �8w�<w&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_W�Y|C�A�Po	=c�탫.ǐN��3��T0 k� �8w�<w&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_W�Y|C�A�Pn	=g�탫.ÐN��3��T0 k� �8v�<v&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_S�Y|C�A�Pn	=g�탫.ÐN��3��T0 k� �8v�<v&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N��A_S�Y|C�A�Pn	=g�탫.��N��3��T0 k� �8v�<v&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N�A_S�Y|C�A�Pn	=g�탫.��N��3��T0 k� �8v�<v&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N�A_S�Y|C�A�Pn�g�탫.��N��3��T0 k� �8v�<v&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N{�A_S�Y|C�A�Pn�k�탫.��N��3��T0 k� �4v�8v&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N{�A_O�Y|C�A�Pn�k�탫.��N��3��T0 k� �4v�8v&�1D"3Q2	4#'Q  ��6   ����c� A]��A���Nw�A_O�Y|C�A�Pn�o�탫.��N��3��T0 k� �4u�8u&�1D"3Q2	4#'Q  ��6    ����c� A]��A���Nw�A_O�Y|C�A�Pm�o�탫.��N��3��T0 k� �4u�8u&�1D"3Q2	4#'Q  ��6    ����c� A]��A���Ns�A_O�Y|C�A�Pm�o�݃�.��N��3��T0 k� �4u�8u&�1D"3Q2	4#'Q  ��6    ����c� A]��A���Ns�A_O�Y|C�A�Pm�s�݃�.��N�3��T0 k� �4u�8u&�1D"3Q2	4#'Q  ��6    ����c� A]��A���No�A_O�Y|C�A�Pm�w�݃�.��N{�3��T0 k� �4u�8u&�1D"3Q2	4#'Q  ��6    ����c� A]��A���No�A_K�Y|C�A�Pmw�݃�.��N{�3��T0 k� �4u�8u&�1D"3Q2	4#'Q  ��6    ����c� A]��A���Nk�A_K�Y|C�A�Pmw�݃�.��Nw�3��T0 k� �4u�8u&�1D"3Q2	4#'Q  ��6    ����c� A]��A���Nk�A_K�Y|C�A�Pm{�݃�.��Ns�3��T0 k� �4u�8u&�1D"3Q2	4#'Q  ��6    ����c� A]��A���Ng�A_K�Y|C�A�Lm{�݃�.��No�3��T0 k� �4t�8t&�1D"3Q2	4#'Q  ��6    ����c� A]��A���Ng�A_K�Y|C�A�Ll{�݃�.��No�3��T0 k� �4t�8t&�1D"3Q2	4#'Q  ��6    ����c� A]��A���Ng�A_K�Y|C�A�Ll{�݃�.��Nk�3��T0 k� �4t�8t&�1D"3Q2	4#'Q  ��6    ����c� A]��A���Nc�A_K�Y|C�A�Ll�݃�.��Ng�3��T0 k� �4t�8t&�1D"3Q2	4#'Q  ��6    ����c� A]��A���Nc�A_G�Y|C�A�Ll�݃�.��Nc�3��T0 k� �4t�8t&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N_�A_G�Y|C�A�Ll�݃�.��Nc�3��T0 k� �4t�8t&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N_�A_G�Y|C�A�Ll� ���.��N_�3��T0 k� �4t�8t&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N_�A_G�Y|C�A�Ll� ���.��N[�3��T0 k� �4t�8t&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N[�A_G�Y|C�A�Ll m� ���.��>[�3��T0 k� �4t�8t&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N[�A_G�Y|C�A�Ll m� ���.��>W�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���N[�A_G�Y|C�A�Ll m� ���.��>S�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NW�A_C�Y|C�A�Lk m� ���.��>S�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NW�A_C�Y|C�A�Lk m� ���.��>O�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NS�A_C�Y|C�A�Lk �� ���.��>K�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NS�A_C�Y|C�A�Lk �� ���.��>K�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NS�A_C�Y|C�A�Lk �� ���.��>G�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NO�A_C�Y|C�A�Lk �� ���.��>C�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NO�A_C�Y|C�A�Lk �� ���.��>C�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NO�A_C�Y|C�A�Lk �� ���.��>?�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NK�A_C�Y|C�A�Lk �� ���.��>;�3��T0 k� �4s�8s&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NK�A_?�Y|C�A�Lk �� ���.��>7�3��T0 k� �4r�8r&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NK�A_?�Y|C�A�Lk �� ���.��>7�3��T0 k� �4r�8r&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NK�A_?�Y|C�A�Lj �� �����>3�3��T0 k� �4r�8r&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NG�A_?�Y|C�A�Lj �� �����>/�3��T0 k� �4r�8r&�1D"3Q2	4#'Q  ��6   ����c� A]��A���NG�A_?�Y|C�A�Lj �� �����>+�3��T0 k� �4r�8r&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NG�A_?�Y|C�A�Lj�� �����>'�3��T0 k� �4r�8r&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NC�A_?�Y|C�A�Lj�� ����N#�3��T0 k� �4r�8r&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NC�A_?�Y|C�A�Lj�� ����N�3��T0 k� �4r�8r&�1D"3Q2	4#'Q  ��6    ����c� A]��A���NC�A_?�Y|C�A�Lj�� �����N�3��T0 k� �4r�8r&�1D"3Q2	4#'Q  ��6    ����c���E�˹B��;�{�E@��ZlC�E�#�%/�rh�D�8e3��T0 k� ������&�1D"3Q2	4#'Q  ��  	   ��� ����E�ӷB��<�{�E0��ZlC�E�+�%3�rx�E�@f3��T0 k� ����&�1D"3Q2	4#'Q  ��  	   ��� ����E�׵E��=�{�E0��ZlC�E�+�%3�r|�E�Dg3��T0 k� ����&�1D"3Q2	4#'Q  ��  	   ��� ����E�۴E��=��E0��ZlC�E�/�%3�r��F�Hg3��T0 k� ����&�1D"3Q2	4#'Q  ��  	   ��� ����E�߳E��>��E0��ZlC�E�3�%!7�r��F�Lh3��T0 k� ����&�1D"3Q2	4#'Q  ��  	   ��� ���E��E��>��E0��ZlC�E�7�%!7�r��G�Ph3��T0 k� ���#�&�1D"3Q2	4#'Q  ��  	   ��� ���E��E��>���E0��ZlC�E�7�%!7�r��G�Th3��T0 k� �'��+�&�1D"3Q2	4#'Q  ��  	   ��� ���E��E��>���E0��b�C�E�;�%!;���H�\i3��T0 k� �3��7�&�1D"3Q2	4#'Q  ��  	   ��� ���E��E��>���E0��b�C�E�?�%!;���I�`i3��T0 k� �;��?�&�1D"3Q2	4#'Q  ��  	   ��� ��'�E��E��>���E0��b�C�E�?�%!;���I�di3��T0 k� �?��C�&�1D"3Q2	4#'Q  ��  	   ��� ��+�E��E��>���E0��b�C�E�?�%!;���J�li3��T0 k� �G��K�&�1D"3Q2	4#'Q  ��  	   ��� ��3�E��E��>���E ��b�C�E�?�%!;���J�pi3��T0 k� �O��S�&�1D"3Q2	4#'Q  ��  	   ��� ��;�E��CB�>���E ��b�C�E�?�%!?����K�ti3��T0 k� �S��W�&�1D"3Q2	4#'Q  ��  	   ��� ��C�E��CB�=���E ��b�C�E�?��?����K�xi3��T0 k� �[��_�&�1D"3Q2	4#'Q  ��  
   ��� ��G�E��CB�=��E ��b�C�E�?��?���%�K�|i3��T0 k� �c��g�&�1D"3Q2	4#'Q  ��  
   ��� ��W�E��CB�<��E ��b�C�E�?��C���%�L��i3��T0 k� �s��w�&�1D"3Q2	4#'Q  ��  
   ��� ��_�E��CB�;��E ��ZlC�E�?��C���%� M��i3��T0 k� �w��{�&�1D"3Q2	4#'Q  ��  
   ��� ��g�E��CB�;��E ��ZlC�E�?��G���%� M��i3��T0 k� �����&�1D"3Q2	4#'Q  ��  
   ��� ��k�E��CB�:Q��E �ZlC�E�;��G���%��M��i3��T0 k� �{���&�1D"3Q2	4#'Q  ��  
   ��� ��s�E��CB�9Q��E �ZlC�E�;��K���%��N��i3��T0 k� �{���&�1D"3Q2	4#'Q  ��  
   ��� ��{�D3�CB�9Q��E {�ZlC�D4;��K���%��N��h3��T0 k� �{���&�1D"3Q2	4#'Q  ��  
   ��� ����D3�CB�8Q��E {�ZlC�D47��O���%��Nr�h3��T0 k� �����&�1D"3Q2	4#'Q  ��  
   ��� � �D3�CR�6��Ew�ZlC�D47��S�� %��Or�g3��T0 k� ������&�1D"3Q2	4#'Q  ��  
   ��� � �D3�CR�5��Ew�ZlC�D43��S��%��Or�g3��T0 k� ������&�1D"3Q2	4#'Q  ��  
   ��� � �D3�CR�4��Es�ZlC�D4/��W��%��Pr�f3��T0 k� ������&�1D"3Q2	4#'Q  ��  
   ��� � £�D3�CR�3��Es�ZlC�D4/��[��%��Pr�f3��T0 k� ������&�1D"3Q2	4#'Q  ��  
   ��� � «�E��CR�2��Es�b�C�D4+��_��%��Pr�e3��T0 k� ������&�1D"3Q2	4#'Q  ��  
   ��� � ¯�E��CR�1A��Es�b�C�D4+��_��%��Qr�d3��T0 k� ������&�1D"3Q2	4#'Q  ��  
   ��� � ·�E��CR�0A��Es�b�C�D4'��c��%��Qr�d3��T0 k� ������&�1D"3Q2	4#'Q  ��  
   ��� � ���E�ۙCR�-A��Es�b�C�D4#��k��$%��Rr�b3��T0 k� ������&�1D"3Q2	4#'Q  �  
   ��� ���E�ۙCR�,A��B�s�b�C�DD��o��(%��R��b3��T0 k� �����&�1D"3Q2	4#'Q  �� 
   ��� ���E�יCb�*A��B�w�b�C�DD�!s��,%��R��b3��T0 k� �s��w�&�1D"3Q2	4#'Q  �� 
   ��� ���E�ӘCb�)��B�w�b�C�DD�!w��0%��Q��b3��T0 k� �g��k�&�1D"3Q2	4#'Q  ��O 
   ��� ���E�ӘCb�'��B�w�b�C�DD�!{��4%��Q��b3��T0 k� �W��[�&�1D"3Q2	4#'Q  ��O 
   ��� ���E�ϙCb�&��B�{�b�C�DD�!��8%��Q��b3��T0 k� �K��O�&�1D"3Q2	4#'Q  ��O 
   ��� ���E�˙Cb�%��E{�b�C�DD�!���<%��P��a3��T0 k� �;��?�&�1D"3Q2	4#'Q  ��O    ��� ���E�˙IR�$��E{�ZlC�DD����@%��P��a3��T0 k� �/��3�&�1D"3Q2	4#'Q  ��O    ��� ���D�ǙIR�#��E�ZlC�DD���sD%��P��`3��T0 k� �#��'�&�1D"3Q2	4#'Q  ��O    ��� ���D���IR� ��E��ZlC�DD���sH%��O��`3��T0 k� ����&�1D"3Q2	4#'Q  ��O    ��� ���D���IR���E���ZlC�DC����sL��O��_3��T0 k� ������&�1D"3Q2	4#'Q  ��O    ��� �#�D���Ib���E���ZlC�DS����sP��N��^3��T0 k� ������&�1D"3Q2	4#'Q  ��O    ��� �#�D���Ib���E���ZlC�DS����cT��N� ^3��T0 k� ������&�1D"3Q2	4#'Q  ��O    ��� �#�D���Ib���E���ZlC�DS���cX��M�\3��T0 k� ������&�1D"3Q2	4#'Q  ��G    ��� �#�D���Ib� ���E���ZlC�DS����c\��L�[3��T0 k� ������&�1D"3Q2	4#'Q  ��G    ��� �#�D���IR� ���E���ZlC�ES����c\��K�[3��T0 k� ������&�1D"3Q2	4#'Q  ��G    ��� �#'�D���IR� ���E���ZlC�ES����c`��J�Y3��T0 k� ������&�1D"3Q2	4#'Q  ��G    ��� �#+�D���IR� ���E���ZlC�ESߜ���cd��I�X3��T0 k� ������&�1D"3Q2	4#'Q  ��G    ��� �#/�D���IR����E���ZlC�ESۜ���Sd��H�W3��T0 k� ������&�1D"3Q2	4#'Q  ��G    ��� �#3�D���E�����E���ZlC�ESם���Sh
��H�V3��T0 k� ������&�1D"3Q2	4#'Q  ��G    ��� �#?�Ec��E�����E���ZlC�ESם���Sh	��F� T3��T0 k� ������&�1D"3Q2	4#'Q  ��G    ��� �#C�Ec��E�����B�ZlC�ESӝ���Sh��E�$S3��T0 k� ����&�1D"3Q2	4#'Q  ��G    ��� �#G�Ec��E��я�B�ǧZlC�ES˝���Sh��D�$Q3��T0 k� ����&�1D"3Q2	4#'Q  ��G    ��� �#K�Ec��E��ы�B�˦ZlC�C�Ǟ���Sh��C�(P3��T0 k� ����&�1D"3Q2	4#'Q  ��G    ��� �#O�Ec��E��ы�B�ϥZlC�C㿞r�Sh��B�,O"���T0 k� ����&�1D"3Q2	4#'Q  ��G    ��� �#W�Ec{�E��ч�E�ۢZlC�C㳟r��h��?�0L"���T0 k� ���#�&�1D"3Q2	4#'Q  ��G    ��� �#[�D3w�E����E�ߡZlC�C㯟r��d��>�0K"���T0 k� �'��+�&�1D"3Q2	4#'Q  ��G    ��� �#_�D3o�E����E��ZlC�C㧠r��d��=�4I"���T0 k� �/��3�&�1D"3Q2	4#'Q  ��G    ��� ��c�D3k�E����E��ZlC�C㟠r#��d��;�8H"���T0 k� �3��7�&�1D"3Q2	4#'Q  ��G    ��� ��k�D3c�E���w�E���ZlC�C㓡r3��`��9�<E"���T0 k� �?��C�&�1D"3Q2	4#'Q  ��G    ��� ��o�D3[�E���s�E���ZlC�C㋡r7��\��7�<D"���T0 k� �G��K�&�1D"3Q2	4#'Q  ��G    ��� ��s�D3W�E���o�B��ZlC�Cモr?��\��6�@B"���T0 k� �O��S�&�1D"3Q2	4#'Q  ��G    ��� ��w�D3S�E���k�B��ZlC�C�{�rC��X��4�@@"���T0 k� �S��W�&�1D"3Q2	4#'Q  ��G    ��� ���D3G�E���c�B��ZlC�C�k�rO��P ��1�H=3��T0 k� �_��c�&�1D"3Q2	4#'Q  ��G    ��� ����D3?�E�� �_�B��ZlC�C�c�rS��P ��0�H;3��T0 k� �c��g�&�1D"3Q2	4#'Q  ��G    ��� ����D3;�E����W�E!�ZlC�C�[�r[��O���.�L:3��T0 k� �k��o�&�1D"3Q2	4#'Q  ��G    ��� ����Ec3�E����S�E!'�ZlC�C�S�r_��O���,�L83��T0 k� �o��s�&�1D"3Q2	4#'Q  ��G    ��� ����Ec'�C����G�E!/�ZlC�C�C�rk��G���)�P43��T0 k� �{���&�1D"3Q2	4#'Q  ��G    ��� �Ó�Ec#�C����C�E!7�ZlC�C�7�bo��G���'�T23��T0 k� �o��s�&�1D"3Q2	4#'Q  ��G    ��� �Ó�Ec�C����;�E;�ZlC�C�/�bs��G���%�T03��T0 k� �k��o�&�1D"3Q2	4#'Q  ��G    ��� �×�Ec�C���7�EC�ZlC�C�'�b{��C���#�X.3��T0 k� �g��k�&�1D"3Q2	4#'Q  ��G    ��� �Û�Ec�C���+�EO�ZlC�C��b{��?�� �\+3��T0 k� �g��k�&�1D"3Q2	4#'Q  �G    ��� �ß�Ec�C���#�ES�ZlC�D�b{��?���\)"s��T0 k� �_��c�&�1D"3Q2	4#'Q  ��    ��� �ß�Eb��C����I[�ZlC�D�b{��?��	�`'"s��T0 k� �[��_�&�1D"3Q2	4#'Q  ��    ��� �ß�Eb��C����I_�ZlC�D��b{�;��	�`%"s��T0 k� �W��[�&�1D"3Q2	4#'Q  ��    ��� �ß�Eb��C���Ik�ZlC�D�b{�;��	�d!"s��T0 k� �S��W�&�1D"3Q2	4#'Q  ��    ��� ����ER��C�� ��Io�ZlC�DۧR{�7��	�d"s��T0 k� �W��[�&�1D"3Q2	4#'Q  ��    ��� ����ER��C�� ��Is�ZlC�DӨRw�7��	�d"s��T0 k� �S��W�&�1D"3Q2	4#'Q  ��    ��� ����ER��C�� ��I!w�ZlC�D˨Rw�3��	�d"s��T0 k� �S��W�&�1D"3Q2	4#'Q  ��'    ��� ����ER��C�� ��I!��ZlC�D��Rs�/��	�h"s��T0 k� �O��S�&�1D"3Q2	4#'Q  ��'    ��� ����ER��EB�� ��I!��ZlC�D��Rs�+��
	�h"s��T0 k� �O��S�&�1D"3Q2	4#'Q  ��'    ��� ����ER��EB�� ��I!��ZlC�D��bo�'��	�h3��T0 k� �C��G�&�1D"3Q2	4#'Q  ��'    ��� ����C���EB�� ��I��ZlC�D��bo�#��sh3��T0 k� �7��;�&�1D"3Q2	4#'Q  ��'    ��� ����C��EB�� ��I��ZlC�D��bg���sh3��T0 k� �+��/�&�1D"3Q2	4#'Q  �'    ��� �ӗ�C��EB����I��ZlC�D��bg��� sd3��T0 k� �#��'�&�1D"3Q2	4#'Q  ��'    ��� �ӗ�C��EB����I��ZlC�Dw�bc����s`3��T0 k� ����&�1D"3Q2	4#'Q  ��'    ��� �ӛ�C��EB����E��ZlC�Do�b_�����\3��T0 k� ����&�1D"3Q2	4#'Q  ��'    ��� ~ӛ�E��EB����E��ZlC�D[�bW�����T
3��T0 k� ����&�1D"3Q2	4#'Q  ��'    ��� zӛ�E��C����E��ZlC�DS�bS������P	3��T0 k� ����&�1D"3Q2	4#'Q  ��'    ��� wӟ�E��C���w�E��ZlC�DK�bO������L3��T0 k� �����&�1D"3Q2	4#'Q  ��'    ��� tӟ�E��C���o�E��ZlC�C�?�bK������L3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� q��E��C���g�E��ZlC�C�7�rC������H3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� n��E�w�C���S�E��ZlC�C�#�r;�������@3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� j��E�w�C����K�E�ÂZlC�C��r7�������<3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� f��E�s�C����C�E�ǂZlC�C��r/�������8 3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� b��E�k�C����;�E�ςZlC�C��r'�������7�3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� ^��D2c�C����3�E�ӂZlC�C���r#�������3�3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� Z��D2c�C����#�E�ۂZlC�C��r����ҟ��/�3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� V��D2_�C�{���E��ZlC�C��r����қ��+�3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� R��D2W�C�w���E��ZlC�C�ۮr����қ��'�3��T0 k� ������&�1D"3Q2	4#'Q  ��'    ��� N                                                                                                                                                                            � � �  �  �  d A�  �K����   �      � \��� ]��� � �!  wj   
	     � �h      wj �h                          �         �     ���   0	&
         ��~�         ��oW�    ����oZ�    ����                  �         �     ���   (	          ��q    	    �g��    ����g��     ,��   	            �         �@  �  ���   0
          ����   $ $       ��W�    ���[����    ��   	             �$               ���   H	$
         ���\          /���    ���9��+j     ���   
              ���$          �     ���   03           ���� ��	      C�S    �����S                             ���E                ���    P		 5              j�P   
    W�Se�     j�>�Si�    ����               ' ���c         �  �  ��H  
	          ���6  � �  k�_E�    ���6�_E�                       	���c         `�   	  ��`  8	 

         ���      �`E�    ����`E�                      	���c         �     ��@   (
	          ���)  > � 
	   ���QH    ���)����      �                	���c         	 � �   
  ��@  0
3
         ��B   D D 
    ����B    ���`���"    ���                C���c         
 ��    ��@  8'
         ��_ ��     � ���    ��_ ���                            ���D             E  ��@    		 5 	                 ��      �                                                                           �                               ��        ���          ��                                                                 �                          rbu  ��        ��M�     rt��M�    ����                   x                j  �       �                          r    ��        ��N       r  �N                                                               �                          ��o�g������S�_�`���� ����M�N    
       	      
     ��� sp�A       )� `t� *D u� �D  n  �� n@ �� 0n` �  n� �D o ���X � �D l� Ƅ �o� Ǆ  p� �� q  �� q@ �  q`���� ���� ���� ����  ����. ����< ����J ����X � G _` G$ _� �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �d �Q����� ����� � 
�\ W� 
�< W� 
�\ X ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����c������ �  ������  
�fD
��L���"����D"� �  " `   J jF��    "�j "���
��
���     �j��  
  �
� �  �  
�  j    ��     ��S      ��    ��     ���       j    ��     ��S          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �6$      �� � �  ���        �t   ��        �        ��        �        ��        �    ��    ������H        ��                         T�) , � �����                                      �                ����             j�S ���&��  ���c���� � $          13 Teemu Selanne                                                                                    4  4     � �
�bE�E�$'KC0 KK))KL �kW� k_� �	ck � � 
ko � �cp � � cr � �cs � �cv � � cx � �c � � c� � �K � � K � �J� � � J� � �c� � � c� � �C � � C# � �c� � � c� � oK/ � K7"�� "�� � � �!
�� �""� � � #"� � �$"� � �%*� �&"�� '"�� �(� �)
��+ *"J }C+") uC  "P }; "= u � ."B }# /"Q }; "= u � 
� � � 
� � �3� � � 
� � 
�6� � 
�
 
�( 9"�:� � 
� �<!� p   "F x@>*9pP  *Hp                                                                                                                                                                                                                         �� P         �     @ 
             Y P E i  ��                    ������������������������������������� ���������	�
���������                                                                                          ��    �\?�� ��������������������������������������������������������   �4, J   * 4� K�� � @���@�A�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 	        @   $ 2    �� �:�J      e�                             ������������������������������������������������������                                                                                                                     	                   ����  ��                                             ��������� ���� � �������� �� ��������������������������������������������� ������� ����� ����������� ��������� �� ������������� �� ����� ��� ���������������������� ��� ��������� ������ �� ��������������������  �  �������������                                       *    �� �R�J                                     ������������������������������������������������������                                                                    	                                                                  ��������                                           ������������� ���� ������������������������������������������� ��� ��������� ����������������������������������������������� ���������������  ������������������������������� ����������� � ��������������������� ��� ���� ��������                                                                                                                                                                                                                                                                                               
                             �              


             �  }�           L+      0�  HC����  8���������������������������������������������������������������������������������  �          @u  J9     M                                                         ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � v�� �\                                                                                                                                                                                                                                                                                       )n)n1n  �              a      m            a            a      k                                                                                                                                                                                                                                                                                                                                                                                                         > �  >�  J�  (�  	(�  F_e�  �̞�X�˖������]�˖���� ]�̎��˖�[����.'                       e        $   �   &  QW  �   �                    �                                                                                                                                                                                                                                                                                                                                        K K           )             !��                                                                                                                                                                                                                            Z��   �� � ��      �� B      ��������� ���� � �������� �� ��������������������������������������������� ������� ����� ����������� ��������� �� ������������� �� ����� ��� ���������������������� ��� ��������� ������ �� ��������������������  �  �������������������������� ���� ������������������������������������������� ��� ��������� ����������������������������������������������� ���������������  ������������������������������� ����������� � ��������������������� ��� ���� ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ?   "   9   "   r                       f     �   �����J���J'      ��     b�   �         �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ��  � ��     � ��  � ��  p �� �� �z  p���� �$ ^h  ��  p  � \ ��   	 ��3h` �� �� �z ��   ��    ��   � �� �� �z   ����� �$ ��   � �� 1 �� �� �� ��  �� �� �  �� �� �z � ��� �$  � �  �� �  �      �       =���� e�����  g��� 	      f ^�         ��Q��      =      ���n���2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                                                  U  T   T   T     T UDUDDUDDDDDDDDDDDDDDDP   E�  DU� DDU�DDDUDDDDDDDDDDDD                UP  E�  E   E                                           ���U�UTD�DDDDDDTDD TDD   �   U_ DEU�DDDUDDDDD��DZT�DDDDDDDDDDDDTDDDDDDDDUTU�����DDDDDDDDDDDEDDDEDDDDTUTU�Ԫ���Z_   P   � �U�UTDUDDDDUTD�DT��D        U_��DEU_DDD_DDDPDDE�DDE  �DD DD DD �DD �UD  �U       DZTDEDDDDE�DDE�DDE�TDDT�DE�TE���DDTU�ZD���������DDTDD��ZT�T���ZTDDE��D��T�T��DUTTT��Z��TQTDDUTD�DDDTDDD�DDDDDDE�DD_TDE�DD_ DDP DDP DD_ DU_ U�  �                                       TE�DDD�UUU                    ���DDDUUUTD  D  D  D  D  U��D�TDDDDEUUDP  DP  DP  DP  UP  TDE�DDDPUUU_                                                    wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwtwwwCwwt1wwCwt1wC�t1��C1����������""""���������������!���""!����,���ww��7����������������wwwwwwwwwwwwwwwwwwww7wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwws��w1wt1�wC�t1��s��s��s������"$��Gw�!������������L���q��"r��������!�����!ww�r�w�ww!�wwrwwwwwwqwwwrwwww�7ww�ww�ww��7w��w���G��'!wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         7v` weV "fff"O�p"��p"��p"�p3�}p-��p=��p|� }�  }�  ��  ��  ��  ��  �  �  �  �  �  "              `  eV  fff O�  ��  ��  �  �} �� �� ��  |�  }�  ��    =   }   =   =              �������}�}�}�ww~r�� ∈�������������������}�� }�� ��� ��� ����   �   �   �   �   �   �   �   C""42""#2""#2""#2""#s3342"""3333    p   p   p   p   p   p   p    ��������� ��� }�� ��  ��  ����  ��  ��  ��  ��  ��  ��  ��                          � �� ��    "               wvf wfU 7Of`w��f"�� "�p-�}p���� ��� ����x��	�� �� �� "�        f  U` f` f` �p w���� `  eV  ff  O�  ��  �� ����}�                �  �  ��  �            �  �  �   �  ��  �                     �  �  �   � `  eV  ff  O�  ��  ��  ����}���������������p	���         `  eV  ff  O�  ��  ��  ���}�     �  �  �   �  ��  �   �            ��  ��  �   ��  �   ���������������p	���                    3333UUUU                        wwww                    333333333333333333333   w  G� ws@ ws� ws$7w@wwww"                               ����������� ��� �� ��  �    `  eV  ff  O�  ��  ��  � ��}�            """"                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                                                �����   �   �   �   ����                                     
�  

  
 � 
 
 
   
   
   
   
  ��                  ��   
   
   
   
   
   
 
 
 � 

  
�                 �   
    �   
    �   
    �   
   
   �  
   �  
   �  
   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "      " ""   "" !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """     " ""   "" !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "      " ""   "" !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        � ��~ ��. �r~ g~  ׮  
�  ��  �� ̾��� ��� ��� �� �� ��� �" "  �                           "   ¨�ˋ��˜��̌������ ��������˻�˻�����D���C��ET��EUZ�U ����Z� ��  �   �        "   "   "       �              �       33  DD3�DD;�3C��34��D� �U��� ��̰ �̰  ̊  ɫ  ��  ""  ""��"� �                                              .   .           �   �   �   �   �   �   �   �"" ""!! ��� �                      �   ��  "   "   �   "  "  "   �                                 �   ���                            �   "                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��                        �          �   � � /  �"" �"  �    "   "   "  �� ��                   �".��".���                                  �   �      ��   �  ��  �  �  �         � ".��".��/����  �                                                                                                                                        �� ��� ��� ww� &'� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                               " "/ �/� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   �".��".���                                ".  ".  ���  �   "  "  "   �                     ""  "".  . �    �                                                                                                                                            �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   �   " � ��      �    �      �                         ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �                    ".  ".  ���                                                                                                                                                                                                  	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��  ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  &'  vv  w                �                        ��"� �"� ����                            ".  ".  ���                                                                                                                                                                                                        �  �  �  �  w  �  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �           �   �     �   �                                                   �   �                               � ����ݼ� ����                                                                                                                                                                 �� ��� ��� ww� &'� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                               " "/ �/� ��    4U� 4U� 4U� 3UXP�EX��U����  ��                    �  ��� ݼ� �    �    �   �                     �         "   "   �                                     �  ��� ݼ� w{� &'� vw�      � ".��".��/����  �                � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                        
���	���̜̽�˽�̈ۻ��ۻ�۽��˲"������"���" ��"                "   "   "                 ���       "   "     ����           �  ��� ݼ� w�� b}� ggp wz�����""H�""T�B"UJ�"UJ�@T�DT�TUJ�  ��.�                           5J� �J� �˻ �˰ ʘ� ̪ ˲"�" ""�"" �  ��                /���"/�  ��                    �                                                                            �               �     "   "                   �     �                                       �   ���                            �   "                      ��   ��                  .  .  "  " ��                                                 �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��r`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   �". ". ����                /���"/�  ��                    �                                                                            �               �     "   "                �   "�  "�  "   /  "   ��  ��                    �   ���                            �   "                                                                                                     �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��  .�"." "."   /�  �  �              � ��         �� �� �� g} &' vw                     ".  ".  ���                   ���                                                                                                                                                                           ̰ ˻ ���wݛb}�gz� w��  ��  ��  ��  ��  ,�  "�  �  ,�  "�  ."  ."  "  "   !                        �   �   ̰  ��  ��  ��� ��� �ܘ �ل@�؊@�4�@�H�@�D �@ �H� "H�""C�"ˋ" �" ��" "��� �  �                     ��  �                            �         �           �       �                                      "  ."  �"    �          �� ̻� ��� ww� &'� vvw    �   �     �     �  �  "   "   "   "�  �                ���                                                                                                                                                                                                                     �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ���������""��""��""�����        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                               � ����ݼ� ����                                                                                                                                                                           2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ D�D D@                     �� ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�GwDGwqwDDwtwwww3333DDDD �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�""""����������A��I��I = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=""""�����A�DA�I��I�    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"��������I���I���I���I��� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(XxMAMAMMMM�M�M����3333DDDD w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xwwD�����MD��M����3333DDDD  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���4���4���4���4���4���43334DDDD �  + � � � � � � � � � � ��	� � � ��� � � � � � � � � � � ��	� � � ��� �� ����(+((�""""wwwwqqqqwGwGGG ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""wwwwwwqqDAwG M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M������������������333DDD � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�M��M��D��M����������3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DD��D�M��D����3333DDDD 5 6  X � �F � � � � � ����� � ����������� � ����� � � � � ��	F ��(X((6(5""""wwwwwwDGqGq x �  l � �G � � � � � � � � � � ������������� � � � � � � � � � ��	G ��l((�x""""wwwwwwwGqGqqD w w x y ������H���������������������������������H�����yxww""""wwwwwwwwGwwGwwGwwGw  � + w�������I�J�K�L�M�N�O � � � � � � � � � � � � � � � � � � � ��O�N�M�L�K�J�I������w(+�(DDwwwqwwGwtDGwwww3333DDDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A e ��A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,GwAqAADqtDGwwwww3333DDDD +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�] � ځ]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+www4www4www4Gww4Gww4www43334DDDD  � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� SA��(( """"���������M�MMM X � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� SA��(Xx""""�������A��AA w � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� )��:	9ww��������������333DDD � � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(I��I����������������3333DDDD  � �!�AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((���A���I��I���I�����3333DDDD m � �!�A�A� � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""������������������������  � �!�AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M""""������D�D��� 
 � �!�AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�""""������������������������ - � �!�!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�wqwwqwwwwwqwwwDwwww3333DDDD 69�:���  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5qqwwwDDwtGwwww3333DDDD x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xwww4www4www4www4www4www43334DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwqwwwqwqwq + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""wwwwwwwDwGwA � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(��A�L�L�L��L���333DDDLDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDD �
�bE�E�$'KC0 KK))KL �kW� k_� �	ck � � 
ko � �cp � � cr � �cs � �cv � � cx � �c � � c� � �K � � K � �J� � � J� � �c� � � c� � �C � � C# � �c� � � c� � oK/ � K7"�� "�� � � �!
�� �""� � � #"� � �$"� � �%*� �&"�� '"�� �(� �)
��+ *"J }C+") uC  "P }; "= u � ."B }# /"Q }; "= u � 
� � � 
� � �3� � � 
� � 
�6� � 
�
 
�( 9"�:� � 
� �<!� p   "F x@>*9pP  *Hp3333DDDDAqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD��������������������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ��������������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ��������������������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE��������������������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD��������������������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD��������������������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD��������������������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� ����7�\�J��<�V�I�P�[�H�P�S�S�L�������8�>�7���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� �� ��>�O�L�V�Y�L�U��1�S�L�\�Y�`�������8�>�7���""""������A�D��I��""""�������D����� ����>�L�L�T�\��=�L�S�H�U�U�L��������>��<���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �8�>�7��� ���A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �>��<�����""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,��,��,�D�,���#333DDDDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II�""""������D""""������IADD���I""""��������D��""""�������I��I�I�I�""""�������A�D�II�I""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            