GST@�                                                           �t�                                                      � ���      �  ��     	      ����e ����J�������ĸ��X�������        �g     #    ����                                d8<n    �  ?     bb����  �
fD�
�L���"����D"� j   " B   J  jF�"    
 �j� � 
 ���
��
�"    "D�j  �
`   "  ��
  ��                                                                              ����������������������������������      ��    bb= QQ0 4 111 44              		 

                     ��� �   � �                 nnn ))	         88�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             ��  )          == �����������������������������������������������������������������������������                                D              @  &   s   �                                                                                 '      )n)n	n  �)�    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    AR�xS��RDA B#��4Q��K��@^��"�C��3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�xS��RDAB#��4Q��K��?^��"�C��3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�xS��RDAB'��4Q��K��?^��"�C��3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�xS��RDAB'��4A��K��>^��"�C��3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�xS��RDAB+��4A��K��>^��"�C��3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�wS��RDAB+��4A��K��>^��"�C��3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�wS��RDAB/��4A{�K��=^��"�C��3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�wS��RDAB/��4As�K��=^��"�C��3��T0 k� �{���e2$ 4e2	d 3  ��H    ��� 8AR�wS��RDAB3��4�k�K��<^��"�C��3��T0 k� �s��w�e2$ 4e2	d 3  ��H    ��� 8AR�wS��RDAB3��4�c�K��<^��"�C��3��T0 k� �k��o�e2$ 4e2	d 3  ��H    ��� 8AR�wS��RDAB3��4�[�K��;^��"�C��3��T0 k� �k��o�e2$ 4e2	d 3 �H    ��� 8AR�wS��RDA B7��4�S�K��;Χ�"�K�3��T0 k� �g��k�e2$ 4e2	d 3 ��O    ��� 8AR�wS��RDA B7��4�K�K��;Σ�"�K�3��T0 k� �c��g�e2$ 4e2	d 3 ��O    ��� 8AR�wS��RHA B;��4�C�K�:Λ�"�K�3��T0 k� �c��g�e2$ 4e2	d 3 ��O   ��� 8AR�vS��RHA�B;��4�;�K�:Γ�"߇K�
3��T0 k� �_��c�e2$ 4e2	d 3 ��O    ��� 8AR�vS��RHA�B;��4�3�K�9Ώ�"߇K�
3��T0 k� �[��_�e2$ 4e2	d 3	 ��O   ��� 8AR�vS��RHA�B?��4�+�K�9·�"߈K�	3��T0 k� �[��_�e2$ 4e2	d 3 ��O    ��� 8AR�vS��RHA�B?��4�#�K�9��"ۈK�3��T0 k� �W��[�e2$ 4e2	d 3 ��O    ��� 8AR�vS��RHA�BC��4��K�8�{�"ۈK�3��T0 k� �S��W�e2$ 4e2	d 3 ��O    ��� 8AR�vS��RDA�BC��4��KЬ8�s�"ۈK�3��T0 k� �S��W�e2$ 4e2	d 3 ��O    ��� 8AR�vS��RDA�BC��4��KШ8�k�"ۈK�3��T0 k� �O��S�e2$ 4e2	d 3 ��O    ��� 8AR�vS��RDA�BG��4��KШ7�g�"׉K�3��T0 k� �O��S�e2$ 4e2	d 3 ��O    ��� 8AR�vS��R@A�BG��4�KФ7�_�"׉K�3��T0 k� �K��O�e2$ 4e2	d 3 ��O    ��� 8AR�vS��R@ A�BG��4 ��KР7�[�"׉K�3��T0 k� �G��K�e2$ 4e2	d 3 ��O    ��� 8AR�uS��R@ A��BK��4 ��KР6�S�"ӉK�|3��T0 k� �G��K�e2$ 4e2	d 3 ��O    ��� 8AR�uS��R< A��BK��4 �C@�6�O�ӉL|3��T0 k� �C��G�e2$ 4e2	d 3 ��O    ��� 8AR�uS��R< A��BK��4 �C@�5�K�ӉLx3��T0 k� �?��C�e2$ 4e2	d 3 ��O    ��� 8AR�uS��R< A��BO��4 �C@�5�C�ӊLx3��T0 k� �?��C�e2$ 4e2	d 3 ��O    ��� 8AR�uS��R< A��BO��4 ۏC@�4�?�ϊLx3��T0 k� �;��?�e2$ 4e2	d 3 ��O    ��� 8AR�uS��R8 A��BO��4 אC@�4�7�ϊLt3��T0 k� �7��;�e2$ 4e2	d 3 ��O   ��� 8AR�uS��R8 A��BS��4 ϐC@�3�3�ϊLt3��T0 k� �7��;�e2$ 4e2	d 3 ��O    ��� 8AR�uS��R7�A��BS��4 ːC@�2�/��ϊLt3��T0 k� 3��7�e2$ 4e2	d 3 ��O    ��� 8AR�uS��R7�A��BS��4 ÐC@�2�+��ˊLp3��T0 k� /��3�e2$ 4e2	d 3  ��O    ��� 8AR�uS��R7�A��BS��4 ��C@�1�#��ˋLp3��T0 k� /��3�e2$ 4e2	d 3" ��O    ��� 8AR�uS��R3�A��BW��4 ��KЈ0���ˋLp3��T0 k� +��/�e2$ 4e2	d 3# ��O    ��� 8AR�uS��R3�A��BW��4 ��KЄ/���ǋLl3��T0 k� +��/�e2$ 4e2	d 3$ ��O    ��� 8AR�tS��R3�A��BW��4 ��KЄ.���ǋLl3��T0 k� �'��+�e2$ 4e2	d 3% ��O    ��� 8AR�tS��R/�A��B[��4 ��KЀ.���ËLl3��T0 k� �#��'�e2$ 4e2	d 3& ��O    ��� 8AR�tS��R/�A��B[��4 ��KЀ-��⿋Ll3��T0 k� �#��'�e2$ 4e2	d 3' ��O    ��� 8AR�tS��R+�A��B[��4 ��K�|,��⿋Ll3��T0 k� ���#�e2$ 4e2	d 3( ��O    ��� 8AR�tS��R+�A��B[��4 ��K�|+��⻋Ll3��T0 k� ����e2$ 4e2	d 3) ��O    ��� 8AR�tS��R+�A��B_��4 ��K�x+���ⷌLh3��T0 k� ���e2$ 4e2	d 3* ��O    ��� 8AR�tS��R'�A��B_��4 ��K�x*���ⷌLh3��T0 k� ���e2$ 4e2	d 3* ��O    ��� 8AR�tS��R'�A��B_��4 ��K�t)]���Lh"s��T0 k� ���e2$ 4e2	d 3+ ��O    ��� 8AR�tS��R'�A��B_��4 ��K�t)]��Ld"s��T0 k� ���e2$ 4e2	d 3, ��O    ��� 8AR�tS��R'�A��Bc��4 ��K�p(]��Ld"s��T0 k� ���e2$ 4e2	d 3- ��O    ��� 8AR�tS��R#�A��Bc��4 �K�p']��Ld "s��T0 k� ����e2$ 4e2	d 3. ��O   ��� 8AR�tS��R#�A��Bc��4 w�K�l']��Ld "s��T0 k� ����e2$ 4e2	d 3. ��O    ��� 8AR�tS��R#�A��Bc��4 s�K�l&]߼�L` "s��T0 k� ����e2$ 4e2	d 3/ ��O    ��� 8AR�tS��R�A��Bc��4 o�K�l%]ۼ�L` "s��T0 k� ����e2$ 4e2	d 30 ��O    ��� 8AR�tS��R�A��Bg��4 k�K�h%]׼�Lc�"s��T0 k� ����e2$ 4e2	d 31 ��O    ��� 8AR�sS��R�A��Bg��4 g�K�h$]Ӽ�L_�"s��T0 k� �����e2$ 4e2	d 31 ��O    ��� 8AR�sS��R�A��Bg��4 c�K�d#]Ӽ�L_�"s��T0 k� �����e2$ 4e2	d 32 ��O    ��� 8AR�sS��R�A��Bg��4 _�K�d#]ϻ�L_�"s��T0 k� ������e2$ 4e2	d 32 ��O    ��� 8AR�sS��R�A��Bk��4 [�K�d"]˻��L_�3��T0 k� ������e2$ 4e2	d 33 ��O    ��� 8AR�sS��R�A��Bk��4 W�K�`"]ǻ��L[�3��T0 k� ������e2$ 4e2	d 33 ��O   ��� 8AR�sS��R�A��Bk��4 S�K�`!]û�L[�3��T0 k� �����e2$ 4e2	d 34 ��O    ��� 8AR�sS��R�A��Bk��4 O�K�\!]��w�L[�3��T0 k� ����e2$ 4e2	d 34 ��O    ��� 8AR�sS��R�A��Bk��4 K�K�\ ]��s�L[�3��T0 k� ����e2$ 4e2	d 35 ��O    ��� 8AR|sS��R�A��Bo��4 G�K�\ ]��o�LW�3��T0 k� ����e2$ 4e2	d 35 ��O    ��� 8AR|sS��R�A��Bo��4 C�K�X]��g�LW�3��T0 k� ����e2$ 4e2	d 36 ��O    ��� 8AR|sS��R�A��Bo��4 ?�K�X]��c�LW�3��T0 k� ����e2$ 4e2	d 36 ��O    ��� 8AR|sS��R�A��Bo��4 ?�K�X]��_�LW�3��T0 k� ����e2$ 4e2	d 36 ��O    ��� 8ARxsS��R�A��Bo��4�;�K�T]��W�LW�3��T0 k� ����e2$ 4e2	d 37 ��O    ��� 8ARxsS��R�A��Bs��4�7�K�T]��S�LS�3��T0 k� �߮��e2$ 4e2	d 37 ��O    ��� 8ARxsS��R�A��Bs��4�3�K�T]��K�LS�"���T0 k� �ۭ�߭e2$ 4e2	d 37 ��O   ��� 8ARxsS��R�A��Bs��4�/�K�P]��G�K�S�"���T0 k� �ۭ�߭e2$ 4e2	d 38 ��O    ��� 8ARxsS��R�A��Bs��4�+�K�P]��?�K�S�"���T0 k� �׭�ۭe2$ 4e2	d 38 ��O    ��� 8ARtsS��R�A��Bs��4�'�K�P]��;�K�S�"���T0 k� �Ӭ�׬e2$ 4e2	d 38 ��O    ��� 8ARtsS��R�A��Bs��4@'�K�L]��3�K�O�"���T0 k� �Ӭ�׬e2$ 4e2	d 38 ��O    ��� 8ARtsS��R�A��Bw��4@#�K�L]��/�K�O�"���T0 k� �ϫ�ӫe2$ 4e2	d 38 ��O   ��� 8ARtsS��R�A��Bw��4@�K�L]��'�K�O�"���T0 k� ϫ�ӫe2$ 4e2	d 38 ��O    ��� 8ARprS��R�A��Bw��4@�K�H]���C�O�"���T0 k� ˪�Ϫe2$ 4e2	d 39 ��O    ��� 8ARprS��R�A��Bw��4@�K�H]���C�O�"���T0 k� Ǫ�˪e2$ 4e2	d 39 ��O    ��� 8ARprS��R�A��Bw��40�K�H]���C�K�"���T0 k� ǩ�˩e2$ 4e2	d 39 ��O    ��� 8ARprS��R�A��Bw��40�K�H]���C�K�"���T0 k� é�ǩe2$ 4e2	d 39 ��O    ��� 8ARprS��R�A��B{��40�K�D]����C�K�3��T0 k� ݿ��èe2$ 4e2	d 39 ��O    ��� 8ARprS��R�A��B{��40�K�D]�����C�G�3��T0 k� ݿ��èe2$ 4e2	d 39 ��O    ��� 8ARlrS��R�A��B{��40�K�@]���C�G�3��T0 k� ݷ����e2$ 4e2	d 38 ��O    ��� 8ARlrS��R�A��B{��4?��K�@]{���C�G�3��T0 k� ݷ����e2$ 4e2	d 38 ��O    ��� 8ARlrS��R�A��B{��4?��K�@]{�QߐC�G�3��T0 k� �����e2$ 4e2	d 38 ��O    ��� 8ARlrS��Q��A��B{��4?��K�@]w�QאC�C�3��T0 k� �����e2$ 4e2	d 38 ��O    ��� 8ARlrS��Q��A��B��4?��K�<]w�QϐC�C�3��T0 k� �����e2$ 4e2	d 38 ��O    ��� 8ARhrS��Q��A��B��4?�K�<]s�QːC�?�3��T0 k� �����e2$ 4e2	d 37 ��O    ��� 8ARhrS��Q��A��B��4?�K�<]o�QÐC�?�3��T0 k� �����e2$ 4e2	d 37 ��O    ��� 8ARhrS��Q��A��B��4?�K�<]o�Q��C�?�3��T0 k� ������e2$ 4e2	d 37 ��O    ��� 8ARhrS��Q��A��B��4/�K�8]k�Q��C�?�3��T0 k� ������e2$ 4e2	d 37 ��O    ��� 8ARhrS��Q��A��B��4/�K�8]k�Q��C�;�3� T0 k� ������e2$ 4e2	d 36 ��O    ��� 8ARhrS��Q��A��B��4/�K�8]g�A��C�;�3� T0 k� ������e2$ 4e2	d 36 ��O    ��� 8ARdrS��Q��A��B��4/�K�8]g�A��C�;�3� T0 k� ������e2$ 4e2	d 35 ��O    ��� 8ARdrS��Q��A��B���4/ߦK�4]c�A��C�;�3� T0 k� ͛����e2$ 4e2	d 35 ��O    ��� 8ARdrS��Q��A��B���4/ߧK�4]c�A��C�7�3� T0 k� ͗����e2$ 4e2	d 35 ��O    ��� 8ARdrS��Q��A��B���4/ۨK�4]_�A��C�7�3� T0 k� ͓����e2$ 4e2	d 34 ��O    ��� 8ARdrS��Q��A��B���4/۩K�4]_�A{�C�7�3� T0 k� ͓����e2$ 4e2	d 34 ��O    ��� 8ARdrS��Q��A��B���4/۪C@4][�As�C�3�3� T0 k� ͏����e2$ 4e2	d 33 ��O    ��� 8ARdrS��Q��A��B���4/۬C@0][�Ak�C�3�3� T0 k� ݏ����e2$ 4e2	d 33 ��O    ��� 8AR`rS��Q��A��B���4׭C@0]W�Ac�C�/�3� T0 k� ݋����e2$ 4e2	d 32 ��O    ��� 8AR`rS��Q��A��B���4׮C@0]W�A[�C�+�3� T0 k� ݇����e2$ 4e2	d 31 ��O    ��� 8AR`rS��Q��A��B���4ׯC@0]S��S�C�'�3� T0 k� ݇����e2$ 4e2	d 31 ��O    ��� 8AR`rS��Q��A��B���4ױK�0]S��K�C�'�3� T0 k� ݃����e2$ 4e2	d 30 ��O    ��� 8AR`rS��Q��A��B���4ײK�,]S��C�C�#�3� T0 k� �����e2$ 4e2	d 3/ ��O    ��� 8AR`rS��Q��A��B���4�׳K�,]O��;�C��3� T0 k� �����e2$ 4e2	d 3/ ��O    ��� 8AR`rS��Q��A��B���4�۴K�,]O��3�C��3� T0 k� �{���e2$ 4e2	d 3. ��O    ��� 8AR`rS��Q��A��B���4�۵K�,]K�A+�C��3� T0 k� �w��{�e2$ 4e2	d 3- ��O    ��� 8AR`rS��Q��A��B���4�۶K�,]K�A#�C��3� T0 k� �w��{�e2$ 4e2	d 3, ��O    ��� 8AR\rS��Q��A��B���4�߷K�,]G�A�C��3� T0 k� �s��w�e2$ 4e2	d 3, ��O    ��� 8AR\rS��Q��A��B���4�߹K�(
]G�A�C��3� T0 k� �o��s�e2$ 4e2	d 3+ ��O    ��� 8AR\qS��Q��A��B���4��K�(
]G�A�C��3� T0 k� �o��s�e2$ 4e2	d 3* ��O    ��� 8AR\qS��Q��A��B���4��K�(	]C�A�C��3� T0 k� �k��o�e2$ 4e2	d 3) ��O    ��� 8AR\qS��Q��A��B���4��K�(	]C�@��C���3� T0 k� �k��o�e2$ 4e2	d 3( ��O    ��� 8AR\qS��Q��A��B���4��K�(]C�@��K���3� T0 k� g��k�e2$ 4e2	d 3' ��O    ��� 8AR\qS��Q��A��B���4��K�(]?�0�K���3� T0 k� c��g�e2$ 4e2	d 3& ��O    ��� 8AR\qS��Q��A��B���4��K�$]?�0�K���3� T0 k� c��g�e2$ 4e2	d 3% ��O    ��� 8AR\qS��Q��A��B���4���K�$];�0ߚK���3� T0 k� _��c�e2$ 4e2	d 3$ ��O    ��� 8ARXqS��Q��A��B���4���K�$];�0ۛK���3� T0 k� [��_�e2$ 4e2	d 3# ��O    ��� 8ARXqS��Q��A��B���4���K�$];�0ӜK���3� T0 k� �[��_�e2$ 4e2	d 3" ��O    ��� 8ARXqS��Q��A��B���4��K�$]7�0˝K���3� T0 k� �W��[�e2$ 4e2	d 3! ��O    ��� 8ARXqS��Q��A��B���4��K�$]7�0ǞK���3� T0 k� �S��W�e2$ 4e2	d 3  ��O    ��� 8ARXqS��Q��A��B���4�K�$]7�0��K���3� T0 k� �S��W�e2$ 4e2	d 3 ��O    ��� 8ARXqS��Q��A��B���4�K� ]3�з�K���3� T0 k� �O��S�e2$ 4e2	d 3 ��O    ��� 8ARXqS��Q��A��B���4�K� 3�г�K���3� T0 k� K��O�e2$ 4e2	d 3 ��O    ��� 8ARXqS��Q��A��B���4�K� 3�Ы�K���3� T0 k� K��O�e2$ 4e2	d 3 ��O    ��� 8ARXqS��Q��A��B���4��K� /�У�L��3� T0 k� G��K�e2$ 4e2	d 3 ��O    ��� 8ARXqS��Q��A��B���4��K� /�П�L��3� T0 k� G��K�e2$ 4e2	d 3 ��O   ��� 8ARXqS��Q��A��B���4��K� /�З�L��3� T0 k� C��G�e2$ 4e2	d 3 ��O    ��� 8ARXqS��Q��A��B���4�'�K� /�Г�L��3� T0 k� �?��C�e2$ 4e2	d 3 ��O    ��� 8ARTqS��Q��A��B���4�+�K�+�Ћ�L��3� T0 k� �?��C�e2$ 4e2	d 3 ��O    ��� 8ARTqS��Q��A��B���4�/�K�+�Ї�L��3� T0 k� �;��?�e2$ 4e2	d 3 ��O    ��� 8ARTqS��Q��A��B���4�7�K�+�Ѓ�L��3� T0 k� �7��;�e2$ 4e2	d 3 ��O    ��� 8ARTqS��Q��A��B���4�;�K� '��{�L��3� T0 k� �7��;�e2$ 4e2	d 3 ��O    ��� 8ARTqS��Q��A��B���4�?�K� -'��w�L��3� T0 k� �3��7�e2$ 4e2	d 3 ��O    ��� 8ARTqS��Q��A��B���4�G�K� -'��o�L��3� T0 k� �/��3�e2$ 4e2	d 3 ��O    ��� 8ARTqS��Q��A��B���4�K�K��-'��k�L��3� T0 k� �/��3�e2$ 4e2	d 3 ��O    ��� 8ARTqS�Q��A��B���4�S�K��-#��g�L��3� T0 k� �+��/�e2$ 4e2	d 3
 ��O    ��� 8ARTqS�Q��A��B���4�W�K��-#��c�L��3� T0 k� �+��/�e2$ 4e2	d 3 ��O    ��� 8ARTqS�Q��A��B���4�_�K��-#��[�L��3� T0 k� �'��+�e2$ 4e2	d 3 ��O    ��� 8ARTqS�Q��A��B���4�c�K��-#��W�L��3� T0 k� �#��'�e2$ 4e2	d 3 ��O    ��� 8ARTqS�Q��A��B���4�k�K��-��S�L��3� T0 k� �#��'�e2$ 4e2	d 3 ��O    ��� 8ARTqS�Q��A��B���4�o�K��-��O�L��3� T0 k� ���#�e2$ 4e2	d 3 ��O    ��� 8ARTqS�Q��A��B���4�w�K����G�L��3� T0 k� ����e2$ 4e2	d 3  ��O   ��� 8ARPqS�Q��A��B���4p{�K����C�L��3� T0 k� ����e2$ 4e2	d 3  ,�O    ��� 8ARPqS�Q��A��B���4p�K����?�L��3� T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARPqS�Q��A��B���4p��K����;�L��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4p��K����7�L��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4p��K����3�L��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4p��K����/�L��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4p��K����'�L��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4p��K����#�L��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4p��K��]���L��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4p��K��]���L��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4���K��]���L��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4���K��]���L��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4���K��]���L��3�T0 k� �����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4���K��]���L��3�T0 k� �����e2$ 4e2	d 3 ��O    ��� 8ARPqS�Q��A��B���4���K��]���L��3�T0 k� �����e2$ 4e2	d 3	 ��O    ��� 8ARPqS�Q��A��B���4���K��]���L��3�T0 k� �����e2$ 4e2	d 3	 ��O    ��� 8ARPqS�Q��A��B���4���K��]���L�3�T0 k� �����e2$ 4e2	d 3
 ��O    ��� 8ARPqS�Q��A��B���4���K��]����L�3�T0 k� ����e2$ 4e2	d 3
 ��O    ��� 8ARPqS�Q��A��B���4���K��]����L{�3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���K��]����L{�3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���C@�]���L{�3�T0 k� ���e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���C@�]���Lw�3�T0 k� ���e2$ 4e2	d 3 ��O   ��� 8ARLqS�Q��A��B���4���C@�]���Lw�3�T0 k� ���e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���C@�]���K�s�3�T0 k� ߁��e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���C@�]���K�s�3�T0 k� ۀ�߀e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���E0�]���K�o�3�T0 k� �ۀ�߀e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���E0�]��߼K�o�3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���E0�]��߼K�o�3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���E0�]��۽K�k�3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���E0�]��׽C�k�3�T0 k� ��~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4���E �]��ӾC�g�3�T0 k� ��~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4��E �]��ӾC�g�3�T0 k� ��}��}e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4��E �]��ϾC�c�3�T0 k� ��}��}e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4��E �]��˿C�c�3�T0 k� ��}��}e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4��E �]��ǿE�_�3�T0 k� ��~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4��B��]��ǿE�_�3�T0 k� ܿ~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4��B��]����E�[�3�T0 k� ܿ~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4��B��]�߿�E�W�3�T0 k� ܻ~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4��B��]�߿�E�S�3�T0 k� ܻ~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4��B��]�߻�E�S�3�T0 k� ܷ~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4��B��]�?��E�O�3�T0 k� �~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4�#�B��]�?��E�K�3�T0 k� �~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4�#�B�#�]�?��E�G�3�T0 k� �~��~e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4�'�B�'�]�?��E�C�3�T0 k� ���e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4�+�B�'�]�?��C�?�3�T0 k� ���e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4�+�C +�\��/��C�;�3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARLqS�Q��A��B���4�/�C /�\��/��C�7�3�T0 k� ����e2$ 4e2	d 3
 ��O    ��� 8ARLqS�Q��A��B���4�3�C /�\��/��C�3�3�T0 k� ����e2$ 4e2	d 3
 ��O    ��� 8ARLqS�Q��A��B���4�3�C 3�\��/��C�/�3�T0 k� ����e2$ 4e2	d 3	 ��O    ��� 8ARLqS�Q��A��B���4�7�C 7�\��/��I�+�3�T0 k� ����e2$ 4e2	d 3	 ��O    ��� 8ARHqS�Q��A��B���4�;�C ;�\�����I�'�3�T0 k� ���e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4q;�C ;�\�����I�#�3�T0 k� ���e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4q?�C ?�\�����I�#�3�T0 k� �����e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4q?�C C�\�����I��3�T0 k� �����e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4qC�C G�\�����I��3�T0 k� �����e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4qG�C K�\�����I��3�T0 k� ܏����e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4qG�CO�\�����I��3�T0 k� ܋����e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4�K�CS�\�����I��3�T0 k� ܋����e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4�O�CW�\����I��3�T0 k� ܇����e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4�O�C[�\����I��3�T0 k� ܇����e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4�S�C_�\����I��3�T0 k� �����e2$ 4e2	d 3 ��O   ��� 8ARHqS�Q��A��B���4�W�Cc�\����I��3�T0 k� ����e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4�W�Ck�\����I��3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�[�Co�\�����I��3�T0 k� {���e2$ 4e2	d 3  ,�O    ��� 8ARHqS�Q��A��B���4�_�Cs�\�����I��3�T0 k� w��{�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�c�Cw�\�����I��3�T0 k� �w��{�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�g�C{�\�����I��3�T0 k� �s��w�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4qg�C ��\�����I��3�T0 k� �s��w�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4qk�C ��\��߻�I��3�T0 k� �o��s�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4qo�C ��\��߻�I��3�T0 k� �k��o�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4qs�C ��\��߿�I��3�T0 k� �k��o�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4qs�C ��\�����I��3�T0 k� �g��k�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4aw�I0��\�����I��3�T0 k� �g��k�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4aw�I0��\�����I��3�T0 k� �c��g�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4a{�I0��\�����AQ�3�T0 k� �_��c�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4a{�I0��\�����AQ�3�T0 k� �_��c�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4a�I0��\�����AQ�3�T0 k� �[��_�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4a�I@��\�����AQ�3�T0 k� �W��[�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�41�I@��\�����AQ�3�T0 k� �W��[�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�41�I@��\�����AQ�3�T0 k� �S��W�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���41��I@��\�����AQ�3�T0 k� �S��W�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���41��I@��\�����AQ�3�T0 k� �O��S�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���41��K�î\�����AQ�3�T0 k� �K��O�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4a��K�í\����AQ�3�T0 k� �K��O�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4a��K�Ǭ\����AQ�3�T0 k� �G��K�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4a��K�˫\���AQ�3�T0 k� �G��K�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4a��K�˪\���AQ�3�T0 k� �C��G�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4a�K�ϩ���AQ�3�T0 k� �?��C�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4a�K�ϩ���AQ�3�T0 k� �?��C�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4a�K�Ϩ���AQ�3�T0 k� �;��?�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B���4Q�K�ϧ���AQ�3�T0 k� 7��;�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4Q{�K�ϧ�p�AQ�3�T0 k� 7��;�e2$ 4e2	d 3 ��O    ��� 8ARHqS�Q��A��B��"�4Q{�K�ϧ�p�AQ�3�T0 k� 3��7�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B��"�4Q{�K�ϧ�p�L�3�T0 k� 3��7�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B��"�4Qw�K�Ϧ�p�L�3�T0 k� /��3�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B��"�4�w�K�ϥ�p�L�3�T0 k� �+��/�e2$ 4e2	d 3  .�O    ��� 8ARHqS�Q��A��B��"�4�s�K�ӥ�p�L�3�T0 k� �+��/�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B��"�4�o�K�Ӥ,�p�L�3�T0 k� �'��+�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B��"�4�o�K�ӣ,�p�L�3�T0 k� �'��+�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B��"�4�k�K�ע,���L�3�T0 k� �#��'�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B��"�4�g�K�ע,���L�3�T0 k� ��#�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B��"�4�c�K�ס,��#�L�3�T0 k� ��#�e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�_�K�נ,��#�L�3�T0 k� ���e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�[�K�۟,��'�L�3�T0 k� ���e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�W�K�۟,��+�L�3�T0 k� ���e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�S�K�۞,��+�L�3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�S�K�ߝ��/�L�3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�S�K�ߝ��3�L!�3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�S�K�ߜ��3�L!�3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�O�K�ߜ��7�L!�3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�O�K����;�L!�3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�O�K����;�L!�3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�O�K����?�L!�3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�O�K����?�L!�3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�K�K����C�L!�3�T0 k� �����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4K�K��\��G�L!�3�T0 k� ������e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4K�K��\��G�L!�3�T0 k� ������e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4K�K��\��K�L!�3�T0 k� ������e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4K�K��\��K�L!�3�T0 k� ������e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4K�K��\��O�L ��3�T0 k� �����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4K�K��\��O�L ��3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4K�K��\��S�L ��3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4K�K��\��S�L ��3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4G�K��\��W�L ��3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4G�K��\��W�L ��3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4C�K��\��[�L ��3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4C�K��\��[�L ��3�T0 k� ����e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4?�K��\��_�L ��3�T0 k� �߈��e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4?�K��\��_�L ��3�T0 k� �߈��e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4;�K��\��c�L ��3�T0 k� �߈��e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���47�K��\��c�L �3�T0 k� �ۉ�߉e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���47�K��\��g�L �3�T0 k� �ۉ�߉e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���43�K��\��g�L �3�T0 k� �׉�ۉe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���43�K���\��g�L �3�T0 k� �׊�ۊe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4/�K���\��k�L �3�T0 k� �׊�ۊe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4/�K���\��k�L �3�T0 k� �ӊ�׊e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4+�K���\��o�L �3�T0 k� �Ӌ�׋e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4+�K���\��o�L �3�T0 k� �Ӌ�׋e2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4+�K���\��o�L �3�T0 k� �ϋ�Ӌe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4+�K���\��s�L �3�T0 k� �ό�ӌe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4'�K���\�ps�L �3�T0 k� �ˌ�όe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4'�K���\�pw�L �3�T0 k� �ˌ�όe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�'�K���\�pw�L �3�T0 k� �ˍ�ύe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�'�K���\�pw�L �3�T0 k� �Ǎ�ˍe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�#�E ��\�p{�L �3�T0 k� �Ǎ�ˍe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�#�E ��\�p{�L �3�T0 k� �Î�ǎe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�#�E ��\���L �3�T0 k� �Î�ǎe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�#�E ��\���L �3�T0 k� �Î�ǎe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4�#�E ��\���L�3�T0 k� ����Ïe2$ 4e2	d 3  ��O    ��� 8ARHqS�Q��A��B���4��E�\�Ѓ�L�3�T0 k� ����Ïe2$ 4e2	d 3  ��O    ��� 8E�X&����g�B��T���4��B�x;���DMB��s���T0 k� �x�|e2$ 4e2	d 3  ��    � 4 �E�h#����w�B��U���4�/�BЌ;����TMB�r���T0 k� �h�le2$ 4e2	d 3  �     � 4 �F�p"�����B��U��4�7�B��:����\LB�r���T0 k� �`
�d
e2$ 4e2	d 3  ��    � 3 �F�x!����B��V��4�C�B��:���dLB�r���T0 k� �\�`e2$ 4e2	d 3  ��    � 2 �F�| ����B��V��4�K�B��:���hLB�$r���T0 k� �T�Xe2$ 4e2	d 3  ��    � 1 �F���õ�B��V��4�S�B��:���pKB�,r���T0 k� �L �P e2$ 4e2	d 3 ��    � 0 �F���˵�B��W�$�4�[�B��:���xKB�4r���T0 k� �G��K�e2$ 4e2	d 3 ��    � / �F���ӵ���B�W�,�4�c�B��9��рJB�<r��T0 k� �?��C�e2$ 4e2	d 3 ��    � . �F���۵���B�W�4�4�k�B��9�'�шJB�Dr��T0 k� �7��;�e2$ 4e2	d 3 ��    � - �F�������B�W�<�4�s�B��9�/�ѐIB�Lr��T0 k� �/��3�e2$ 4e2	d 3 ��    � + �F�������B�X�D�4��E�9�3�єIB�Tr��T0 k� �'��+�e2$ 4e2	d 3 ��    � ) �F�������B�(X�L�4���E�9�;��HB�\r��T0 k� ���#�e2$ 4e2	d 3 ��   � ' �F��������B�0X�T�4���E�8�C��HB�dr��T0 k� ����e2$ 4e2	d 3 ��    � % �Fø�����B�8X�\�4���E 8�K��GB�hr��T0 k� ����e2$ 4e2	d 3 ��    � # �F�������B�@Y�d�4���E8�O��FB�pr��T0 k� ����e2$ 4e2	d 3  ��    � ! �F�������B�HY�l�4���E8�W��FB�xr��T0 k� ����e2$ 4e2	d 3  ��    �  �F�������B�PY�t�4���E8�_���EB��r��T0 k� ������e2$ 4e2	d 3  ��    �  �F���#����B�XY�|�4���E$7�c���DB��r��T0 k� ������e2$ 4e2	d 3  ��    �  �F���+���B�dZބ�4�ÎE07�k���DB��r��T0 k� ������e2$ 4e2	d 3  ��    �  �F���3���B�lZތ�4�ˎE87�s���CB��r��T0 k� ������e2$ 4e2	d 3  ��    �  �F���;���B�tZޔ�4�ӏE�D7�w���BB��r��T0 k� ������e2$ 4e2	d 3  ��    �  �F���K��+�B΄[ޤ�4��E�X7�����AE��r��T0 k� ������e2$ 4e2	d 3  ��    �  �F���O��3�BΌ[ެ�4�E�`7A����@E��r��T0 k� ������e2$ 4e2	d 3  ��    �  �F���W��;�BΔ[޴�4�E�h6A����?E��r��T0 k� ������e2$ 4e2	d 3  ��    �  �F���_��C�BΜ[޼�4��E�t6A���?E��r��T0 k� ������e2$ 4e2	d 3  ��    � 	 �F���g��K�BΨ[���4�E�|6A���>E��r��T0 k� ������e2$ 4e2	d 3  ��    �  �F���k��S�Bް\���4�E��6A���=E��r��T0 k� ������e2$ 4e2	d 3  ��   �  �F��
�s��[�B޸\���4�E��7A���<E��r��T0 k� ������e2$ 4e2	d 3  ��    �   �F��
�{��c�B��\���4�E��7A��� <E��q��T0 k� ������e2$ 4e2	d 3  ��    ��� �F��	����g�B��\���4'�DѤ7A���(;E��q��T0 k� ������e2$ 4e2	d 3  ��    ��� �F��	����o�B��\���4/�DѬ7A���0:E��q��T0 k� ������e2$ 4e2	d 3  ��    ��� �F������w�B��]���47�DѸ7A���89E��q��T0 k� ������e2$ 4e2	d 3  ��    ��� �F�����Ã�B��]� �4�K�D��8AǪ�D7E�q��T0 k� �w��{�e2$ 4e2	d 3  ��    ��� �E#����Ë�B��]�4�S�E��8Q˫L7E�q��T0 k� �o��s�e2$ 4e2	d 3  ��    ��� �E#����Ï�B��]�4�[�E��9QϬT6E�q��T0 k� �g��k�e2$ 4e2	d 3  ��    ��� �E#����Ï�B�^�4�c�E��9Q׭\5E�$q��T0 k� �_��c�e2$ 4e2	d 3  ��    ��� �E#����Ï�B�^ �4�k�E��9Qۮ`4E�,q��T0 k� �W��[�e2$ 4e2	d 3  ��    ��� �E����Ó�B� ^�0�4�{�E�:���p2E�<p��T0 k� �K��O�e2$ 4e2	d 3  ��    ��� �E����×�B�(^�8�4���E�;���x1E�Dp3��T0 k� �C��G�e2$ 4e2	d 3  ��    ��� �E����Ô B�0_�@�4���E�;���|0B�Hp3��T0 k� �;��?�e2$ 4e2	d 3  ��    ��� �E����Ӕ E�8_�H�4��E� <����/B�Po3��T0 k� �3��7�e2$ 4e2	d 3  ��    ��� �E����ӔE�@_�P�4��E�(<�����/B�Xo3��T0 k� �/��3�e2$ 4e2	d 3  ��   ��� �E����ӘE�P_�`�4��Er<=�����-B�hnc��T0 k� �~�#~e2$ 4e2	d 3  ��    ��� �E� b��ӘE�\_�h�4��ErD>����,E�pnc��T0 k� �{�{e2$ 4e2	d 3  )�    ��� �E�� b���E�d_�p�4��ErP?����+E�xnc��T0 k� 2{�{e2$ 4e2	d 3  ��    ��� �E�� b���E�l`�x�4˖ErX?����*E��mc��T0 k� 2|�|e2$ 4e2	d 3  ��   ��� �E�  b���E�|`߈�4ۗErhA����(E��lc��T0 k� 1�~��~e2$ 4e2	d 3  ��    ��� �E���E��`ߐ�4�ErpB��r�'E��lc��T0 k� 1�~��~e2$ 4e2	d 3  ��    ��� �E���E��`ߘ�4	�ErxC��r�&E��kc��T0 k� ����e2$ 4e2	d 3  ��    ��� �E�	��E��`ߠ�4	�Er�D��r�%E��kc��T0 k� ����e2$ 4e2	d 3  ��    ��� �E�
��E��aߨ�4	��Er�E�#�r�#E��jc��T0 k� �߁��e2$ 4e2	d 3  ��    ��� �E�'��E��a߬�4	�Er�F�'�r�"E��jc��T0 k� �ہ�߁e2$ 4e2	d 3  ��    ��� �E��3��E��aߴ�4	�Er�G�'�r�!E��ic��T0 k� �ӂ�ׂe2$ 4e2	d 3  ��    ��� �E��K��E��a�� �4	�Eb�J�/�r�E��hc��T0 k� �Ǆ�˄e2$ 4e2	d 3  ��    ��� �Et�W��E��a�� �4�Eb�K�/�r�E��gc��T0 k� ����Åe2$ 4e2	d 3  ��    ��� �Et�c��E��a����4'�Eb�L�3���E��fc��T0 k� ������e2$ 4e2	d 3  ��    ��� �Et�o��E��`����4/�Eb�N�3�� E��fc��T0 k� ������e2$ 4e2	d 3  ��    ��� �Et�{��|B��`����47�Eb�O�3��E��ec��T0 k� ������e2$ 4e2	d 3  ��    ��� �Et����xB��`����4;�Eb�P�7��E��dc��T0 k� ������e2$ 4e2	d 3  ��    ��� �Et ����p	B��`����4�K�Eb�S�7��E��bc��T0 k� ������e2$ 4e2	d 3  ��    ��� �D�$����l	B�`���4�S�Eb�S�7��CC bc��T0 k� ������e2$ 4e2	d 3  ��    ��� �D�$����h	B�_���4�[�Eb�S�7��$CCac��T0 k� ������e2$ 4e2	d 3  ��    ��� �D�$���d
B�_���4�c�Eb�S�7��(CCac��T0 k� ������e2$ 4e2	d 3  ��    ��� �D�( ���d
B�(^�#��4�s�ER�T�7��(CC `c��T0 k� �s��w�e2$ 4e2	d 3  ��    ��� ~Et,"���d
B�0^�+��4�{�ER�T�7��(CC(`c��T0 k� �o��s�e2$ 4e2	d 3  ��    ��� |Et,$���d	B�8^�/��4���ER�U�7��(CC0`c��T0 k� �g��k�e2$ 4e2	d 3  ��    ��� zEt,&���h	B�@]�7��4r��ER�U�3��(CC8_c��T0 k� �_��c�e2$ 4e2	d 3  ��    ��� xEt0(���hC L]�?��4r��ER�U�3��(CC@^c��T0 k� �[��_�e2$ 4e2	d 3  ��    ��� vEt4,��hC \\�O��4r��ER�V�/��(CCL]c��T0 k� �K��O�e2$ 4e2	d 3  ��    ��� tEt4.��ChC d\�W��4r��C��V�/��(
CCT]c��T0 k� �G��K�e2$ 4e2	d 3  ��    ��� rEt40��ChC l[�_��4r��C��W�+��(CS\\c��T0 k� �?��C�e2$ 4e2	d 3  ��    ��� pEt82�+�ChE�t[ c��4r��C��W�+��(CSd[c��T0 k� �7��;�e2$ 4e2	d 3  ��    ��� nEd84 3�ChE�|Z k��4rÒC��W�'��(CShZc��T0 k� �3��7�e2$ 4e2	d 3  ��    ��� lEd86 ;�ChE��Z s��4r˒C��W2'��(CSpYc��T0 k� �+��/�e2$ 4e2	d 3  ��    ��� jEd8; K�ChE��Y ���4rےC��X2��$CS|Wc��T0 k� ���#�e2$ 4e2	d 3  ��    ��� hEd<= W�ChE��X ���4r�C��X2��$CS�Vc��T0 k� ����e2$ 4e2	d 3  ��    ��� fEd<?S�ChE��X����4r�C��Y2��$CS�Uc��T0 k� ����e2$ 4e2	d 3  ��    ��� dEd<BO�ChE��W����4b�C��Y2��$ CS�Tc��T0 k� ����e2$ 4e2	d 3  ��    ��� bEd<DO��hE��V����4b��C��YR��'�CS�Sc��T0 k� ����e2$ 4e2	d 3  ��O    ��� `Ed8FO��hE��V����4b��C��YR��'�CS�Rc��T0 k� �����e2$ 4e2	d 3  ��O    ��� ^Ed8K�K��dE��U����4c�C��ZR��'�Cc�Pc��T0 k� ����e2$ 4e2	d 3  ��O    ��� \Ed8M�K��dE��T����4c�C��ZR��'�Cc�Nc��T0 k� ����e2$ 4e2	d 3  ��O    ��� ZEd8O�G��`E��S����4c�C��[R��#�Cc�Mc��T0 k� ����e2$ 4e2	d 3  ��O    ��� XET8R�G��`E��R����4c�C��[Q���#�Cc�Lc��T0 k� �ߞ��e2$ 4e2	d 3  ��O    ��� VET4T�G��\E��Q����4c�C��[����#�Cc�Jc��T0 k� �מ�۞e2$ 4e2	d 3  ��O    ��� TET4V�G��\E��P����4c�C��[����#�E��I3��T0 k� �ϟ�ӟe2$ 4e2	d 3  ��O    ��� RET0X�C��XE��O����4c#�C��\����#�E��H3��T0 k� �ˠ�Ϡe2$ 4e2	d 3  ��O    ��� PET0Z�C��TE�N����4S'�C��\����#�E��F3��T0 k� �à�Ǡe2$ 4e2	d 3  ��O    ��� NET,\�C��PE�M����4S+�C��\����#�E��E3��T0 k� ����áe2$ 4e2	d 3  ��O    ��� LET,^�C��PE�L����4S/�C��\����#�E��C3��T0 k� ������e2$ 4e2	d 3  ��O    ��� JET(`dC��LE�K����4S3�D�\���#�E��B3��T0 k� ������e2$ 4e2	d 3  ��O    ��� HC�$dd?��DE�(I���4�7�D�]���#�E��?3��T0 k� ������e2$ 4e2	d 3  ��O    ��� FC� fd?��@E�,G���4�;�D�]���#�E��=3��T0 k� ������e2$ 4e2	d 3  ��O    ��� DC�hd;��<E�0F���4�;�D�]1��#�E��<3��T0 k� ������e2$ 4e2	d 3  ��O    ��� BC�jd;��8E�8EA��4�?�D�^1��#�E��:3��T0 k� ������e2$ 4e2	d 3  ��O    ��� @C�lT7��4E�<DA��4�?�D�^1��'�E��93��T0 k� ������e2$ 4e2	d 3  ��O    ��� >C�nT7��0E�@BA#��4�?�D�^1��'�E��73��T0 k� ������e2$ 4e2	d 3  ��O    ��� <C�oT3��,E�HAA+��4�?�D�^1���'�E� 53��T0 k� �����e2$ 4e2	d 3  ��O    ��� :C�qT3��$E�L@A/��4�C�D�^1���+�E�43��T0 k� �w��{�e2$ 4e2	d 3  ��O    ��� 9C� sT/�� E�P>A7��4�C�D�_1���+�E�23��T0 k� �s��w�e2$ 4e2	d 3  ��O    ��� 8C��uT+��E�T=A;��4�C�D�_1���+�E�03��T0 k� �k��o�e2$ 4e2	d 3  �O    ��� 8AS�vT'�SE�X<A?��4�C�D�_!���/�E�/3��T0 k� �g��k�e2$ 4e2	d 3  �O    ��� 8AS�xT'�SE�\:AG��4�?�D|_!���/�E�-3��T0 k� �_��c�e2$ 4e2	d 3  ��O    ��� 8AS�zT#�SE�`9AK��4�?�Dx_!��/�E�+3��T0 k� �[��_�e2$ 4e2	d 3  ��O    ��� 8AS�{T�SE�d8AO�"�4�?�Dp`!s��3�E�)3��T0 k� �S��W�e2$ 4e2	d 3  ��O    ��� 8AS�}T�SE�h6AW�"�4�?�ERh`!k��3�E�(3��T0 k� �K��O�e2$ 4e2	d 3  ��O    ��� 8AS�~T�R�E�l5A[�"�4�;�ER``!_��7�E�&3��T0 k� �G��K�e2$ 4e2	d 3  ��O    ��� 8AS�T�R�Ap4A_�"�4�;�ER\`!W�s7�E�$3��T0 k� �?��C�e2$ 4e2	d 3  ��O    ��� 8AS�T�R�At3Ac�"�4�;�ERT`!O�s7�E�"3��T0 k� �;��?�e2$ 4e2	d 3  ��O    ��� 8AS�T�R�Ax2Ak�"�4�7�ERL`!C�s;�E� 3��T0 k� �3��7�e2$ 4e2	d 3  ��O    ��� 8AS�T�R�A|0Ao�"�4�3�EBDa!;�s;�E�3��T0 k� �/��3�e2$ 4e2	d 3  ��O    ��� 8AS�T�R�A|/As�"�4�3�EB<a!3�s?�E�3��T0 k� �'��+�e2$ 4e2	d 3  ��O    ��� 8AS�T�R�A�.Aw�"�4�/�EB4a!+�s?�E�3��T0 k� �#��'�e2$ 4e2	d 3  ��O    ��� 8AS�T�R�A�-A{�"�4�+�EB,a!�s?�E�3��T0 k� ����e2$ 4e2	d 3  ��O    ��� 8AS�T�R�A�,A�"�4+�EB$a!�cC�E�3��T0 k� ����e2$ 4e2	d 3  ��O   ��� 8AS�T�R�A�+A���4'�EBa!�cC�E�3��T0 k� ����e2$ 4e2	d 3  ��O    ��� 8AS�T�R�A�*A���4#�EB`!�cC�C�3��T0 k� ����e2$ 4e2	d 3  ��O    ��� 8AS�S��R�A�)A���4�EB` ��cC�C�3��T0 k� ����e2$ 4e2	d 3  ��O    ��� 8AS�S��R�A�(A���4�EB` ��cG�C�3��T0 k� �����e2$ 4e2	d 3  ��O    ��� 8AS�S��R�A�'A���4�EB ` ��cG�C�3��T0 k� ������e2$ 4e2	d 3  ��O    ��� 8AS�S��R�A�&A���4�EA�_ ��cG�C�3��T0 k� �����e2$ 4e2	d 3  ��O    ��� 8AS�S��R�A�%A���4�E1�_ ��cG�C�3��T0 k� ����e2$ 4e2	d 3  ��O    ��� 8AS�S��R�A�$A���4�E1�_ ��cG�C�3��T0 k� ����e2$ 4e2	d 3  ��O    ��� 8AS�S�R�A�#A���4�E1�^ ��cG�C�3��T0 k� �ߺ��e2$ 4e2	d 3  ��O   ��� 8ASxS�R�A�"A���4��E1�^ ��SG�C� 3��T0 k� �ۻ�߻e2$ 4e2	d 3  ��O    ��� 8AStS�R�A�!A���4��E1�] ��SG�C��3��T0 k� �ӻ�׻e2$ 4e2	d 3  ��O    ��� 8ASpS�R�A� A��"�4��E1�\ ��SC�C�� 3��T0 k� �ϼ�Ӽe2$ 4e2	d 3  ��O    ��� 8ASlS�R�A�A��"�4�E1�\P��SC�C�� 3��T0 k� �ǽ�˽e2$ 4e2	d 3  ��O    ��� 8ASdS�R�A�A��"�4�E1�[P��SC�C�� 3��T0 k� �ý�ǽe2$ 4e2	d 3  ��O    ��� 8AS`�S�R�A�A��"�4�E1�ZP��SC�C�� 3��T0 k� ����þe2$ 4e2	d 3  ��O    ��� 8AS\S�R�A�A��"�4߂E1�YP��S?�C��!3��T0 k� ������e2$ 4e2	d 3  ��O    ��� 8ASXS�R�A�A��"�4ׂCA�XP���?�C��!3��T0 k� ������e2$ 4e2	d 3  ��O    ��� 8ASTS�R�A�A��"�4ӃCA�XP���?�C��!3��T0 k� ������e2$ 4e2	d 3  ��O    ��� 8ASPS�R�A�A��"�4˃CA�WP���;�C��"3��T0 k� ������e2$ 4e2	d 3  ��O    ��� 8ASL~S߲R�A�A��"�4ÃCA�VP��;�C��"3��T0 k� ������e2$ 4e2	d 3  ��O    ��� 8ASH~S߱R�A�A��"�4��CA�U�o��7�D�"3��T0 k� ������e2$ 4e2	d 3  ��O    ��� 8ASD~S۱R�A�A��"�4ⷃKфT�c��3�D�"3��T0 k� ������e2$ 4e2	d 3  ��O    ��� 8AS@~S۱R�A�A���4⯄KрS�S��3�D�#3��T0 k� ������e2$ 4e2	d 3  ��O    ��� 8AS<}S۰R�A�A���4⧄K�xS�G�/�D�#3��T0 k� ������e2$ 4e2	d 3  ��O   ��� 8AS8}SװR�A�A���4⣄K�tR�7�+�D�#3��T0 k� ������e2$ 4e2	d 3  ��O    ��� 8AS4}SװR�A�A���4⛄K�lQ�+�+�EC�#3��T0 k� �����e2$ 4e2	d 3  ��O    ��� 8AS0}SӯR�A�A���4ⓄK�hP��'�EC�#3��T0 k� �w��{�e2$ 4e2	d 3  ��O    ��� 8AS,|SӯR|A�A���4⋅K�`P��'�EC�#3��T0 k� �s��w�e2$ 4e2	d 3  ��O    ��� 8AS(|SӯR|A�A���4⃅K�\O��#�EC�#3��T0 k� �k��o�e2$ 4e2	d 3  ��O    ��� 8AS$|SϯRxA�A���4�{�K�XN���#�EC�#3��T0 k� �g��k�e2$ 4e2	d 3  ��O    ��� 8AS |SϮRtA�A���4�s�K�PM����EC�#3��T0 k� �_��c�e2$ 4e2	d 3  ��O    ��� 8AS|SϮRtA�A���4�k�K�LM����EC�#3��T0 k� �[��_�e2$ 4e2	d 3  ��O    ��� 8AS{SˮRpA�A���4�c�K�HL����C��"3��T0 k� �W��[�e2$ 4e2	d 3  ��O    ��� 8AS{S˭RlA�A���4�[�K�@K����C��"3��T0 k� �O��S�e2$ 4e2	d 3  ��O    ��� 8AS{S˭RlA�A���4�S�K�<K߻��C��"3��T0 k� �K��O�e2$ 4e2	d 3  ��O    ��� 8AS{SǭRhA�A���4�G�K�8J߯��C�x!3��T0 k� �C��G�e2$ 4e2	d 3  ��O    ��� 8AS{SǭRhA�A���4�?�K�4Iߣ��C�p!3��T0 k� �?��C�e2$ 4e2	d 3  ��O    ��� 8AS{SǬRdA�A���4�7�K�,Iߛ�#�C�l!3��T0 k� �;��?�e2$ 4e2	d 3  ��O    ��� 8ASzSìR`A�B��4�/�K�(Hߏ�#�C�d 3��T0 k� �3��7�e2$ 4e2	d 3  ��O    ��� 8ASzSìR`A�B��4�'�K�$H߃�#�C�\ 3��T0 k� �/��3�e2$ 4e2	d 3  ��O    ��� 8AS zSìR\A�B��4��K� G�{�#�C�X3��T0 k� �/��3�e2$ 4e2	d 3  ��H    ��� 8AR�zSëR\A�B��4��K�F�o�#�C�P3��T0 k� �+��/�e2$ 4e2	d 3  ��H    ��� 8AR�zS��RXA�
B��4��K�F�g�#�C�H3��T0 k� �#��'�e2$ 4e2	d 3  ��H    ��� 8AR�zS��RXA�
B��4��K�E�[�#�C�D3��T0 k� ����e2$ 4e2	d 3  ��H    ��� 8AR�yS��RTA�	B��4��K�E�S�#�C�<3��T0 k� ����e2$ 4e2	d 3  ��H    ��� 8AR�yS��RTA�	B��4�K�D�G�"��C�43��T0 k� ����e2$ 4e2	d 3  ��H    ��� 8AR�yS��RPA�B��4�K�Do?�"��C�,3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�yS��RPA�B��4�K� Co3�"��C�(3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�yS��RLA�B��4ۈK��Bo+�"��C� 3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�yS��RLA�B��4QψK��Bo#�"��C�3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�yS��RHA�B��4QǈK��Ao�"��C�3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�xS��RHA B��4Q��K��A_�"��C�3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8AR�xS��RDA B#��4Q��K��@_�"��C�3��T0 k� ������e2$ 4e2	d 3  ��H    ��� 8                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��n� ]�(�(� 
� �� qgo   W    � �-     qgo �-                      n <          �     ���   
	          ����    )     � �2�    ���� �2�           	        #               ��     ���   0&         ��'�           j�O    ��'� j��      ��   
            �� :         +�     ���   8	
         ���          h}n    ��� h}n                     
   �$          p     ���   @

          ����   $ $      . ��|    ���� ���                    	 	����          P@     ���   8
4

          >�  ��       B��r     >���r                             ���\              �  ���     

 0            ��<�  > >      V G�     ��N� HCJ    ���b            �� 8�        �P�     ��@    	
          ��;� Q Q      j @LF    ���� ?�0    �n�               �� 8          Gb     ��@ 
0
&
 
          �� #   |	     ~�:��    �� #�:�      ��           �� 8         r     ��H   8

	         ����  M M     �  Vk    ���� �:    ���             V�� 8         	 ���     ��@  8


         ���� � � 
	   � 8o�    ��}� 8�x     ��[            
	�� 8         
 ��    ��`  03 	           :� ��
	      � �s�     :� �s�                              ���]               ��@   

 0
 
                 ��      �                                                                           �                               ��        ���          ��                                                                 �                         ���  ��        ���s�  ����G���Ԭ  ����M                  x                j  �   �   �                         ��    ��        ���      ��  ��           "                                                �                          � � j h �� G @�:   8 �������   
 	             
   �   � �� ����       7� `m@ 8� @n  :d n� ��  s� �D v  �d v@ ? @k� ?� l  H 0u� Hd u� H� v ���X � J v  J$ v@ 
�\ V  $ `r@ � s   s  
�| W� 
�| W� 
�| W� �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� �R� � }`���� ����� � 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���� 8 ������  ������  
�fD
��L���"����D" � j  "  B   J jF�"     
�j � � 
��
��
��"    "D�j  
� `  "  �
� �  �  
� ����  ��     ���  �   ��    ��     � �      ����  ��     ��:          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �O	4	      �� � �  ��        � �T ��        �        ��        �        ��        �    ��    ��������        ��                         ���   
� ��                                    �         
        ����           ���� ���%��  �� 8 2                7 Neal Broten ll  k   0:01                                                                        5  3     � �
"� �C
� � �c� � � c� � �k� � � k� � �	kj � �kp � � 	kt � �
cV � � c\ � �K �K" �C* � C2 fC. � v C6 � �"� � � "� � {"� � {*� � x!� | � "J � � "  |8  "J � x!� | � "J � � "  |8  "J � x!� | � "E �8  "E �8  "E �8  "E �8  "J � � $"  |8  "J �8  "J �8  "E � � ("& � �)". |@  "K � �+". |@  "K �8  "E �8  "E � �/!� | � 0"J �,  "  | � 2"@ | � 3"P �  4"& |0  "* |2 )�|L 7*Pd\  *HdX  *HjX  *KyX  *Hy �<*<g=*2w#>*:g3  *Pw                                                                                                                                                                                                                         d� P         �    @ 
         �     ^ P E _  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    �`~�l� ��������������������������������������������������������   �4, =�
 * �
@��@�
�@؂�O�������                                                                                                                                                                                                                                                                                                                               ��
                                                                                                                                                                                                                                                    H    4    ��   :�J      E�  	                           ������������������������������������������������������                                                                                                                               
           �    �    �        �      ��                  
     ��� �� ����� �  ����������������������� ������ ���� �������� ���� �� �������������� ��������� ����� ���� �� ����������������������� ��������������� ������������������� ����������������������������������������� ������������������� ���             x                    6    .    ��  !N�J      he  	                           ������������������������������������������������������                                                                                                                                    �  �  �     �                ��                	   	 	  ���������������������������������������� ���������������� ���� ������������������������������ ������������������������������ ���������������� � �������������� ����������������� ������� ��� ������ ���   ������ ����� �����������                                                                                                                                                                                                                                                              	                                                           �             


             �  }�         ������������  *���������  +����������������  '�   ������������  'q������������������������������������                         '�                              N�  N�                     ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" < D <                                 � +� �t�                                                                                                                                                                                                                                                                                       )n)n	n  �)�                k            a            a                                                                                                                                                                                                                                                                                                                                                                                                                j          > �  
>�   7  #�  C#�  Fa�  ��� ��:�Y��v�������˖�D��8�������������                ���E :�� 
         �   & AG� �  �   
              �                                                                                                                                                                                                                                                                                                                                        K C    z                     !��                                                                                                                                                                                                                            Y��   �� � Ѱ��      �� 7      ��� �� ����� �  ����������������������� ������ ���� �������� ���� �� �������������� ��������� ����� ���� �� ����������������������� ��������������� ������������������� ����������������������������������������� ������������������� ��� ���������������������������������������� ���������������� ���� ������������������������������ ������������������������������ ���������������� � �������������� ����������������� ������� ��� ������ ���   ������ ����� �����������             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    B   !   @     ��                       7     �   ���������J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p����      � �N     `d  �@���6 ��  �@���6 �$ ^$ �r@  �@  �r@      4 
�V   �     ����� ��   ����� �$ ^$  )   �                       ��  t� �D �� t� �D Q �� � ���� �  �      �  ��   ���� e�����  g���        f ^�         �� L��            ��o���2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                               	                 �  ��� �UU���U              �	���UUU�UUUUUU      	� ��U�UUUUUUUUUUUUUUUUUUU    ��� U^��UUU�UUU^UUUUUUUUUUUU            �   �   ^�  U�  UY�    � 	UU 	��  	�  	�  �^ 	��    �	UY�������UUUUUUU��UU��UU�U�UUUUUUUUUUUUUUUUUUUUUUUUUUUU^UUUYUU^�U^� U� ^�  �  ��  �   �   ��UU ��U �U  �U  ��            U^� UU� UU� UU� ���                    	   �       	   	   	    �UUU�UU���U  	�� �����U�UUU�UUUUUUYUUUYUUUYUUU^UUU^UUUUUUUUUUUU�   �   �   �   �   � �^���U^��            	����UUU�UUU�UUUUUU^            ��  U�  Y�  �  �      �   �   �   	                ���Y���U��Y�^�U��U ��^ 	� 	� UUUU�UUUUUUUU^�U^����� �        UUUUUUUUUUUUUUUUUUUU�������    UUU�UU^�UU�U� Y�  ��          �                               wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  " ! " ""      " ""   "" !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                        "!  "! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                            �� ������}����zvw� w
�  ��  �� 	�� �� ��� ��� ��� ��� �� ɘ�̾ �˰ +�  �                   ��   �    �                            ��  �ɨ �݋������������������������˼�̹�˸�븙� �UU X�U X�U U�U D�T �K ̸ �� �� "�  " ��   �                    �   �   �   T   T   T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ���� ��� ����                            �   O   T     ��                                 � ���� ��   � � �                                                                                                                                                         
   �   �  
�  �  ��  ��� ��� ���ཉ��=  
3  �D  �C  �T  �U  �T  ��  �� 
� �,� ,�  �"             �  �˰ ̻� �ݰ �w� ��� ��� ����������˚�̸���ۛ��ݻ�˽�̹� ��" �3: DDJ 33C 334�CET0�4K� ��� 	�� 
�� �  �/ "�������  �                 �   �           ɪ  ��� ټ� �̰ �̰ ��� ��  ��     �   � � �  ��� ��  �                       �   �                      �������  ���    �                      �    �                    ��                 � ���� ��   � � �                                                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��   "  " "  ��  �              �   � � �  ��� ��  �             "  �"     �                            �    ���  ��                    ��  ��  ���     �     �                                                                                                                                                                                                  �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �   ��/ ""� "!� "�"�!�  ��                    � �������� �              ��  ����� ��                           �   ���         �     �                                                                                                                                                                                         �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   �   �"  ""  !� �� ��  �               �   ������  ��   ����   �       �                                   �    ���  ��                    ��  ��  ���                                                                                                                                                                                                   �� ̽ �� �� w}  �� 
�� ��� ��� ��� ��� ��  �� �� �� 	�� �� 4U 33 �3= ݘ� �۽������ʸ�	˽��� "��                                  ��  ��  �ˀ ��� ͚���ػ��ۻ�̽��˸.���"��� 	��M UJ��ET��UM��D��߈ۛ�ۋ�ٰ ��� ����-�������"��� �           �   ��                     �   �   �  �  "  �         �   �   �   �            �        � ����� ��     �  �  �          �   �  �  �   �               �   �                               � ����ݼ� ����                                                                                 �  �  ��  �                                                                     � 
��	�˽���w��{k��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            �  �  �  ��  �            ��  ��                                �  �� �  �  �   �     "  "  "                       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����            �����                                  �  �˰ ��� �wp ���                       ����     �   �  �  �  ��  �   �                           ��   ��                  �  �  �� � ���    �  �                                 �  	�  ˹ ˹ �̹ ��� ̽� ̽�̽�	�ͺ������J�CT�T UJ� UT� EU� T� J�  ��  ��  ʩ ̰ �  "" "" ""    ��   ��  ��  ��  �w  �p  ��  ��  ��  ̰  Ȱ  ��  ��  ��  ��  "�  0"� 3 � 30�C0 �C  Ƞ  ��  ��  ݻ ��"/""""""/"��� ��� ��             �� ������ ����  �   �  �   �  �     �                                       ��        �        �   �     �       �   �   �   �   �      �                    ��� ���� ��    ��   �  ��  �  �  �         � �������������  �                                                                                                                                        �����̬̽��̽��̽���ת
wz� ��� ��� ˙� �) "+ .# 32� 33� �3> �3> �� � "  " "" "   "/� �  �                            �   ˰  ��  �̰ ��� �̻���ː�۹������̅�̙U�����
�ŀ���̵�̵K�D��"L�"  ""  "" ��.����������     �  ��  �   ��  ��            "   "   "   "   ��   ��  �  �   �    �                            �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                ��  ��  ��� ���                                                                                                                                                                                              ˰ ̻ ̻ �� {�  �� 
�� ��� ��� ������
���	��ܻ̍ݻ���"� 8"  8  �  D�  H�  X�  ��  �   �          "  "     �                        ��  ��� �̺�̻����ۻ�˽��̽��̝ ̙� �30 �EP �U@ �T0 EC0 T3  C:  K�  �"  �"/ ����˽� �"� "" �""� � �� ��      �   �� ��  �"  �                   
 "� ""� ""� "                       �                             ���                         �  ��                    �����                                  �  �˰ ��� �wp ���                                                                                                                                                                   �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                        � ��                  �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                          �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��                  �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                         @  @  @  @  @  @                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""��������������������""""������DDM�D��""""�������MM�M�M""""��������DD�A��""""�������MAA�MA""""��������AA�A""""����������M�MA""""������������M���M���M���"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUQUUQUUUUUUQUUUUUUUU3333DDDDUUUUDEEDDTEUUUU3333DDDDAEAEQQUDTDUUUU3333DDDDQUQUQDUDDUUUU3333DDDDAADAUAUEDUTUUUU3333DDDDADAEAQAUEDUTUUUU3333DDDDUDUQEUQUUQUEUDUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwDGqGq""""wwwwwwqwDqq""""wwwwwwGwGwGwGw""""wwwwwwwGwqGwGwDGw""""wwwwwqwDqqq""""wwwwwwwGwwDGwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD������������������������3333DDDDJ�JDJ�DD�����3333DDDDADAJ�J��J�D����3333DDDDJ�J��DD�����3333DDDDJ�J�DJJDD�J����3333DDDDA�AA�����D�D����3333DDDD���J��J��J��D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=""""��������AA�A    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ADA�LL��L�D����3333DDDD x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(XxLL����������D����3333DDDD w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""����������A������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(""""�������I�I������ �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�""""�������I��D���I������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`�D�M�D���M������3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(MD�M�A�����MD�����3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(�""""�����AMAD������ � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(�""""������������������ � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(�""""�������DAADAI � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(��A�AM�M�DM��M334CDDDD 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5DD����M��DM�����3333DDDD x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x""""wwwwwwDGqGq w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwwGwwDGwwwwwwww + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+ADAH�DJ�H�H�����3333DDDD � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(��H��J�AD�DH�D����3333DDDD � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(�""""�������DD����� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
"� �C
� � �c� � � c� � �k� � � k� � �kj � �kr � � 	kt � �
cV � � c\ � �K �K" �C* � C2 fC. � v C6 � �"� � � "� � {"� � {*� � x!� | � "J � � "  |8  "J � x!� | � "J � � "  |8  "J � x!� | � "E �8  "E �8  "E �8  "E �8  "J � � $"  |8  "J �8  "J �8  "E � � ("& � �)". |@  "K � �+". |@  "K �8  "E �8  "E � �/!� | � 0"J �,  "  | � 2"@ | � 3"P �  4"& |0  "* |2 )�|L 7*Pd\  *HdX  *HjX  *KyX  *Hy �<*<g=*2w#>*:g3  *Pw3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������$��7�O�Q�K��7�U�J�G�T�U� � � � � � � � � �.�+�6�����������������������������������������!��;�[�Y�Y��-�U�[�X�Z�T�G�R�R� � � � � � �.�+�6�����������������������������������������"��8�K�G�R��,�X�U�Z�K�T� � � � � � � � � �.�+�6�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������.�+�6� �� �������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�1�B� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            