GST@�                                                           �e�                                                      8  /                       �������r�	 J�����������H���z���        �h     #    z���                                d8<n    �  ?     b`����  �
fD�
�L���"����D"��   " `  J  jF��    "�j "����
��
��     �j�� 
   ��
  k                                                                               ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������?  0b  5  81                      
     
              �  4    �                  Yn  1          := �����������������������������������������������������������������������������                                �   *       �   @  &   �   �                                                                                 '       )n)n1n  Y1n    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��L���Eo�^O�K�c�Y|8]'� m�P]l@H mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������M��Es�^O�K�c�Y|8]'� m�P]l@H mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��   �������M��Ew�^O�K�c�Y|8]'� m�P]l@H mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������M��B�w�^O�K�g�Y|8]'� m�P]l@H mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������M��B�{�^O�K�g�Y|8]'� m�P]l@H mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������M��B��^O�K�g�Y|8]'� m�P]l@H mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������M��B���^O�K�g�Y|8]'� m�P]l@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������M��B���^O�K�g�Y|8]#� m�P]l@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������M��B���^O�K�k�Y|8]#� m�P]l@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������M��B���^O�K�k�Y|8]#� m�P]l@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���B���^S�K�k�Y|8]#� m�P]h@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���B���^S�K�k�Y|8]#� m�P]h@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���B���^S�K�k�Y|8]#� m�P]h@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���B���^S�K�k�Y|8]#� m�P]h@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���B���S�K�o�Y|8]#� m�P]h@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���B���S�K�o�Y|8]#� m�P]h@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���B���W�K�o�Y|8]#� m�P]h@L mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���B���W�K�o�Y|8]#� m�P]h@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��   �������L���B���W�K�o�Y|8]#� m�P]h@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������A��B���W�K�o�Y|8]#� m�P]h@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������A��B�âW�K�s�Y|8]#� m�P]h@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������A��B�ǡW�K�s�Y|8]#� m�P]h@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������A��B�ϠW�K�s�Y|8]#� m�P]h@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������A��B�ӟW�K�s�Y|8]#� m�P]d@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������A��B�ӟW�K�s�Y|8]#� m�P]d@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������A��B�מ[�K�s�Y|8]#� m�P]d@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������A��B�מ[�K�w�Y|8]#� m�P]d@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ����� n�A��Eם[�K�w�Y|8]#� m�P]d@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ����� n�A��Eۜ._�K�w�Y|8]#� m�P]d@P mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ����� n�A��Eߛ._�K�w�Y|8]#� m�P]d@T mg�c��T0 k� �����&�1D"3Q	2�D 3Q  ��    ����� n�A��Eߛ._�K�w�Y|8]#� m�P]d@T mg�c��T0 k� �����&�1D"3Q	2�D 3Q  ��    ����� n�A��E�._�K�w�Y|8]#� m�P]d@T mg�c��T0 k� �{���&�1D"3Q	2�D 3Q  ��    �������A��E�._�K�w�Y|8]#� m�P]d@T mg�c��T0 k� �{���&�1D"3Q	2�D 3Q  ��    ������#�A��E��.c�K�{�Y|8]#� m�P]d@T mg�c��T0 k� �w��{�&�1D"3Q	2�D 3Q  ��    ������#�A��E��.c�K�{�Y|8]#� m�P]d@T mg�c��T0 k� �w��{�&�1D"3Q	2�D 3Q  ��    ������'�A��E��.c�K�{�Y|8]#� m�P]d@T mg�c��T0 k� �s��w�&�1D"3Q	2�D 3Q  ��    ������'�A��E��.g�K�{�Y|8]#� m�P]d@T mg�c��T0 k� �s��w�&�1D"3Q	2�D 3Q  ��   ������'�A��E��.g�K�{�Y|8]#� m�P]d@T mk�c��T0 k� �o��s�&�1D"3Q	2�D 3Q  ��    ������+�A��E���.g�K�{�Y|8]#� m�P]d@T mk�c��T0 k� �o��s�&�1D"3Q	2�D 3Q  ��    ������+�A��E���.g�K��Y|8]#� m�P]d@T mk�c��T0 k� �k��o�&�1D"3Q	2�D 3Q  ��   ������+�A��E���.g�K��Y|8]#� m�P]d@T mk�c��T0 k� �k��o�&�1D"3Q	2�D 3Q  ��    ������+�A��E}��.g�K��Y|8]#� m�P]`@T mk�c��T0 k� �g��k�&�1D"3Q	2�D 3Q  ��    ������+�A��E}��.g�K��Y|8]#� m�P]`@T mk�c��T0 k� �g��k�&�1D"3Q	2�D 3Q  ��    ������+�A��E}��.g�K��Y|8]#� m�P]`@T mk�c��T0 k� �c��g�&�1D"3Q	2�D 3Q  ��    ������+�A��E}��.k�K��Y|8]#� m�P]`@T mk�c��T0 k� �c��g�&�1D"3Q	2�D 3Q  ��    ������/�A��E~�.k�K��Y|8]#� m�P]`@X mk�c��T0 k� �_��c�&�1D"3Q	2�D 3Q  ��    ������/�A��D��.k�Kރ�Y|8]#� m�P]`@X mk�c��T0 k� �_��c�&�1D"3Q	2�D 3Q  ��    ������/�A��D��.o�Kރ�Y|8]#� m�P]`@X mk�c��T0 k� �[��_�&�1D"3Q	2�D 3Q  ��    ������/�A��D��.o�Kރ�Y|8]#� m�P]`@X mk�c��T0 k� �[��_�&�1D"3Q	2�D 3Q  ��    ������/�A��D��.s�Kރ�Y|8]#� m�P]`@X mk�c��T0 k� �W��[�&�1D"3Q	2�D 3Q  ��    ������3�A��D��.s�CN��Y|8]#� m�P]`@X mk�c��T0 k� �W��[�&�1D"3Q	2�D 3Q  ��    ������3�A��L^�.s�CN��Y|8]#� m�P]`@X mk�c��T0 k� �S��W�&�1D"3Q	2�D 3Q  ��    ������3�A��L^�.w�CN��Y|8]#� m�P]`@X mk�c��T0 k� �S��W�&�1D"3Q	2�D 3Q  ��    ������3�A��L^�.w�CN��Y|8]#� m�P]`@X mk�c��T0 k� �O��S�&�1D"3Q	2�D 3Q  ��    ������3�A��L^�.w�CN��Y|8]#� m�P]`@X mk�c��T0 k� �O��S�&�1D"3Q	2�D 3Q  ��    ������7�A��L^�.{�@���Y|8]� m�P]`@X mk�c��T0 k� �O��S�&�1D"3Q	2�D 3Q  ��    ������7�A��L^�.{�@���Y|8]� m�P]`@X mk�c��T0 k� �K��O�&�1D"3Q	2�D 3Q  ��    ������7�A��L^�.{�@���Y|8]� m�P]`@X mk�c��T0 k� �K��O�&�1D"3Q	2�D 3Q  ��    ������;�A��L^#�.�@���Y|8]� m�P]`@X mk�c��T0 k� �G��K�&�1D"3Q	2�D 3Q  ��    ������;�A��L^#�.�@���Y|8]� m�P]`@X mk�c��T0 k� �G��K�&�1D"3Q	2�D 3Q  ��    ������;�A��L^'�.�E·�Y|8]� m�P]`@X mk�c��T0 k� �C��G�&�1D"3Q	2�D 3Q  ��    ������;�A��Ln+�.��E·�Y|8]� m�P]`@X mk�c��T0 k� �C��G�&�1D"3Q	2�D 3Q  ��    ������?�A��Ln+�.��E·�Y|8]� m�P]`@X mk�c��T0 k� �?��C�&�1D"3Q	2�D 3Q  ��    ������?�A��Ln/�.��E·�Y|8]� m�P]`@X mk�c��T0 k� �?��C�&�1D"3Q	2�D 3Q  ��    ������?�A��Ln/�.��E·�Y|8]� m�P]`@\ mk�c��T0 k� �;��?�&�1D"3Q	2�D 3Q  ��   ������C�A��Ln3�.��E·�Y|8]� m�P]`@\ mk�c��T0 k� �;��?�&�1D"3Q	2�D 3Q  ��    ������C�A��Ln3�.��E·�Y|8]� m�P]`@\ mk�c��T0 k� �7��;�&�1D"3Q	2�D 3Q  ��    ������C�A��Ln7�.��E·�Y|8]� m�P]\@\ mk�c��T0 k� �7��;�&�1D"3Q	2�D 3Q  ��    ������G�A��Ln7�.��E·�Y|8]� m�P]\@\ mk�c��T0 k� �3��7�&�1D"3Q	2�D 3Q  ��    ������G�A��Ln;���E·�Y|8]� m�P]\@\ mk�c��T0 k� �3��7�&�1D"3Q	2�D 3Q  ��    ������G�A��Ln;���E·�Y|8]� m�P]\@\ mk�c��T0 k� �3��7�&�1D"3Q	2�D 3Q  ��    ������G�A��Ln?���E·�Y|8]� m�P]\@\ mk�c��T0 k� �/��3�&�1D"3Q	2�D 3Q  ��    ������K�A��Ln?���A��Y|8]� m�P]\@\ mk�c��T0 k� �/��3�&�1D"3Q	2�D 3Q  ��    ������K�A��LnC���A��Y|8]� m�P]\@\ mk�c��T0 k� �+��/�&�1D"3Q	2�D 3Q  ��    ������K�A��LnC���A��Y|8]� m�P]\@\ mk�c��T0 k� �+��/�&�1D"3Q	2�D 3Q  ��    ������K�A��LnG���A��Y|8]� m�P]\@\ mk�c��T0 k� �'��+�&�1D"3Q	2�D 3Q  ��   ������O�A��LnG���A��Y|8]� m�P]\@\ mk�c��T0 k� �'��+�&�1D"3Q	2�D 3Q  ��    ������O�A��LnG���C���Y|8]� m�P]\@\ mk�c��T0 k� �#��'�&�1D"3Q	2�D 3Q  ��    ������O�A��LnG���C���Y|8]� m�P]\@\ mk�c��T0 k� �#��'�&�1D"3Q	2�D 3Q  ��    ������O�A��LnG���C���Y|8]� m�P]\@\ mk�c��T0 k� ���#�&�1D"3Q	2�D 3Q  ��    ������O�L���LnG���C���Y|8]� m�P]\@\ mk�c��T0 k� ���#�&�1D"3Q	2�D 3Q  ��    ������O�L���LnG���C���Y|8]� m�P]\@\ mk�c��T0 k� ���#�&�1D"3Q	2�D 3Q  ��    ������O�L���LnK���C���Y|8]� m�P]\@\ mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ������O�L���LnK���C���Y|8]� m�P]\@\ mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ������O�L���LnK�^��C���Y|8]� m�P]\@\ mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ������O�L���LnK�^��C���Y|8]� m�P]\@\ mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ������O�L���LnK�^��C���Y|8]� m�P]\@\ mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ������O�L���LnK�^��C��Y|8]� m�P]\@\ mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ������O�L���LnO�^��C��Y|8]� m�P]\@\ mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ������O�L���LnO�C�{�Y|8]� m�P]\@\ mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ������O�M��LnO�C�{�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ������O�M��LnO�C�{�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� nO�M��LnO�C�w�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� nO�M��LnO�C�w�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� nO�M��LnS���C�w�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� nO�M��LnS���C�w�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� nO�M��LnS���C�w�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� nO�M��LnS���C�w�Y|8]� m�P]\@` mk�c��T0 k� �����&�1D"3Q	2�D 3Q  ��    ����� nO�M��LnS���C�s�Y|8]� m�P]\@` mk�c��T0 k� �����&�1D"3Q	2�D 3Q  ��    ����� nO�L���LnS���C�s�Y|8]� m�P]\@` mk�c��T0 k� �����&�1D"3Q	2�D 3Q  ��    ����� nO�L���LnS���C�s�Y|8]� m�P]\@` mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ����� �O�L���LnW���C�s�Y|8]� m�P]\@` mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ����� �O�L���L^W���C�s�Y|8]� m�P]\@` mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ����� �O�L���L^W���C�s�Y|8]� m�P]\@` mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ����� �O�L���L^W���C�s�Y|8]� m�P]\@` mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ����� �O�L���L^W���CNs�Y|8]� m�P]\@` mk�c��T0 k� �����&�1D"3Q	2�D 3Q  ��    ����� �O�L���L^W�.��CNs�Y|8]� m�P]\@` mk�c��T0 k� �����&�1D"3Q	2�D 3Q  ��    ����� �O�L���L^W�.��CNs�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� �O�A��D�[�.��CNs�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� �O�A��D�[�.��CNs�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� �O�A��D�[�.��CNs�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� �O�A��D�[�.��CNs�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ����� �O�A��D�[�.��CNs�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��CNs�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��C^s�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��C^s�Y|8]� m�P]\@` mk�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��C^s�Y|8]� m�P]\@` mk�c��T0 k� �߫��&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��C^s�Y|8]� m�P]\@` mk�c��T0 k� �ߪ��&�1D"3Q	2�D 3Q  ��   �����O�A��D�[�.��C^s�Y|8]� m�P]\@` mk�c��T0 k� �ߪ��&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��C^s�Y|8]� m�P]\@` mk�c��T0 k� �۪�ߪ&�1D"3Q	2�D 3Q  ��   �����O�A��D�[�.��C^s�Y|8]� m�P]\@` mk�c��T0 k� �۪�ߪ&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��C^s�Y|8]� m�P]\@` mk�c��T0 k� �ת�۪&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��@�s�Y|8]� m�P]\@` mk�c��T0 k� �ש�۩&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��@�s�Y|8]� m�P]\@` mk�c��T0 k� �ש�۩&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��@�s�Y|8]� m�P]\@` mk�c��T0 k� �ө�ש&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��@�s�Y|8]� m�P]\@d mk�c��T0 k� �ө�ש&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��@�s�Y|8]� m�P]\@d mk�c��T0 k� �ϩ�ө&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��C�s�Y|8]� m�P]\@d mk�c��T0 k� �Ϩ�Ө&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��C�s�Y|8]� m�P]\@d mk�c��T0 k� �Ϩ�Ө&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��C�s�Y|8]� m�P]\@d mk�c��T0 k� �˨�Ϩ&�1D"3Q	2�D 3Q  ��    �����O�A��D�[�.��C�s�Y|8]� m�P]\@d mk�c��T0 k� �˨�Ϩ&�1D"3Q	2�D 3Q  ��    �����O�A��A�[�.��C�o�Y|8]� m�P]\@d mk�c��T0 k� �ǧ�˧&�1D"3Q	2�D 3Q  ��    �����O�A��A�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� �ǧ�˧&�1D"3Q	2�D 3Q  ��    �����O�A��A�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� �ǧ�˧&�1D"3Q	2�D 3Q  ��    �����O�A��A�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� �ç�ǧ&�1D"3Q	2�D 3Q  ��   ������O�A��A�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� �ç�ǧ&�1D"3Q	2�D 3Q  ��    ������K�A��D�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� ����æ&�1D"3Q	2�D 3Q  ��    ������K�A��D�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� ����æ&�1D"3Q	2�D 3Q  ��    ������K�A��D�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� ����æ&�1D"3Q	2�D 3Q  ��    ������K�A��D�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������K�A��D�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������K�A��D�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������K�A��D�[�.��C�o�Y|8]� m�P]X@d mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������K�A��D�[�.��K�o�Y|8]� m�P]X@d mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������G�A��D�_�.��K�o�Y|8]� m�P]X@d mk�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������ fC�#�E엛�	C���`�����hfM߽w���c��T0 k� <�����&�1D"3Q	2�D 3Q ��_    ����:�fC�#�E����	C���`�����\eM׽o���c��T0 k� ������&�1D"3Q	2�D 3Q ��_    ����9�fC��E����	C��`������TeM˽g���c��T0 k� ������&�1D"3Q	2�D 3Q ��_    ����8�fC��E���	C�w�`������LeM���_���c��T0 k� ������&�1D"3Q	2�D 3Q ��_    ����8	��fC��E�w��x	E�o�`�����DdM���[���c��T0 k� ������&�1D"3Q	2�D 3Q ��_    ����8	��fC���E�o��l	E�g�`�����<dm���S���c��T0 k� ������&�1D"3Q	2�D 3Q ��_    ����8	��fOM��E�k��d	E�_�`�����4dm���K���c��T0 k� ������&�1D"3Q	2�D 3Q ��_    ����8	��fOM�E�[��T	E�O�`���ג�$cm���;����c��T0 k� ������&�1D"3Q	2�D 3Q ��_    ����8	��fOM۾E�S��L	E�G�`���ϓ�bm���3����"���T0 k� ������&�1D"3Q	2�D 3Q ��_    ����8	��fOMӽE�O��D	E�?�`���˓�b}{��+����"���T0 k� ������&�1D"3Q	2�D 3Q ��_    ����8	��fOM˼E�G��<	E�7�`���Ó�a}o��#����"���T0 k� L���ë&�1D"3Q	2�D 3Q	 ��_    ����8	��fOMûE�G��0	E�/�`��뿔�a}g������"���T0 k� Lì�Ǭ&�1D"3Q	2�D 3Q	 ��_    ����8	��fOM��FG��(	E�'�`��뷔��`}_������"���T0 k� LǬ�ˬ&�1D"3Q	2�D 3Q	 ��_    ����8	��fOM��FC�� 	E��`��볔��_}S������"���T0 k� Lˬ�Ϭ&�1D"3Q	2�D 3Q	 ��_    ����8	��fOM��FC��	E��`��믕��_�K������"���T0 k� LϬ�Ӭ&�1D"3Q	2�D 3Q
 ��_    ����8	��fOM��FC��	E��`��맕��^�C�������"���T0 k� ,ӭ�׭&�1D"3Q	2�D 3Q
 ��_    ����8	��fOM��F?��	E��`���맖��]�;�������"���T0 k� ,׭�ۭ&�1D"3Q	2�D 3Q
 ��_    ����8	��fOM��F?�� 	E���`���룗��\�3������"���T0 k� ,ۭ�߭&�1D"3Q	2�D 3Q
 ��_    ����8	��fOM��E�?���	E���`���룘��[�'������"���T0 k� ,߮��&�1D"3Q	2�D 3Q
 ��_    ����8	��fOM��E�?���	E]�`���럙��Z���ۂ���c��T0 k� ,���&�1D"3Q	2�D 3Q
 ��_    ����8	��fOM�E�?���	E]�`��럚�Y���ӂ���c��T0 k� <���&�1D"3Q	2�D 3Q
 ��_    ����8	��fOMw�E�?���	E]ߍ`��뛛�X���˂���c��T0 k� <���&�1D"3Q	2�D 3Q
 ��_    ����8	��fOMs�E�?���	E]׎`��뛜�W���Ã ��c��T0 k� <���&�1D"3Q	2�D 3Q
 ��_    ����8	��fOMk�B�?��	E]ώ`��뗝�V���� ��c��T0 k� <���&�1D"3Q	2�D 3Q
 ��_    ����8	��fOMc�B�?��	E]ǎ`��;���U���� ��c��T0 k� <����&�1D"3Q	2�D 3Q
 ��_    ����8	��fOM_�B�C��	E]��`��;���T���� ��c��T0 k� ������&�1D"3Q	2�D 3Q
 ��_    ����8	��fOMW�B�C��	E]��`�߯;���S���� ��c��T0 k� ������&�1D"3Q	2�D 3Q
 ��_    ����8	��fEMO�B�C��	E�`�߯;��ۘR���� ��c��T0 k� �����&�1D"3Q	2�D 3Q
 ��_    ����8	�xfEMC�B�G��	Eퟏ`�׮+��ېO|ӵ�� ��c��T0 k� ����&�1D"3Q	2�D 3Q
 ��_    ����8	�xfEM?�B�K��	E헏`�Ӯ+��یN|ϵ� ��"���T0 k� ����&�1D"3Q	2�D 3Q	 ��_    ����8	�tfEM7�B�K��	E퓏`�Ӯ+��ۈM|ǵw� ��"���T0 k� ����&�1D"3Q	2�D 3Q	 ��_    ����8	�tfE=3�B�O�|	E틐`�Ϯ+��ۄK|��o� ��"���T0 k� ����&�1D"3Q	2�D 3Q	 ��_    ����8	�pfE=+�B�S�t	E탐`�Ϯ+��ۀJ|��g���"���T0 k� ����&�1D"3Q	2�D 3Q	 ��_    ����8	�pfE='�B�W�l	E�{�`�˭����|Il��[��"���T0 k� ����&�1D"3Q	2�D 3Q ��_    ����8	�pfE=�B�W�d	E�s�`�˭����xHl��S�w�"���T0 k� M���&�1D"3Q	2�D 3Q ��_    ����8	�lfE=�B�[�\	E�k�`�˭����xFl��K�o�"���T0 k� M��#�&�1D"3Q	2�D 3Q ��_    ����8	�lfE=�B�_�T	E�c�`�˭����tEl��C�k�"���T0 k� M#��'�&�1D"3Q	2�D 3Q ��_    ����8	�lfE=�B�_�@	E�S�`�ǭ+��pBl��3�[�"���T0 k� M+��/�&�1D"3Q	2�D 3Q ��_    ����8	�hfE=�B�_�8	E�K�`�Ǯ+��lAl��+�S�"���T0 k� -/��3�&�1D"3Q	2�D 3Q ��_    ����8	�hfE,��B�_�0	E�C�`�Ǯ+��l?l��#�O�c��T0 k� -3��7�&�1D"3Q	2�D 3Q ��    ����8	�hfE,��B�[�(	E�;�`�Ǯ+��h>l���G�c��T0 k� -7��;�&�1D"3Q	2�D 3Q �� 	   ����8	�hfE,�B�[� 	E�3�`�Ǯ+��h<l���< c��T0 k� -?��C�&�1D"3Q	2�D 3Q ��D 	   ����8	�hfE,�B�[�	E�/�`�î+��l;����4c��T0 k� -;��?�&�1D"3Q	2�D 3Q ��D 	   ����8	�hfE,�B�[��	E�/�`�î+��l9�����,c��T0 k� �7��;�&�1D"3Q	2�D 3Q ��D 	   ����8	�hfE,�B�[��	E�+�`�î+��l7�����(c��T0 k� �7��;�&�1D"3Q	2�D 3Q ��D 	   ����8	�hfE,ߕB�[���	E�#�`�î��p6����� c��T0 k� �3��7�&�1D"3Q	2�D 3Q ��D 	   ����8	�hfE,ۓB�[���	E��`�î���p4�����c��T0 k� �+��/�&�1D"3Q	2�D 3Q ��D 	   ����8�hfE,ϐB�_���	E��`������t1<���ӈ�c��T0 k� �#��'�&�1D"3Q	2�D 3Q  ��D 	   ����8�hfE,ˏB�_���	F�^{�����x0<���ˈ� c��T0 k� �'��+�&�1D"3Q	2�D 3Q  ,�D 	   ����8�hfE,ǍB�_���	F�^{�����x.<��PÈ��c��T0 k� -+��/�&�1D"3Q	2�D 3Q  ��D 	   ����8�hfE,ËB�_���	F�^{î���|-<��P����c��T0 k� -+��/�&�1D"3Q	2�D 3Q  ��D 	   ����8�hfE��B�_���	F�^{ï����+<��P����c��T0 k� -+��/�&�1D"3Q	2�D 3Q  ��D 	   ����8�hfE��B�c��	F�^{ï����*<��P����c��T0 k� -+��/�&�1D"3Q	2�D 3Q ��D 	   ����8�hfE��B�c��	F��`;ï����),��P����	c��T0 k� -+��/�&�1D"3Q	2�D 3Q ��D 	   ����8�hfE��B�c���	B\��`;ǰ�����&,��P����
c��T0 k� �#��'�&�1D"3Q	2�D 3Q ��D 
   ����8�hfE��B�c���	B\��`;˰�����$,��P����c��T0 k� ����&�1D"3Q	2�D 3Q ��D 
   ����8MhfE��B�c���	B\��`;˱�����#,��P���c��T0 k� ����&�1D"3Q	2�D 3Q ��D 
   ����8MhfE�B�c���	B\�`;ϲ�����",��@w���c��T0 k� ����&�1D"3Q	2�D 3Q ��D 
   ����8MhfE�Jc��|	B\�_�ϲ�����!,��@o���c��T0 k� ����&�1D"3Q	2�D 3Q ��D 
   ����8MhfE��Jc��t	B\�_�ӳ����,��@g���c��T0 k� ����&�1D"3Q	2�D 3Q ��D 
   ����8MhfE��Jc��l	B\�_�Ӵ������@[���c��T0 k� ����&�1D"3Q	2�D 3Q ��D 
   ����8 hfE���J_��\	B\�_�۶������@K���c��T0 k� -���&�1D"3Q	2�D 3Q ��D 
   ����8 hfE���B�_��P	B\�`۷������@C��c��T0 k� -���&�1D"3Q	2�D 3Q ��D 
   ����8 hfE���B�_�H	B\�`߸������@;��c��T0 k� -���&�1D"3Q	2�D 3Q ��D 
   ����8 lfE���B�_�@	B\�`߹������@3�xc��T0 k� -���&�1D"3Q	2�D 3Q ��D 
   ����8 lfE���B�_�8	Bl�`���������+�tc��T0 k� -���&�1D"3Q	2�D 3Q ��D    ����8�pfE���B�_�(	Bl�`�����������dc��T0 k� =���&�1D"3Q	2�D 3Q ��D    ����9�pfE���B�c�� 	Bl�`����������\c��T0 k� =���&�1D"3Q	2�D 3Q ��D    ����:�tfE���B�c��	Bl�`[������������Tc��T0 k� =���&�1D"3Q	2�D 3Q ��D    ����;�tfE���B�c��	F�`[������ �������Lc��T0 k� =���&�1D"3Q	2�D 3Q ��D    ����<�xfE���B�g��	F�`[������ �������Dc��T0 k� =���&�1D"3Q	2�D 3Q  ��D    ����=�|fE���B�k���	F�`[������!������4c��T0 k� -���&�1D"3Q	2�D 3Q  ��D    ����>��fB���B�k�<�F�`[������!ܻ��ߐ�,c��T0 k� -���&�1D"3Q	2�D 3Q  /�D    ����?��fB���B�o�<�F�`[�����"ܿ��ב�$c��T0 k� -���&�1D"3Q	2�D 3Q  ��D    ����@��fB���B�s�<�F�`\����#����ǒ�c��T0 k� -���&�1D"3Q	2�D 3Q  ��D    ����A��fB���B�w�<�F��Y|�����#������	�c��T0 k� M���&�1D"3Q	2�D 3Q  ��D    ����C��fB�ÉB�{�	��E���Y|���� $������	�c��T0 k� M���&�1D"3Q	2�D 3Q  ��D    ����E��fB�ǊB��	��E���Y|��#��$������	� c��T0 k� M���&�1D"3Q	2�D 3Q  ��D    ����H��fB�ϊB���	��E���Y|��3��%������	��c��T0 k� M��#�&�1D"3Q	2�D 3Q  �D    ����K��fB�ӋB���	��E��Y���;��%���O��	��c��T0 k� �#��'�&�1D"3Q	2�D 3Q  ��O    ����N��fB�׋B���	̠g��Y���C�� &���O��	��c��T0 k� �'��+�&�1D"3Q	2�D 3Q  ��O    ����QͬfB�یB̓�	̜g��Y���K��(&���O��	��c��T0 k� �+��/�&�1D"3Q	2�D 3Q  ��O    ����T͸fB��B̟�	̐g��Y�#��W��4'���Os�	��c��T0 k� �3��7�&�1D"3Q	2�D 3Q  ��O    ����WͼfB��Ḅ�	̈g��Y�'��_��<'���Ok�	��c��T0 k� �7��;�&�1D"3Q	2�D 3Q  ��O    ����Y��fB��B̧��g��Y�+��g��D(���Oc���c��T0 k� �;��?�&�1D"3Q	2�D 3Q  ��O    ����[��fB���B̯��|g�#�Y�+��s��H(��O[���c��T0 k� �?��C�&�1D"3Q	2�D 3Q  ��O   ����]��fB��B̻��pg�/�Y�3����X)��OK��c��T0 k� �G��K�&�1D"3Q	2�D 3Q  ��O    ����_��fB��B̿��hg�3�Y�3����`)��?C��c��T0 k� �K��O�&�1D"3Q	2�D 3Q  ��O    ����a��eB��B�ǭ�dg�7�Y�7����d*��?;��c��T0 k� �O��S�&�1D"3Q	2�D 3Q  ��O    ����c��eB��B�˭�\g�;�Y�7����l+��?3��c��T0 k� �S��W�&�1D"3Q	2�D 3Q  ��O    ����e��eB�#�B�ۭ�Pg�C�Y�7����|,�'�?'��c��T0 k� �[��_�&�1D"3Q	2�D 3Q  ��O    ����g��eB�+�B�߭�Hg�G�Y|;������-�+�?�>�c��T0 k� �_��c�&�1D"3Q	2�D 3Q  ��O    ����i�dB�3�B���@g�K�Y|;������-�/�?�>�c��T0 k� �c��g�&�1D"3Q	2�D 3Q  ��O    ����k�dB�?�B����4g�W�Y|;������/�;�?�>|c��T0 k� �k��o�&�1D"3Q	2�D 3Q  ��O    ����m�cB�G�E����,g�[�Y|;������0�?�?�>tc��T0 k� �o��s�&�1D"3Q	2�D 3Q  ��O    ����o� cE�O�E���$g�_�Y|;�	�����1�C�>��>pc��T0 k� �s��w�&�1D"3Q	2�D 3Q  ��O    ����q�$bE�W�E��� g�c�Y|;�	�����2�G�>�>hc��T0 k� �w��{�&�1D"3Q	2�D 3Q  ��O    ����s�,bE�_�E���g�g�Y|;�	�����2�O�.�>`c��T0 k� �{���&�1D"3Q	2�D 3Q  ��O    ����u~<`E�o�E�#���g�o�Y|;�	�����4�W�.߭>Pc��T0 k� ������&�1D"3Q	2�D 3Q  ��O    ����w~D`E�w�D�+���g�s�Y|;�
���5�[�.ۮ�Lc��T0 k� ������&�1D"3Q	2�D 3Q  ��O    ����y~H_E��D�/���g�w�Y|;�
���6�_�.Ӱ�Dc��T0 k� ������&�1D"3Q	2�D 3Q  ��O   ����{~P^E���D�7����g�w�Y|;�
���7�_�.ϱ�<c��T0 k� ������&�1D"3Q	2�D 3Q  ��O    ����|~\]Dݗ�D�G����g��Y|;�
��9�k�.ô�,c��T0 k� ������&�1D"3Q	2�D 3Q  ��O    ����~~d\Dݟ�D�O����Q=��Y|;�	�#��:�o�.���$c��T0 k� ������&�1D"3Q	2�D 3Q  ��O   ����~l[Dݧ�D�W���Q=��Y|;�	�'��;�o�.��� c��T0 k� ������&�1D"3Q	2�D 3Q  ��O    �����~pZDݯ�D�_���Q=��Y|;�	�+�<�w�.���c��T0 k� ������&�1D"3Q	2�D 3Q  ��H    �����~|WDݿ�D�o���Q=��Y|;�	�7��>��.���c��T0 k� ������&�1D"3Q	2�D 3Q  ��H    �����~�VD�ǜE�{���Q=��Y|;�
;��?���.��� c��T0 k� ������&�1D"3Q	2�D 3Q  ��H    �����~�UD�ϝE������Q=��Y|;�
?��$@�������c��T0 k� ������&�1D"3Q	2�D 3Q  ��H    �����n�RE�ߞE������Q=��Y|;�
K��4B�������	c��T0 k� ������&�1D"3Q	2�D 3Q  ��(    �����n�QE��E������Q=��Y|;�
O��<C�������c��T0 k� ������&�1D"3Q	2�D 3Q  ��(    �����n�PE��E������Q=��Y|;��S�	=@D�������c��T0 k� ������&�1D"3Q	2�D 3Q  ��(    �����n�ME���E�����Q=��Y|;��[�	=PF�������c��T0 k� ������&�1D"3Q	2�D 3Q  ��(    �����>�LE��E�����Q=��Y|;��_�	=XF�������c��T0 k� ������&�1D"3Q	2�D 3Q  ��(    �����>�JE��E�����Q=��Y|;��g�	=\G�������c��T0 k� ������&�1D"3Q	2�D 3Q  ��(    �����>�IE��Dݻ���Q=��Y|;��k�	=dH�������c��T0 k� ������&�1D"3Q	2�D 3Q  ��(    �����>�FE�'�D�˿��Q=��Y|;��s�	MpI�������c��T0 k� ������&�1D"3Q	2�D 3Q  ��(    �����>�DE�/�D�����Q=��Y|;��{�	MtJ������� c��T0 k� �����&�1D"3Q	2�D 3Q  ��(    �����>�CE~7�D�����Q=��Y|;���	M|K���������c��T0 k� ����&�1D"3Q	2�D 3Q  ��(    �����>�@E~C�D����Q=��Y|;����	M�L���������c��T0 k� ����&�1D"3Q	2�D 3Q  ��(    �����n�>E~K�D����Q=��Y|;�}��	=�L��������c��T0 k� ���#�&�1D"3Q	2�D 3Q  ��(    �����n�<E~S�D�����Q=��Y|;�}��	=�M��������c��T0 k� �'��+�&�1D"3Q	2�D 3Q  ��(    �����n�9E~c�D����Q=��Y|;�}��	=�N�����c��T0 k� �7��;�&�1D"3Q	2�D 3Q  ��(    �����n�7E~g�D����Q=��Y|;�}��	=�N�#���w�c��T0 k� �3��7�&�1D"3Q	2�D 3Q  ��(    �����n�6E~o�E����Q=��Y|;�}��	M�N�+���s�c��T0 k� �3��7�&�1D"3Q	2�D 3Q  ��(    �����n�4E~w�E�+���Q=��Y|;�}��	M�O�3���o�c��T0 k� �3��7�&�1D"3Q	2�D 3Q  ��(   �����n�0E~��E�;���Q=��Y|;�}��	M�O�?���c�c��T0 k� �?��C�&�1D"3Q	2�D 3Q  ��(    �����n�/E~��E�C���Q=��Y|;�}��	M�O�G���_�c��T0 k� �?��C�&�1D"3Q	2�D 3Q  ��(    �����n�-E~��E~K��#�Q=��Y|;�}��	=�O�O����[�c��T0 k� �@ �D &�1D"3Q	2�D 3Q  ��(    �����^�+En��E~S��'�Q=��Y|;�m��	=�P�W����W�c��T0 k� �H�L&�1D"3Q	2�D 3Q  ��(    �����^�'En��E~c��/�Q=��Y|;�m��	=�P�c����O�c��T0 k� �T�X&�1D"3Q	2�D 3Q  ��(    �����^�&En��E~k��3�Q=��Y|;�m��	=�P�k����O�c��T0 k� �X�\&�1D"3Q	2�D 3Q  ��(    �����^�$En��E~s��7�Q=��Y|;�m��	M�P�s�ާ��K�c��T0 k� �`�d&�1D"3Q	2�D 3Q  ��(    �����^�"D>��E~{��?�Q=��Y|;�m��	M�P�{�ާ��G�c��T0 k� �h�l&�1D"3Q	2�D 3Q  ��(    �����^�!D>��E~���C�Q=��Y|;�m��	M�P��ޫ��C�c��T0 k� �l�p&�1D"3Q	2�D 3Q  ��(    �����^�D>��E~���K�Q>�Y|;�m��	M�P΋�޳��?�c��T0 k� �t
�x
&�1D"3Q	2�D 3Q  ��(    �������D>��E~���S�Q>�Y|;�]��	=�PΓ�޷��?�c��T0 k� �x
�|
&�1D"3Q	2�D 3Q  ��(    �������En��E~���W�Q>�Y|;�]��	=�PΗ�޻��;�c��T0 k� ��
��
&�1D"3Q	2�D 3Q  ��(    �������En��E~���[�Q>�Y|;�]��	=�PΛ�޿��;�c��T0 k� ����&�1D"3Q	2�D 3Q  ��(    �������En��E~���g�Q>�Y|;�]��	=�PΤ ����;�c��T0 k� ����&�1D"3Q	2�D 3Q  ��(    �������En��E~���k�Q>�Y|;�]��	M�PΨ����7�c��T0 k� ����&�1D"3Q	2�D 3Q  ��(    �������En��E~���s�Q>�Y|;�]��	M�Pά����7�c��T0 k� ����&�1D"3Q	2�D 3Q  ��(    �������En��E~���w�Q>�Y|;�]��	M�Pά����7�c��T0 k� ����&�1D"3Q	2�D 3Q  �(    ������En��En�����Q>�Y|;�]��	M�P^�����7�c��T0 k� ����&�1D"3Q	2�D 3Q  ��(    ������En��En�����Q>#�Y|;���	=�P^�����7�c��T0 k� ����&�1D"3Q	2�D 3Q  ��(    ������En��En�����Q>#�Y|;���	=�P^�����7�c��T0 k� �|	��	&�1D"3Q	2�D 3Q  ��(    ������En��En�����Q>'�Y|;���	=�P^�����;�c��T0 k� �x�|&�1D"3Q	2�D 3Q  ��(    �����.�E^��En��L��Q>+�Y|;���	=�P^�����;�c��T0 k� �p�t&�1D"3Q	2�D 3Q  �(    �����.�E^��En��L��Q>/�Y|;�]�� m�P^���� m;�c��T0 k� �l�p&�1D"3Q	2�D 3Q  �(    �����.�E^��En��L��Q>3�Y|;�]�� m�P^�O� m;�c��T0 k� �h�l&�1D"3Q	2�D 3Q  ��(    �����.�E^��En��L��Q>3�Y|;�]�� m�P^�O� m;�c��T0 k� �d�h&�1D"3Q	2�D 3Q  ��(    �����.�E^��D.��L��Q>7�Y|;�]�� m�P^�O� m?�c��T0 k� �`�d&�1D"3Q	2�D 3Q  ��(    ������E^��D.��,��Q>7�Y|;�]�� m�Pn� O� m?�c��T0 k� �X�\&�1D"3Q	2�D 3Q  ��(    ������E^��D.��,��Q>;�Y|;�]�� m�Pn�O� m?�c��T0 k� �X �\ &�1D"3Q	2�D 3Q  �/    ������E^��D.��,˥Q>?�Y|;�]�� m�Pn�O#� m?�c��T0 k� �P �T &�1D"3Q	2�D 3Q  ��/    ������E^��On��,ϥQ>C�Y|;�]�� m�Pn�O+� m?�c��T0 k� �O��S�&�1D"3Q	2�D 3Q  ��/    ������E^��On��,ץQ>C�Y|;�]�� m�P�O/� m?�c��T0 k� �O��S�&�1D"3Q	2�D 3Q  ��/    ������EN��On��,ۥQ>G�Y|;�]�� m�P�O3� mC�c��T0 k� �K��O�&�1D"3Q	2�D 3Q  ��/    ������EN��On��,�Q>G�Y|;�]�� m�P�O7� mC�c��T0 k� �G��K�&�1D"3Q	2�D 3Q  ��/    ������EN��On���Q>K�Y|;�]�� m�P|O;� mC�c��T0 k� �C��G�&�1D"3Q	2�D 3Q  ��/    ������EN��On���Q>O�Y|;�]�� m�PxO?� mC�c��T0 k� �C��G�&�1D"3Q	2�D 3Q  ��/    ������EN��On����Q>O�Y|;�]�� m�P.tOG� mC�c��T0 k� �?��C�&�1D"3Q	2�D 3Q  ��/    ������EN��On����Q>S�Y|;�]�� m�P.pOK� mC�c��T0 k� �;��?�&�1D"3Q	2�D 3Q  ��/    ������EN��On���Q>S�Y|;�]�� m�P.lOO� mC�c��T0 k� �7��;�&�1D"3Q	2�D 3Q  ��/    ������EN��On����Q>W�Y|;�]�� m�P.dOS� mG�c��T0 k� �7��;�&�1D"3Q	2�D 3Q  ��/    ������E>��On����Q>W�Y|;�]�� m�P.`OW� mG�c��T0 k� �3��7�&�1D"3Q	2�D 3Q  ��/    ������E>��On����Q>[�Y|;�]�� m�P.\O[� mG�c��T0 k� �/��3�&�1D"3Q	2�D 3Q  ��/    ������E>��On����Q>[�Y|;�]�� m�P>XO_� mG�c��T0 k� �+��/�&�1D"3Q	2�D 3Q  ��/    ������E>��On���#�Q>_�Y|;�]�� m�P>TOc� mG�c��T0 k� �+��/�&�1D"3Q	2�D 3Q  ��/    ������E>��On���+�Q>_�Y|;�]�� m�P>POg� mG�c��T0 k� �'��+�&�1D"3Q	2�D 3Q  ��/    ������E>��On���/�Q>_�Y|;�]�� m�P>LOh  mG�c��T0 k� �#��'�&�1D"3Q	2�D 3Q  ��/    ������E>��On���7�Q>c�Y|;�]�� m�P>HOl  mG�c��T0 k� �#��'�&�1D"3Q	2�D 3Q  ��/    ������E>��On���;�Q>c�Y|;�]�� m�P>DOp  mK�c��T0 k� ���#�&�1D"3Q	2�D 3Q  ��/    ������E>��On� �C�Q>g�Y|;�]� m�P>@Ot mK�c��T0 k� ����&�1D"3Q	2�D 3Q  ��/    ������CN��On� �G�Q>g�Y|;�]� m�P><Ox mK�c��T0 k� ����&�1D"3Q	2�D 3Q  ��/    ������CN��On��O�Q>k�Y|;�]{� m�P>8O| mK�c��T0 k� ����&�1D"3Q	2�D 3Q  ��/    ������CN��On��S�Q>k�Y|;�]{� m�P>4O� mK�c��T0 k� ����&�1D"3Q	2�D 3Q  ��/    ������CN��On��[�Q>k�Y|;�]{� m�P>4O� mK�c��T0 k� ����&�1D"3Q	2�D 3Q  ��/    �����^�CN��On��_�Q>o�Y|;�]w� m�P>0O� mK�c��T0 k� ����&�1D"3Q	2�D 3Q  ��/    �����^|CN��On��c�Q>o�Y|;�]w� m�P>,O� mK�c��T0 k� ����&�1D"3Q	2�D 3Q  ��/    �����^|CN��En��k�Q>s�Y|;�]s� m�P>(O� mK�c��T0 k� ����&�1D"3Q	2�D 3Q  ��/    �����^xCN��En��o�Q>s�Y|;�]s� m�P>$O� mO�c��T0 k� ����&�1D"3Q	2�D 3Q  ��/    �����^tCN��En��s�Q>s�Y|;�]s� m�P> O� mO�c��T0 k� ����&�1D"3Q	2�D 3Q  ��/    �����^tCN��En��w�Q>w�Y|8 ]o� m�P> O� mO�c��T0 k� �����&�1D"3Q	2�D 3Q  ��/    �����^pCN��En���Q>w�Y|8 ]o� m�P>O� mO�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����^pCN��E^����Q>{�Y|8 ]o� m�P>O� mO�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����^lC^��E^����Q>{�Y|8 ]k� m�P>O� mO�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����^hC^��E^����Q>{�Y|8 ]k� m�P>O� mO�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����^hC^��E^����Q>�Y|8 ]k� m�P>O� mO�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����^dC^��E^����Q>�Y|8 ]g� m�P>O� mO�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����^dC^��C�����Q>�Y|8 ]g� m�P>O� mO�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����^`C^��C�����QN��Y|8 ]g� m�P>O� mO�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n`C^��C�����QN��Y|8 ]c� m�P>O� mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n\C^��C�����QN��Y|8 ]c� m�P> O� mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n\C^��C�����QN��Y|8 ]c� m�P=�O� mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nXC^��C�����QN��Y|8 ]c� m�P=�O� mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nTC^��C�����QN��Y|8 ]_� m�P=�O� mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nTCn��C�����QN��Y|8 ]_� m�P=�O� mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nPCn��C�����QN��Y|8 ]_� m�P=�O� mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nPCn��C�����QN��Y|8 ][� m�P=�O� mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nLCn��C���æU��Y|8 ][� m�P=�O� mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nHCn��C���ǦU��Y|8 ][� m�P=�O� mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nHCn��C���˦U��Y|8 ][� m�P=�O�	 mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nDCn��C���ϦU��Y|8 ]W� m�P=�O�	 mS�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nDCn��C���ϦU��Y|8 ]W� m�P=�O�	 mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n@Cn��C�|�ӦU��Y|8 ]W� m�P=�O�	 mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n<E���C�x�צU��Y|8 ]W� m�P=�O�	 mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n<E���C�t�ۦU��Y|8 ]S� m�P=�O�
 mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n8E���C�p�ߦU��Y|8 ]S� m�P=�	O�
 mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n8E���C�l��E���Y|8 ]S� m�P=�	O�
 mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n4E���C�h��E���Y|8 ]S� m�P=�	O�
 mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n0E���C�d��E���Y|8 ]S� m�P=�	O�
 mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n0E���C�`��E���Y|8 ]O� m�P=�	O� mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n,E���C�\��E���Y|8 ]O� m�P=�	O� mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n,E���C�X ��K���Y|8 ]O� m�P=�	O� mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n(E���C�W���K���Y|8 ]O� m�P=�	O� mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n(C���C�S����K���Y|8 ]O� m�P=�	O� mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/   �����n$C���C�K����K���Y|8 ]K� m�P=�	O� mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n$C���K�G����K���Y|8 ]K� m�P=�	O� mW�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n C���K�C����K���Y|8]K� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����n C���K�?���K���Y|8]K� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nC���K�;���K���Y|8]K� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��/    �����nC���K�7���K���Y|8]G� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �����nE���K�/���K���Y|8]G� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��   �����nE���K�+���K���Y|8]G� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �����nE���K�'���K���Y|8]G� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �����nE���K�#���K���Y|8]G� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �����nE���K����K���Y|8]C� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��   �����nE���K����K΃�Y|8]C� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �����nE���K����K΃�Y|8]C� m�P=�
O� m[�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �����nE���K���#�K΃�Y|8]C� m�P=�
@  m[�c��T0 k� �����&�1D"3Q	2�D 3Q  ��    �����nE���K���'�K��Y|8]C� m�P=�
@  m[�c��T0 k� �����&�1D"3Q	2�D 3Q  ��    �����nE���L��'�K��Y|8]C� m�P=�@ m[�c��T0 k� �{���&�1D"3Q	2�D 3Q  ��    �����^AÿL��+�K��Y|8]?� m�P=�@ m[�c��T0 k� �w��{�&�1D"3Q	2�D 3Q  ��    �����^AþL��/�K��Y|8]?� m�P=�@ m[�c��T0 k� �w��{�&�1D"3Q	2�D 3Q  ��    �����^A��L���/�K�{�Y|8]?� m�P=�@ m[�c��T0 k� �s��w�&�1D"3Q	2�D 3Q  ��    �����^A��L���3�K�{�Y|8]?� m�P=�@ m[�c��T0 k� �s��w�&�1D"3Q	2�D 3Q  ��    �����^ A��L���7�K�{�a�8]?� m�P=�@ m_�c��T0 k� �o��s�&�1D"3Q	2�D 3Q  ��   �����^ A��L���7�K�{�a�8]?� m�P=�@ m_�c��T0 k� �k��o�&�1D"3Q	2�D 3Q  ��    ������ A��L���;�K�w�a�8]?� m�P=�@ m_�c��T0 k� �k��o�&�1D"3Q	2�D 3Q  ��    �������A��L���;�K�w�a�8];� m�P=�@ m_�c��T0 k� �g��k�&�1D"3Q	2�D 3Q  ��    �������A��L���;�K�w�a�8];� m�P=�@ m_�c��T0 k� �c��g�&�1D"3Q	2�D 3Q  ��    �������A��L���?�K�w�a�8];� m�P=�@ m_�c��T0 k� �c��g�&�1D"3Q	2�D 3Q  ��    �������A��L���?�K�s�a�8];� m�P=�@ m_�c��T0 k� �_��c�&�1D"3Q	2�D 3Q  ��    �������A��L���?�K�s�a�8];� m�P=�@ m_�c��T0 k� �_��c�&�1D"3Q	2�D 3Q  ��    �������A��L���?�K�s�a�8];� m�P=�@ m_�c��T0 k� �[��_�&�1D"3Q	2�D 3Q  ��    �������A��L���C�K�s�a�8];� m�P=�@ m_�c��T0 k� �W��[�&�1D"3Q	2�D 3Q  ��    �������L���L���C�K�s�a�8];� m�P=�@ m_�c��T0 k� �W��[�&�1D"3Q	2�D 3Q  ��    �������
L���L���C�K�o�Y|8]7� m�P=�@ m_�c��T0 k� �S��W�&�1D"3Q	2�D 3Q  ��    �������
L���L���C�K�o�Y|8]7� m�P=�@ m_�c��T0 k� �O��S�&�1D"3Q	2�D 3Q  ��    �������	L���L���C�K�o�Y|8]7� m�P=�@ m_�c��T0 k� �O��S�&�1D"3Q	2�D 3Q  ��    �������L���L���C�K�o�Y|8]7� m�P=�@ m_�c��T0 k� �K��O�&�1D"3Q	2�D 3Q  ��    �������L���L���C�K�o�Y|8]7� m�P=�@ m_�c��T0 k� �K��O�&�1D"3Q	2�D 3Q  ��    �������L���L�� C�K�k�Y|8]7� m�P=�@ m_�c��T0 k� �G��K�&�1D"3Q	2�D 3Q  ��    �������L���L�� C�K�k�Y|8]7� m�P=�@ m_�"���T0 k� �C��G�&�1D"3Q	2�D 3Q  ��    �������L���L�� C�K�k�Y|8]7� m�P=�@  m_�"���T0 k� �C��G�&�1D"3Q	2�D 3Q  ��    �������L���L�� C�K�k�Y|8]7� m�P=�@  m_�"���T0 k� �?��C�&�1D"3Q	2�D 3Q  ��    �������M��L�� C�K�k�Y|8]3� m�P=�@  m_�"���T0 k� �?��C�&�1D"3Q	2�D 3Q  ��    �������M��L�� nC�K�g�Y|8]3� m�P=�@  m_�"���T0 k� �;��?�&�1D"3Q	2�D 3Q  ��    �������M��L�� nC�K�g�a�8]3� m�P=�@$ m_�"���T0 k� �7��;�&�1D"3Q	2�D 3Q  ��    ������� M��L�� nC�K�g�a�8]3� m�P=�@$ m_�"���T0 k� �7��;�&�1D"3Q	2�D 3Q  ��    ��������M��L�� nC�K�g�a�8]3� m�P=�@$ m_�"���T0 k� �3��7�&�1D"3Q	2�D 3Q  ��    ��������M��L�� nC�K�g�a�8]3� m�P=�@$ mc�"���T0 k� �3��7�&�1D"3Q	2�D 3Q  ��    ��������M��L�� nC�K�g�a�8]3� m�P=�@( mc�"���T0 k� �/��3�&�1D"3Q	2�D 3Q  ��    ��������M��L�� nC�K�c�a�8]3� m�P=�@( mc�"���T0 k� �+��/�&�1D"3Q	2�D 3Q  ��    ��������M��L�� nC�K�c�a�8]3� m�P=�@( mc�c��T0 k� �+��/�&�1D"3Q	2�D 3Q  ��    ��������L���L�� nC�K�c�a�8]3� m�P=�@( mc�c��T0 k� �'��+�&�1D"3Q	2�D 3Q  ��    ��������L���L�� �C�K�c�a�8]3� m�P=�@, mc�c��T0 k� �'��+�&�1D"3Q	2�D 3Q  ��    ��������L���L�� �C�K�c�a�8]/� m�PM�@, mc�c��T0 k� �#��'�&�1D"3Q	2�D 3Q  ��    ��������L���L�� �C�K�c�a�8]/� m�PM�@, mc�c��T0 k� ���#�&�1D"3Q	2�D 3Q  ��    ��������L���L�� �C�K�c�Y|8]/� m�PM�@, mc�c��T0 k� ���#�&�1D"3Q	2�D 3Q  ��    ��������L���L�� �C�K�_�Y|8]/� m�PM�@, mc�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ��������L���L�� �C�K�_�Y|8]/� m�PM�@0 mc�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ��������L���K��� �C�K�_�Y|8]/� m�PM�@0 mc�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ��������L���K��� �C�K�_�Y|8]/� m�PM�@0 mc�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ��������A��K��� �C�@n_�Y|8]/� m�PM�@0 mc�c��T0 k� ����&�1D"3Q	2�D 3Q  ��    ��������A��K��� �C�@n_�Y|8]/� m�PM�@0 mc�"���T0 k� ����&�1D"3Q	2�D 3Q  ��    ��������A��K��� �C�@n_�Y|8]/� m�P]�@4 mc�"���T0 k� ����&�1D"3Q	2�D 3Q  ��    ��������A��K��� �C�@n_�Y|8]/� m�P]�@4 mc�"���T0 k� ����&�1D"3Q	2�D 3Q  ��    �������A��EM��C�@n_�Y|8]/� m�P]�@4 mc�"���T0 k� ����&�1D"3Q	2�D 3Q  ��    �������A��EM��C�CN_�Y|8]/� m�P]�@4 mc�"���T0 k� ����&�1D"3Q	2�D 3Q  ��    �������A��EM��C�CNc�Y|8]+� m�P]�@4 mc�"���T0 k� ����&�1D"3Q	2�D 3Q  ��    �������A��EM��C�CNc�Y|8]+� m�P]|@4 mc�"���T0 k� ����&�1D"3Q	2�D 3Q  ��    �������A��EM��C�CNc�Y|8]+� m�P]|@8 mc�"���T0 k� �����&�1D"3Q	2�D 3Q  ��    ��������A��E=��C�CNc�Y|8]+� m�P]|@8 mc�"���T0 k� �����&�1D"3Q	2�D 3Q  ��    ��������A��E=�C�CNc�Y|8]+� m�P]|@8 mc�"���T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E={�C�CNc�Y|8]+� m�P]|@8 mc�"���T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E={�C�CNc�Y|8]+� m�P]|@8 mc�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E=w�C�CNc�Y|8]+� m�P]x@8 mc�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E=w�C�CNc�Y|8]+� m�P]x@< mc�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E=s�C�@�c�Y|8]+� m�P]x@< mc�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E=o�^C�@�c�Y|8]+� m�P]x@< mc�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E-k�^C�@�c�Y|8]+� m�P]x@< mc�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E-k�^C�@�c�Y|8]+� m�P]x@< mc�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E-k�^C�CNc�Y|8]+� m�P]t@@ mc�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E-g�^C�CNc�Y|8]+� m�P]t@@ mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E-g�^C�CNc�Y|8]'� m�P]t@@ mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������A��E-g�^C�CNc�Y|8]'� m�P]t@@ mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������A��B�g�^C�CNc�Y|8]'� m�P]t@@ mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������A��B�c�^C�CNc�Y|8]'� m�P]t@@ mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ������A��B�c�^C�CNc�Y|8]'� m�P]t@@ mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������A��B�c�^C�CNc�Y|8]'� m�P]t@@ mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������A��B�c�^C�K�c�Y|8]'� m�P]p@D mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������A��E-c�^C�K�c�Y|8]'� m�P]p@D mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    ��������L���E-g�^C�K�c�Y|8]'� m�P]p@D mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���E-g�^C�K�c�Y|8]'� m�P]p@D mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���E-g�^C�K�c�Y|8]'� m�P]p@D mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���E-g�^C�K�c�Y|8]'� m�P]p@D mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���E-g�^G�K�c�Y|8]'� m�P]p@D mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���E-k�^G�K�c�Y|8]'� m�P]p@D mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���E-k�^K�K�c�Y|8]'� m�P]p@H mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���Ek�^K�K�c�Y|8]'� m�P]p@H mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �������L���Eo�^O�K�c�Y|8]'� m�P]l@H mg�c��T0 k� ������&�1D"3Q	2�D 3Q  ��    �����                                                                                                                                                                            � � �  �  �  d A�  �K����   �      6 \��7  ]�";": � �����   � �	    ����    ��|���]    ��|               	����           ��     ���   0	&


         ��6Q        ���I    ��H�����    ��_               +����          K0     ���   (	 
          ��g�  H H	     ���    ��'�����    �               J ����           �      ���   0
          ��l   � �
	   ����    ��V����    �� �                N����          ��    ���   H$
         ���l  � �	   /���    ���l��d      �^                Q	����          �p�   	  ���  03 
           	� ��	      C��     	���                            ���a              3  ���    P		 5             ���6          W�G�>    ���6�G�>                     
  I �         �     ��@   (
	           PH        k�u"     PH�u"                      
   �         �     ��@   8	 

          �<        �V�     �<�V�y      ��                  �         �     ��H    		�           �  $ $       � eQ     | `�      G               �� �         	 T`     ��@   H


         ����         ��Z:�    �����Z:�                      
    �         
 @     ��@   0
3
         ��d/ ��     � ��    ��d/ ��                            ����                ��@    		 5 	                 ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��C�  ��        �����    ��xg��;�    ���- "                 x                j  �   �   �                         ��    ��       ���      ��  ��           "                                                �                         ������������G�u�V �Z �������   	  
            
  S   i?� {��B       �� �e� �� f� �� 0g  �D  g` �� g� �d d� �D g���� ���� ����  ����. ����< ����J ����X � �D ]  (� `t� )D  u� 
�| V  
�� V  
�\ V@ 
�| W� 
�� W� 
�\ X  �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  � �c` � d` ބ �`�  � �^` � _` � }� � �j� � k�  � �m` � n`���� � ;� `j� <� k� <� k� <�  k� H� �^` I�  _� J _� J$ _� 
�\ V  
�< V  
� V@ 
�\ W� 
�< W� 
� X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������������ k  ������  
�fD
��L���"����D"� �  " `   J jF��    "�j "���
��
���     �j��  
  �
� �  �  
�       ��     ���  �   ��    ��     ���           ��     ��V          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  ���      �� �  ���        � � �  ���        �        ��        �        ��        �    ��     n������        ��                         ��q <   ��                                      �                ����             �� ���&��  ������               20 Luc Robitaille                                                                                   3  3     �[KC#d KK3]KL)cW �I c_ �c0: c�8c� �!	c� � �
ckrcs� �B� � � B� � �B� � �B� � � B� � �K � � K � �K � �K/ � � K7 � �K8 � �K; � � K= � �C � � C# � � C$ � � C% � � C& � � C' � �J� � � J� � R!c�8 b "c�0 �#"� � � $"� � �%"� � �&*� �:'"�,: ("�>*)�(**
�7 � +"K q ,"P � -"K q ."L �-  "C �- 0"B �U  "Q � 2"H �- 3"B �U  "Q �U  "Q �- 6"B �U  "Q �Y  "Q �G 9" |W :"Q �W "+ | � 
� �=� � � 
� � !� y; 
� �                                                                                                                                                                                                                 �� P         �     @ 
        �     U P E c  ��                    ������������������������������������� ���������	�
���������                                                                                          ��    �R�� ��������������������������������������������������������   �4, 9   0 #  �� �@3@�@������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ,    +    ��  �D�J      /�  	                           ������������������������������������������������������                                                                                                                                        ����  ��                                              �������������������� ��� ������ �������������������������� ���������������������� �������� ���� ���������������������������������������������������� ���������� �������� � ���� ����������  ��������������� �������� ��� �� ���� ������ ��� ���                                  E    -    �� �\�J      (E                             ������������������������������������������������������                                                                                                                      
                   ���� ��  �                                           ������������� ������������������������� �����  ��� ������������������������� ������� ��������������� ���� ������������ ��� ��������������� ��������� �������������������������������������������� ���� ������� �� �� ��������������  �                                                                                                                                                                                                                                            
                                                                                �              


             �   }�         ���          N"     8�                                                              !2  ,�      6�������������  J������������������������������������������������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � \3 �e�                                                                                                                                                                                                                                                                                           )n)n1n  Y1n        k      f      k      m      m            d      e                                                                                                                                                                                                                                                                                                                                                                                                          > �  >�  J�  <�  � #��  Cm�  ��B����f����� 6�̎�� �N ����������a�����w                       ���        $   �   & QW  �   �                  �                                                                                                                                                                                                                                                                                                                                        K K   �                      !��                                                                                                                                                                                                                            Z   �� �� ����      �� I       �������������������� ��� ������ �������������������������� ���������������������� �������� ���� ���������������������������������������������������� ���������� �������� � ���� ����������  ��������������� �������� ��� �� ���� ������ ��� ���������������� ������������������������� �����  ��� ������������������������� ������� ��������������� ���� ������������ ��� ��������������� ��������� �������������������������������������������� ���� ������� �� �� ��������������  �             $����������������˪�������������������������������������f��ff��ff�������̺�ff�fffffffffffffffffff����ƹ��ffʻfff�fffjffffffffffff��������������������ʺ��l���f˪������������������������������������������������������������������fff�fff�fff�ffk�ffi�ff��ff��ff�ffffffff�fff�x�����w��xx�������wfffffff�ffff�fffww��ww�x����wx��fk��ff��ff��ffʹffj��fʪ�f�ˊ�k������������ʚ��������������������������������������������˫��ʫ��ff��fl��fl��ff̫fff�ffʬ�f���f�����������wu���w��l������f����W��������xww��Wy�l����x������k���W�fi���j���j���f����˘�����y�y�y����������������������������������������������������ʻ����ʫɚ�����l���ƨ�lƘ�j���k���̜i���j���kxx���wx������wx������������ƈx����������������wW����w�������������������������z����������˫��̺������������������������������������������������������������ʺ������k������������������������������������������x�j���˙�x�˘��̩�x������x���xx�x������x������wx���˫��ʫ����������˪�����ʻ��������������������������������������ʻ�ʻ�����ʪ̫����˺��������������������˪�����f���k��f��fǶW�g���k���̻���f������������������x�������˩f̺�����uw�����w��x�wXx��˪�����������l����l���i��ƹx�f�������������������ʫUW��UUU�UUUX      ;      9   � ��                       f     �  �����J���J'      ��     p   �               �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��  � ��     � ��   	 ��  p �� �� ��     	Z  ��  n >�������� J  n 	Z  ��  n   )  �1   ��   ��  �� ��  � �� �� �z     &   ��� ��     ��   	 ��  c` ��  �� �� e� �� �� �z e� �� �$ 8/  ��8 /      �  ��   "�����������J  g��� 
       f ^�         �� ��      "      ��7��������J���J��a����      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                                                  U  T   T   T     T UDUDDUDDDDDDDDDDDDDDDP   E�  DU� DDU�DDDUDDDDDDDDDDDD                UP  E�  E   E                                           ���U�UTD�DDDDDDTDD TDD   �   U_ DEU�DDDUDDDDD��DZT�DDDDDDDDDDDDTDDDDDDDDUTU�����DDDDDDDDDDDEDDDEDDDDTUTU�Ԫ���Z_   P   � �U�UTDUDDDDUTD�DT��D        U_��DEU_DDD_DDDPDDE�DDE  �DD DD DD �DD �UD  �U       DZTDEDDDDE�DDE�DDE�TDDT�DE�TE���DDTU�ZD���������DDTDD��ZT�T���ZTDDE��D��T�T��DUTTT��Z��TQTDDUTD�DDDTDDD�DDDDDDE�DD_TDE�DD_ DDP DDP DD_ DU_ U�  �                                       TE�DDD�UUU                    ���DDDUUUTD  D  D  D  D  U��D�TDDDDEUUDP  DP  DP  DP  UP  TDE�DDDPUUU_                                                    wwwwtDDDt""$t"""t"w"t"w"t"w"t""$wwwwtDGtD"GtD"GtD"GtD"GtD"GtD"GtwwwwDDDD"D"""D"""DD""Gt""Gt""Gt"wwwwDDDD"B"""B""DDD"GwD"GwB$GtB$wwwwDwww$www$wwt$wwtGwwtGwwwwwwwwwwwtDDDD�DLL�D���D�D�D�t�D�t�D�wwwwDDww��Gw��Gww�Gww�Gww�Gww�Gwt"""t"w"t"w"t"w"t"""t""$tDDDwwwwD"GtD"GtD"GtD"DDD""$D""$DDDDwwww"Gt""Gt""Gt""Gt""Gt""Gt"DGtDwwwwGt"DGD"DGB$GGB$DGB""GB""GDDDwwwwwwwwwwwwwwwwDwww$www$wwwDwwwwwwwt�D�t�D�t�D�t�D�t�D�t�DMtDDDwwwww�Gww�Gww�Gww�Gw��Gw��GwDDwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "! " ""  "!  " ! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  "! ""! " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "! " ""  "!  " ! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         w 
�� ɚ� ���
�˻Ɋ�����������-� �"+ ". "$ "$ �U  Z�  Z�  J�  J�  �D  ��  ��  ɘ ˰ "  �"/�"" "  �  �            g���z��ȩ�����ة�� ���  ̰  ̰  ˰  ��  �  N�� T4�CD  CD0 C40 C30 3;� ܰ �� �� �  �  "  �""�"" �"/���  � �  �      �     �   �   ��  �"" �""  ""   "                 �   ��   �                            � "�"                  .  ".  "               �                                           � ��                  �  �˰ ��� �wp �&                     �   ���                            �   "                                                                                                                 �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp��& ��vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �" �"" �"   �                    .   .   �        �� ۼ�����wp�& vvp�ww�             �                          ��"� �"� ����                                    � ��       "   "   "�  �                            �   ���                            �   "                                                                                                   ̰ �� ̻ {��'��vz� w��  ��  ��  ̘  	�  
� "��,̻�"�� "#3  34  D  
�  �  " "" """ ! ��  ��                               ˹� �ɩ ��� �͋ ��� ��� ��̀��Ȑ���лܹнȝ0ݙ�@43�PCD�@@E�@ E�@ U�� H�  K�  �   ��    �� "�" ���                             "   "   .  ��                �   �   �   "   "   "  !�    ��                ����                         � "            � "�",�"+� ",                       "  .���"    �     �                         � ".��".��/����  �                                                                                                                                             �   �   �   r�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  bp gp �'������ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     "  �           �   �   �                     .  ". "  ""                              	�                                                                                                                                                                                                  w 
�� ɚ� ���
�˻Ɋ�����������-� �"+ ". "$ "$ �U  Z�  Z�  J�  J�  �D  ��  ��  ɘ ˰ "  �"/�"" "  �  �            g���z��ȩ�����ة�� ���  ̰  ̰  ˰  ��  �  N�� T4�CD  CD0 C40 C30 3;� ܰ �� �� �  �  "  �""�"" �"/���  � �  �      �     �   �   ��  �"" �""  ""   "                 �   ��   �                            � "�"                  .  ".  "               �                                           � ��                  �  �˰ ��� �wp �& ���������������������  ��  ��  ��  �   �    �          �         �                                �  �  "�  "   "                                                  �  �  �  �  w  �  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �           �   �     �   �             �  �� Ș ��  ��  �    �   �                               �   �   ��   ��  �   ��   �                                                                                 �  �  "   "                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��    "  "  "                       �  ��  ��  ww  &'  vv  w                �                        ��"� �"� ����                            �"  �""� "�    ��   �  ��  �  �  �         � ".��".��/����  �                                                                                                                                                              	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           "� /���  �       �   �   �                                                   ��  "   "   "  �� ��                   �".��".���                                �   O   T     ��                                 � "�"  �    � � �                           �   "                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��               �   �   "           �   �   �                                       �  ���   �                          �   �   �"  �""��� �   �      �       �                            ""  "".  . �    �                                                                                                                                            �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   �   " � ��      �    �   �   �"  ""  !� �� ��  �               �   " ��.�  ��      �    � �  �                     �         "   "   �           � ��                    ���� �                                           �   ���                            �   "                                                                                                                         	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           "� /���  �       �   �   �                       ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �                    ".  ".  ���                   ���                � ".��".��/����  �                                                                                                                                        ����������ݼ�����))�����.(����M���M D � ��� �"( ��� �� �� �  �  �   �   �  �   ��  ��� ؼ̰ڛ�˺������ɪ�۸��Ȕ͙̄̄͜Mڜ��̩U�̴@��ݿ��������ɉ��ɋ�������������𻻲  "/  ��   �   �   �   �           ��  �     "            �   �   �   ��      �   ��                          �   �   �   �   �   �   �   �   �  ��  �     ��         "  "   �"  "   �                .   .   �    �                             �          �                                                                                                                                                                                                   2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ DD D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�GwDGwqwDDwtwwww3333DDDD �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�""""����������A��I��I = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=""""�����A�DA�I��I�    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"��������I���I���I���I��� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(XxMAMAMMMM�M�M����3333DDDD w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xwwD�����MD��M����3333DDDD  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���4���4���4���4���4���43334DDDD �  + � � � � � � � � � � ��	� � � ��� � � � � � � � � � � ��	� � � ��� �� ����(+((�""""wwwwqqqqwGwGGG ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""wwwwwwqqDAwG M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M������������������333DDD � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�M��M��D��M����������3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DD��D�M��D����3333DDDD!�!�!�!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���rs��ww""""������DH�H�!�!�!�))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�tu���(+""""�������H�H��D!�!�!�5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�vw��(W(�""""��������H��H��H��H�� !�!�AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���&2�(a(�DD������L��DL����3333DDDD;'(!�AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(�L�A�AAD��DL�����3333DDDD<34!�AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� SA��l(=���4���4���4L��4L��4���43334DDDD  � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� SA��(( """"���������M�MMM X � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� SA��(Xx""""�������A��AA w � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� )��:	9ww��������������333DDD � � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(I��I����������������3333DDDD  � �!�AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((���A���I��I���I�����3333DDDD m � �!�A�A� � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""������������������������  � �!�AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M""""������D�D��� 
 � �!�AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�""""������������������������ - � �!�!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�wqwwqwwwwwqwwwDwwww3333DDDD 69�:���  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5qqwwwDDwtGwwww3333DDDD x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xwww4www4www4www4www4www43334DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwqwwwqwqwq + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""wwwwwwwDwGwA � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(��A�L�L�L��L���333DDDLDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDD[KC#d KK3]KL)cW �I c_ �c0: c�8c� �!	c� � �
ckrcs� �B� � � B� � �B� � �B� � � B� � �K � � K � �K � �K/ � � K7 � �K8 � �K; � � K= � �C � � C# � � C$ � � C% � � C& � � C' � �J� � � J� � R!c�8 b "c�0 �#"� � � $"� � �%"� � �&*� �:'"�,: ("�>*)�(**
�7 � +"K q ,"P � -"K q ."L �-  "C �- 0"B �U  "Q � 2"H �- 3"B �U  "Q �U  "Q �- 6"B �U  "Q �Y  "Q �G 9" |W :"Q �W "+ | � 
� �=� � � 
� � !� y; 
� �AqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD��������������������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ��������������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ��������������������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE��������������������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD��������������������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD��������������������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD��������������������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� ����>�L�L�T�\��=�L�S�H�U�U�L��������>��<���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� ��$��/�L�U�P�Z��=�H�]�H�Y�K���������>��<���""""������A�D��I��""""�������D����� ����7�\�J��<�V�I�P�[�H�P�S�S�L�������8�>�7���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �8�>�7������A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �>��<���!��""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,�����������DDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II�������������������������������������������������������������������������������������������������������������������������������������-�.��/�0�1�2�3������ �������������������!�"�#�4�5�$�$�$�$�$�$�$�$�%������������������&�'�(�)�*�*�*�*�*�*�*�*�*�*�+�,������������������6�7���8�9�:�;�<�=�>�?�@� �������������������!�"�#�$�$�$�$�$�$�$�A�5�$�%������������������&�B�C�D�E�F�G�H�I�J�K�L�M�N�O�P�����������������Q�R�S�T�U�V�W�X�Y�Z�X�[�\�]�^�_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            