GST@�                                                           �t�                                                      �   �   �  n  0      
      � 2�����	 ʳ����������`���t���        vh      #    t���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     "�j  " ���
��
�"    
 �j�
�
  
  ��
   �                                                                              ����������������������������������      ��    =oo 0 4gg 1                 ��                      � � � �                 �� 
         88�����������������������������������������������������������������������������������������������������������������������������oo    oo      ++    ''           ��                		  77  VV  		                              :: �����������������������������������������������������������������������������                                �?  ?       �   @  #   �   �                                                                                '"    
��      H   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E ? �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    �hU]c�A�YAd?�S�|,4hK��nLT(X�K��ZӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]_�A�YAd@�S�|,DhK��nLT(X�K��ZӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU][�A�YAd@�S�|,DhK��nLT(X�K��[ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]W�A�YAh@�S�|,DhK��nLT(X�K��[ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]S�A�YAh@�S�|,DhK��nLT(X�K��\ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]O�A�YAh@�S�|,DhK��nLT(X�K��\ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �lT]K�A�YAhA�S�|,�hK��nLT(X�K��]ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �lT]C�A�YAlA�S�|,�hK��nLT(X�K��]ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �lT]?�A�YAlA�S�|,�hK��nLT,X�L��^ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �lT];�A�YAlA�S�|,�hK��nLT,X�L��^ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �lT]7�A�YAlA�S�|,�hK��oLT,X� L��^ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �lT]3�A�YAlA�S�|,4hK��oLd,X� L��^ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �lT]/�A�YApB�S�|,4hK��oLd,X� M c�_ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �lT]+�A�YApB�S�|,4hK��oLd,X� M c�_ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �lT]'�A�YApB�S�|,4hK��oLd,X� M c�_ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �pT]#�A�YApB�S�|,4hK��oLd,Y� M c�_ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �pT]�A�YAtB�S�|,4hK��oLd,Y� N c�_ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �pT]�A�YAtB�S�|,4hK��oLd,Y� N �_ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �pT]�A�YAtC�S�|,4hK��oLd,Y� N �_ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; 	���ac�Ep�2F � �|,R|I2@-E��.A#��K�3��T0 k� ����(%2't �1"t'%  ��3    � % i	���1k�Ep�2F � �|,�|I2H,E��-A+��S�3��T0 k� ����(%2't �1"t'%  ��3    � % k	���1o�Ep�3F � �|,�|I2L,E��+Q/��[�3��T0 k� ����(%2't �1"t'%  ��3    � % m	���1s�Ep�4F � �|,�|I2T+E��)Q/��_�3��T0 k� ��� (%2't �1"t'%  ��3    � % o	���1w�Ep�4F � �|,�xI2X+E��(Q3��g�3��T0 k� ��(%2't �1"t'%  ��3    � % q	���1{�Ep�5BP� �|,�xIB\+E��&Q;��o�3��T0 k� ��(%2't �1"t'%  ��3    � % s	���a�Ep�6BP�	 �|,RxIBd*E��$Q?��s�3��T0 k� ��(%2't �1"t'%  ��3    � % u	���a��Ep�8BP� �|,RtIBl*E��!Q?����3��T0 k� �� (%2't �1"t'%  ��3    � % w	���a��D��9BQ �|,RpIBp*E��QC����3��T0 k� � �$(%2't �1"t'%  ��3    � % y	���a��D��:F �|,RlI2t)E��QG����3��T0 k� �,�0(%2't �1"t'%  ��3    � % {	���a��D� ;F �|,Bl
I2x)E��QO����3��T0 k� �8�<(%2't �1"t'%  ��3    � % }	���a��D�<F �|,Bh
I2|)E��QS����3��T0 k� �D�H(%2't �1"t'%  ��3    � % 	���a��D�>F$ �|,Bd	I2�)E��a[����3��T0 k� �P�T(%2't �1"t'%  ��3    � % � ��a��D�@F4 �|,B`E��(E��ac����3� T0 k� �`�d(%2't �1"t'%  ��3    � % � ��Q��D�$BF< �|,B\E��(E��ak����3� T0 k� �h �l (%2't �1"t'%  ��3    � % � ��Q��D�,CFD �|,BXE��(E��as����3� T0 k� �p!�t!(%2't �1"t'%  ��3    � % � ��Q��D�0DFL �|,BXE��(E��aw����3� T0 k� �x"�|"(%2't �1"t'%  ��3    � % � ��Q��D�8FFP �|,2TE��(E��a����3� T0 k� �#��#(%2't �1"t'%  ��3    � % ���Q��D�@HFX �|,2PE��(C��a���ú3� T0 k� �$��$(%2't �1"t'%  ��3    � % ���Q��D�LKFh��|,2HE��'C��	���˹3� T0 k� �&��&(%2't �1"t'%  ��3    � % ���Q��D�PLFp��|,2D@b�'C�����Ϲ3� T0 k� �'��'(%2't �1"t'%  ��3    � % ���Q��D�XNFx��|,2D@b�'C�����Ӹ3� T0 k� �(��((%2't �1"t'%  ��3    � % ���Q��D�\PF���|,2@@b�'E�����׸3�T0 k� �)��)(%2't �1"t'%  ��3    � % ���ủD�dRF���|,2<@b�'E�����۸3�T0 k� �*��*(%2't �1"t'%  ��3    � % ���ῤFpUF���|,"8E"�&E������3�T0 k� ��,��,(%2't �1"t'%  ��3    � % ��#�ῢFtWF� ��|,"4E"�&E���ú��3�T0 k� ��-��-(%2't �1"t'%  ��3    � % ��'�ῡF|YE��!��|,"4E"�&E���˹��3�T0 k� ��*��*(%2't �1"t'%  ��3    � % ��+��F�[E��"��|,"0E"�&E���ӹ��3�T0 k� ��(��((%2't �1"t'%  ��3    � % ��7��F�^E��$��|,",E"�&E���߸���3�T0 k� ��(��((%2't �1"t'%  ��3    � % ��;��F�`E��%��|,",E"�&Eѿ����3�T0 k� ��'��'(%2't �1"t'%  ��3    � % ��?��ØF�bE��&��|,�(E��&E�����3�T0 k� ��'��'(%2't �1"t'%  ��3    � % ��C��ÖF�cE��'��|,�(	E��&E������3�T0 k� ��'��'(%2't �1"t'%  ��3    � % ��K��ÒF�gE��(��|,�(
E��&E�����3�T0 k� � (�((%2't �1"t'%  ��3 	   � % ��S��ÐE��i@!�)��|,�$
E��%E��R��'�3�T0 k� �)�)(%2't �1"t'%  ��3 	   � % ��W��ÎE��j@!�*��|,"$E��%E��R��/�3�T0 k� �,*�0*(%2't �1"t'%  ��3 	   � % � [��ÏE��l@!�+��|,"$E��%E��R��3�3�T0 k� �<*�@*(%2't �1"t'%  ��3 	   � % � c�ÏE��n@",��|,"$E��%E��R#��;�3�T0 k� �L+�P+(%2't �1"t'%  ��3 	   � % � k�ǐE��qE�.��|,"$E��%E��R/��K�3�T0 k� �P-�T-(%2't �1"t'%  ��3 	   � % � s�ǑE��rE�/��|,"$E��%E��R3��S�3�T0 k� �P.�T.(%2't �1"t'%  ��3 	   � % � w�ǑE��tE�$/��|,$E"�%E��R7��W�3�T0 k� �P.�T.(%2't �1"t'%  ��3 	   � % � �ˑE��uE�,0��|,(E"�%E��R;��_�3�T0 k� �T/�X/(%2't �1"t'%  ��3 	   � % � ��˒E��wE�41� |,(E"�%E��R?��g�3�T0 k� �X0�\0(%2't �1"t'%  ��3 	   � % � ���ϒE��xE<2�|,(E"�$E��RC��o�3�T0 k� �\2�`2(%2't �1"t'%  ��3 	   � % � ���ϒE��zED3�|,(E"�$E�{�BG��w�3�	T0 k� �`4�d4(%2't �1"t'%  ��3 
   � % � ���ӓE�}ET4�|,,E"�$E�s�BO�Ї�3�	T0 k� �l7�p7(%2't �1"t'%  ��3 
   � % ����דE�~E\5�|,�0E# $E�o�BS�Ћ�3�
T0 k� �p8�t8(%2't �1"t'%  ��3 
   � % ����דE�E�d6�|,�0E# $E�k�BS�Г��
T0 k� �x=�|=(%2't �1"t'%  ��3 
   � % ����ۓE�$�E�l7�$|,�4E#$E�g�BW�Л��
T0 k� �A��A(%2't �1"t'%  ��3 
   � % ����ߔE�,�E�t7�(|,�4@c$E�c�B[�У��T0 k� �D��D(%2't �1"t'%  ��3 
   � % �����E�8E��9�4|,�8@c$F[�2_�г��T0 k� �H��H(%2't �1"t'%  ��3 
   � % �����E�@E��:�8|,�<@c$FW�2c�л��T0 k� �J��J(%2't �1"t'%  ��3 
   � % �����E�LE��;�@|,r@@c$FS�2c��î�T0 k� �K��K(%2't �1"t'%  ��3    � % �����E�T~E��<�D|,r@@c$FO�2g��Ǯ�T0 k� �M��M(%2't �1"t'%  ��3    � % �����E"\~E��=�L|,rD@c$FO�2g��Ϯ�T0 k� �O��O(%2't �1"t'%  ��3    � % ������E"d}E��=�T|,rH@c$FK�Bk��׮�T0 k� ��P��P(%2't �1"t'%  ��3    � % � ����E"t|E��?�`|,L@c#FG�Bo����T0 k� ��R��R(%2't �1"t'%  ��3    � % � ����E"|{E��@�d|,P@c#D�C�Bo����T0 k� ��S��S(%2't �1"t'%  ��3    � % � ����E"�{Er�A�l|,P@c#D�C�Bs�����T0 k� ��U��U(%2't �1"t'%  ��3    � % � ����E"�zEr�B�t|,T@c#D�G�Bs�����T0 k� ��W��W(%2't �1"t'%  ��3    � % � ����E"�yEr�C�||,X@c #D�G�Bw����T0 k� ��X��X(%2't �1"t'%  ��3    � % �!���E"�xEr�D��|,\@c #D�K�Bw����T0 k� ��Y��Y(%2't �1"t'%  ��3    � % �!���E�wEr�E��|,�`@c$#D�O�R{����T0 k� ��Z� Z(%2't �1"t'%  ��3    � % �!��+�E�vEr�H��|,�d@c(#D�S�R��#��T0 k� �]�](%2't �1"t'%  ��3    � % �!��3�E�uEs I��|,�h@c(#D�W�R��+��T0 k� �_�_(%2't �1"t'%  ��3    � % ����7�E�tEsJ��!�,�l@c(#D�[�R���3��T0 k� �`�`(%2't �1"t'%  ��3    � % ����?�E�sEsL��!�,�t@c,#D�_�R���;��T0 k� �a� a(%2't �1"t'%  ��3    � % ����C�E�sEsM��!�,�x@c,#D�c�R���?��T0 k� �$c�(c(%2't �1"t'%  ��3    � % ����K�E�rEcN��!�,�|@c0#D�g�R���G��T0 k� �b� b(%2't �1"t'%  ��3    � & ����S�E�qEc P��!�,��@c0#D�k�R���O��T0 k� �c�c(%2't �1"t'%  ��3    � ' �!#��_�E pEc,R��!�,��@c4#D�s�R���_��T0 k� �d�d(%2't �1"t'%  ��3    � ( �!'��g�EoEc0T��!�,��@c4#D�w�b���g��T0 k� �e�e(%2't �1"t'%  ��3    � ) �!+��k�EnEc8U��!�,��@c8#D�{�b���o��T0 k� �e�e(%2't �1"t'%  ��3    � * �!3��s�E�nEc<W��!�,��@c8#D� b���w��T0 k� �g�g(%2't �1"t'%  ��3    � + �!7��{�E�$mEc@Y��!�,��@c8"D�b���{��T0 k� �i� i(%2't �1"t'%  ��3    � , �8 �E�,mEcDZ��|,�@c<"D�b������T0 k� �j� j(%2't �1"t'%  ��3    � - �@�E�<lEcDZ�|,�@c<"D�2������T0 k� � l�$l(%2't �1"t'%  ��3    � . �D�E�DmEcL[�|,�E�@"D�2������T0 k� � l�$l(%2't �1"t'%  ��3    � / �L£�E�LmEcP[� |,�E�@"D�	2������T0 k� �$k�(k(%2't �1"t'%  ��3    � 0 ��P«�E�TnEST\�(|,��E�D"D�
2������T0 k� �0e�4e(%2't �1"t'%  ��3    � 1 ��T³�E�\oESX\�0|,��E�D!D�2������T0 k� �4a�8a(%2't �1"t'%  ��3    � 2 ��`
�ÛD�pqES`^�@|,��E�H!D�2������T0 k� �<^�@^(%2't �1"t'%  ��3    � 3 ��h�˛D�xrESd^�H|,��E�H I�2���Ǩ�T0 k� �@[�D[(%2't �1"t'%  ��3    � 4 ��l�כDӀsESh_�P|,��E�L I�2���Ϩ�T0 k� �DZ�HZ(%2't �1"t'%  ��3    � 5 ��t�ߛDӈtESl_�X!�,�E�LI��2���ר�T0 k� �HY�LY(%2't �1"t'%  ��3    � 6 ��x��DӐuESl`�`!�,�E�LI��2���ߨ�T0 k� �LY�PY(%2't �1"t'%  ��3    � 7 �����DӠwESta�p!�,�API��	R�����T0 k� �PY�TY(%2't �1"t'%  ��3    � 8 �����DӨwECta�x!�,�APJ�	R��	���T0 k� �TV�XV(%2't �1"t'%  ��3    � 9 ����DӰxECxa߀!�,ATJ�	R��	���T0 k� �TU�XU(%2't �1"t'%  ��3    � 9 ����DӼyECxb߈!�,ATJ�	R��	��T0 k� �XS�\S(%2't �1"t'%  ��3    � : ����D��{ECxbߐ!�,ATJ�	R��	��T0 k� �XR�\R(%2't �1"t'%  ��3    � : ���#�D��zEC|bߘ!�,AXJ�	R��	��T0 k� �XQ�\Q(%2't �1"t'%  ��3    � : ���+�D��yEC|bߠ!�,A\I��	b��	��T0 k� �\Q�`Q(%2't �1"t'%  ��3    � : ���7�D��xEC|cߨ!�,A`I��	b��	"��T0 k� �\Q�`Q(%2't �1"t'%  ��3    � ; ���G�D��wEC�c߸|, AhI��!	b��	"'��T0 k� �\Q�`Q(%2't �1"t'%  ��3    � ; ���O�D��vA�c��|,$ AlI� "	b�	"+��T0 k� �TQ�XQ(%2't �1"t'%  ��3    � ; ���W�I��uA�c��|,, ApJ#"�	"3��T0 k� �PQ�TQ(%2't �1"t'%  ��3    � ; ���_�I��uA�c��|,0!ApJ#"�	7��T0 k� �LQ�PQ(%2't �1"t'%  ��3    � ; ���g�I��tA�c��|,4"AtJ$"�	;��T0 k� �HQ�LQ(%2't �1"t'%  ��3    � ; ���s�I� sA�b��|,8"AxJ%"�	?��T0 k� �HQ�LQ(%2't �1"t'%  ��3    � ; ���{�I�rA�b��|,@#A|J&"�	C��T0 k� �PQ�TQ(%2't �1"t'%  ��3    � ; �����JqA|b��|,H$A�I�'"�	K��T0 k� �TQ�XQ(%2't �1"t'%  ��3    � ; �����JpA|b|,P%A�I� '"�	"O��T0 k� �XQ�\Q(%2't �1"t'%  ��3    � ; �����JoA|a|,T%A�I�$("�	"S��T0 k� �XP�\P(%2't �1"t'%  ��3    � ; �����JoEC|a|,�\&A�I�,)"�	"W��T0 k� �XO�\O(%2't �1"t'%  ��3    � ; �� ���JnECx`|,�`'A�I�0*"�	"W��T0 k� �XN�\N(%2't �1"t'%  ��3    � ; ��!���I�nECx`$|,�h'A�Er4+�	"[��T0 k� �XM�\M(%2't �1"t'%  ��3    � ; ��"�ǣI� mECt_4|,�t(A�Er<-�	c��T0 k� �TL�XL(%2't �1"t'%  ��3    � ; � "�ϣI�$lE3t^<|,	x)A�Er@.�	c��T0 k� �\K�`K(%2't �1"t'%  ��3    � ; �#�פI�(lE3t^D|,	|)A�ErD/�	g��T0 k� �`J�dJ(%2't �1"t'%  ��3    � ; �#�ߥJ(kE3t]L|,	�)A�ErH1�	g��T0 k� �`I�dI(%2't �1"t'%  ��3    � ; �$��J,kE3p\�T|,	�*A�ErP2�	k��T0 k� �dH�hH(%2't �1"t'%  ��3    � ; �$��J,kE3p[�\|,	�*EäErT3�	"k��T0 k� �dG�hG(%2't �1"t'%  ��3    � ; �(%���J0j@�pZ�l|,	#�*EèEb\6�"	"o��T0 k� �`E�dE(%2't �1"t'%  ��3    � ; �0&��I�0j@�lY�t|,	#�+EìEb\7�#	"o��T0 k� �`D�dD(%2't �1"t'%  ��3    � ; �8&��I�0j@�lX�||,	#�+EìEb`9�%	"s��T0 k� �`C�dC(%2't �1"t'%  ��3    � ; �<'��I�4j@�lW��|,	#�+EìEbd:�&	s��T0 k� �`B�dB(%2't �1"t'%  ��3    � ; �D'��I�4j@�lV��|,	#�+EðEbh<��(	s��T0 k� �\A�`A(%2't �1"t'%  ��3    � ; �T(�+�@4i@�hS��|,�+EӰ	Ebl?��*	s��T0 k� �\>�`>(%2't �1"t'%  ��3    � ; �\(�3�@4h@�hRФ|,�+EӰ	Ebp@��+	w��T0 k� �\=�`=(%2't �1"t'%  ��3    � ; �d)�7�@4h@�hQЬ|,�+EӰEbpB��-	"w��T0 k� �X<�\<(%2't �1"t'%  ��3    � ; �l)�?�@4g@�hPд|,�,EӰEbpC��.	"w��T0 k� �X;�\;(%2't �1"t'%  ��3    � ; �t*�C�@4g@�dNм|,�,EӰEbtE�/	"w��T0 k� �X9�\9(%2't �1"t'%  ��3    � ; 	|*�K�E�4f@�dM��|,�,EӰEbtG�0	"w��T0 k� �X8�\8(%2't �1"t'%  ��3    � ; 	�*�S�E�4e@�dJ��|,�,E�ERxJ�1 w��T0 k� �T5�X5(%2't �1"t'%  ��3    � ; 	�+�[�E�4d@�dI��|,��,E�ERxL�2 w��T0 k� �T3�X3(%2't �1"t'%  ��3    � ; 	�+�_�E�4c@�`G��|,��,E�ERxM�3 w��T0 k� �T2�X2(%2't �1"t'%  ��3    � ; 	"�+�c�E�4b@�`F��|,��,E�ERxO�$4 w��T0 k� �T0�X0(%2't �1"t'%  ��3    � ; 	"�+�k�E�4a@�`B��|,��,E�ERxR�05 w��T0 k� �P-�T-(%2't �1"t'%  ��3    � ; 	"�+�o�E�4`@�`A�|,��,ES�ERxS�05 w��T0 k� �P+�T+(%2't �1"t'%  �3    � ; 	"�+�s�E�8_@�`@�|,��,ES�ERtU�44 w��T0 k� �T+�X+(%2't �1"t'%  ��3    � ; 	�+�w�E�8]@�d?q|,��,ES�ERtV�44 bw��T0 k� �`(�d((%2't �1"t'%  �3    � ; 	�+�{�E�8[@�l>q$ |,�-ES�ERpY�83 bw��T0 k� �x#�|#(%2't �1"t'%  ��?    � ; 	�+��E�8Z@�l=q/�|,�.E�ERpZ�<2 bw��T0 k� � �� (%2't �1"t'%  ��?    � ; 	�+��E�8X@�p<q7�|,�/E�EBl\s@1 bw�"C�T0 k� ���(%2't �1"t'%  ��?    � ; 	"�+ԃ�E�8WGt<q;�|,�/E�EBl]s@1�w�"C�T0 k� ���(%2't �1"t'% ��?    � ; 	"�+ԋ�E�4TGx:qK�|,t0E�EBh_sD/�{�"C�T0 k� ���(%2't �1"t'% $�?    � ; 	"�+ԋ�E�4SG|:qS�|,t 1E�EBdasH.�{�"C�T0 k� #���(%2't �1"t'% ��?    � ; 	"�+ԏ�E�4RG�9�W�|,t$1E�EB`bsL-�{���T0 k� #���(%2't �1"t'% ��?    � ; ��+ԓ�E�4PF�8�_�|,t(2D3|EB`csL,���T0 k� #���(%2't �1"t'% ��?    � ; ��+ē�E�0OF�8�g�|,t,2D3xEB\csP+���T0 k� #���(%2't �1"t'%  ��    � ; �+ě�E�0LF�6�s�|,t04D3pEBTesT)����T0 k� #���(%2't �1"t'%  ��    � ; �+ě�E�,JF�6�{�|,t44D3hEBPfcX(����T0 k� ����(%2't �1"t'%  ��    � ; �+ė�E�,IF�5��|,t85ESdEBLgc\'�����T0 k� ����(%2't �1"t'%  �    � ; +ԏ�E�(GF�5���|,t<5ES`E2Hgc`%�����T0 k� ����(%2't �1"t'%  ��    � ;  +ԇ�E�$FF�4���|,t@6ES\E2Hhcd$�����T0 k� ����(%2't �1"t'%  ��3    � ; ,+�w�C�$FF�3���|,dH6ESPE2@i�l"�����T0 k� ����(%2't �1"t'%  ��3    � ; 0,�o�C�$EF�2���|,dL6I�LE2<i�p �����T0 k� 3���(%2't �1"t'%  ��3    � ; 8,�g�C� DF�2���|,dP6I�HE28i�x�����T0 k� 3���(%2't �1"t'%  ��3    � ; <,�c�C�DF�1���|,dT6I�DE24j�|�����T0 k� 3���(%2't �1"t'%  ��3    � ; @,�[�C�CF�1���|,dX6I�@E20j��r����T0 k� 3���(%2't �1"t'%  ��3    � ; L,�K�C�AF�0���|,d\6ES8E2,j��r����T0 k� ����(%2't �1"t'%  ��3    � ; P,�C�C�@F�/q��|,d`6ES4E"(j��r����T0 k� ����(%2't �1"t'%  ��3    � ; T,�;�C�@F�.q��|,T`6ES,E"$j��r����T0 k� ����(%2't �1"t'%  ��3    � ; \,�3�C�?F�.q��|,Td5ES(E"$j��r����T0 k� ����(%2't �1"t'%  ��3    � ; `,�+�C�>F�-q��|,Th5ES$E" j��r����T0 k� ����(%2't �1"t'%  ��3    � ; h,��C�=F�-q��|,Th5ESE�i��r����T0 k� ����(%2't �1"t'%  ��3    � ; p,��C�=F�,q��|,Tl5ESE�i��b����T0 k� ����(%2't �1"t'%  ��3    � ; p,��C�<F�,q��|,Tl5ESE�h��bå��T0 k� ����(%2't �1"t'%  ��3    � ; t,��C�<F�+q��|,Tl5ECE�h��bǤ��T0 k� ����(%2't �1"t'%  ��3    � ; t,��C�;E��+q��|,�l4EC E�g��bǣ��T0 k� ����(%2't �1"t'%  ��3    � ; |,���C�;E��)q��|,�l4EB�E�f��bˢ��T0 k� ����(%2't �1"t'%  ��3    � ; �,���C�:E��)a��|,�l4EB�CBf��bϡ��T0 k� ����(%2't �1"t'%  $�3    � ; �,���C�:E��(b�|,�l4E��CBe��bϠ��T0 k� ô��(%2't �1"t'%  ��     � ; �,���C�:E��(b�|,�l4E��CBd��Rϟ��T0 k� ô��(%2't �1"t'%  ��     � ; �,���C�:E��&b�|,�l4E��CB b��Rӝ�T0 k� ô��(%2't �1"t'%  ��     � ; �-���C�9E��&b�|,�l3E��CA�a��
RӜ�T0 k� ð��(%2't �1"t'%  ��     � ; �-���C�9E��%b�|,�h3E��CA�`��	RӜ�T0 k� ����(%2't �1"t'%  ��     � ; �-ӻ�C�9E��#b�|,Td3EҰCA�^���Ӛ�
T0 k� �� �� (%2't �1"t'%  ��     � ; �-ӳ�C�9E��"b�|,Td3EҨCA�]���ә�
T0 k� ��!��!(%2't �1"t'%  �     � ; �-ӫ�A9E��"b�|,T`3EҠE!�\���Ә�	T0 k� ��"��"(%2't �1"t'%  �     � ; ��-ӛ�A9E�� b'�|,T\3EҐE!�Z���ϗ�T0 k� ����(%2't �1"t'%  ��     � ; ��-ӓ�A9E��b'�|,D\3E�E!�X��Rϖ�T0 k� ����(%2't �1"t'%  ��     � ; ��-ӏ�A9E��b+�|,DX3E�|E!�W��R˕�T0 k� ����(%2't �1"t'%  ��     � ; ��-��A9E��b/�|,DP3E�lE!�T��Rǔ�T0 k� ����(%2't �1"t'%  ��     � ; ��-Sw�A9E��b3�|,DP3E�dE!�S��RǓ�T0 k� ����(%2't �1"t'%  ��     � ; ��-So�A9A�b7�|,4L4E�XE!�R��BÒ�T0 k� ����(%2't �1"t'%  ��     � ; ��-Sg�A9A��7�|,4L4E�PE!�P��BÒ�T0 k� ����(%2't �1"t'%  ��     � ; ��-S_�A9A��;�|,4L4E�HE!�O�� B���T0 k� ����(%2't �1"t'%  ��     � ; ��-S[�A9A��;�|,4H5E�<E!�M���B����T0 k� ����(%2't �1"t'%  ��     � ; ��-SK�A:A��C�|,4H5E�,E�J���B����T0 k� ����(%2't �1"t'%  $�     � ; ��-SC�A:A��C�|,4D6E� E�I���B����T0 k� ����(%2't �1"t'%  ��    � ; ��-S;�A:A��G�|,4D6E�E�G���B����T0 k� ����(%2't �1"t'%  ��    � ; ��,S3�A;A��G�|,4D7E�E�F���2��3�T0 k� ����(%2't �1"t'%  ��    � ; ��,S'�A;A��K�|,4D7E��E�C���2��3�T0 k� ����(%2't �1"t'%  ��    � ; 	�,S�A<A��O�|,DD8E��E�B���2��3�T0 k� ����(%2't �1"t'%  ��    � ; 	�+S�A <A��S�|,DD8E��B��@���2��3�T0 k� ����(%2't �1"t'%  ��    � ; 	�+S�A =A��S�|,D@9E��	B��?���B��s�T0 k� ����(%2't �1"t'%  ��    � ; 	�+S�A =A��W�|,D@:E��
B��>���B��s�T0 k� ����(%2't �1"t'%  ��    � ; 	�+S�A =A��W�|,D@;E��
B� =���B��s�T0 k� ����(%2't �1"t'%  ��    � ; 	�*R��A�>A��[�|,�<<E��B�:���B��s�T0 k� ��
��
(%2't �1"t'%  ��    � ; 	�*R��A�>A��_�|,�<=E�B�9���2��s�T0 k� ��
��
(%2't �1"t'%  ��    � ; 	�*R��A�?A��_�|,�<>E�B�8���2��C�T0 k� ��
��
(%2't �1"t'%  ��    � ; 	 *R��A�?A��_�|,�<>E�B�6���2��C�T0 k� ��
��
(%2't �1"t'%  ��    � ; 	 *R��A�?A��_�|,�<?F�B�5���2��C�T0 k� ��
��
(%2't �1"t'%  ��    � ; 	)R��A�@A��_�|,�<@F�B�4���2��C�T0 k� ��
��
(%2't �1"t'%  ��    � ; 	*R��A�@A��_�|,�8AF�B�3���"��C�T0 k� ��
��
(%2't �1"t'%  ��    � ; 	*R��A�@A��_�|,�8BF�B�$2���"��C�T0 k� ��
��
(%2't �1"t'%  ��    � ; 	+R��A�AA��_�|,�4DF�B�,0���"���T0 k� ����(%2't �1"t'%  ��    � ; 	+R��A�AA��_�|,�0EF�B�4/���"���T0 k� ����(%2't �1"t'%  ��    � ; 	+R��A�BA��[�|,�0GFxB�8-�������T0 k� ����(%2't �1"t'%  ��    � ; 	,R��A�BA��[�|,�,HFtE<,�������T0 k� ����(%2't �1"t'%  ��    � ; 	,R��A�BA��[�|,�,IFpED+�������T0 k� ����(%2't �1"t'%  ��    � ; 	,R��A�CA��[�|,�(JFlEH*�������	T0 k� ����(%2't �1"t'%  ��    � ; �-R��A�CA��[�|,	t(JE�dEP)�������	T0 k� ����(%2't �1"t'%  ��    � ; �-R��A�CA��[�|,	t(KE�` EX(�������	T0 k� ����(%2't �1"t'%  ��    � ; �-R{�A�CA��[�|,	t(LE�`"E\'�������
T0 k� ����(%2't �1"t'%  ��    � ; �.Ro�A�DA��[�|,	t$ME�X%El%�������T0 k� ����(%2't �1"t'%  ��    � ; �.Rg�A�DA��[�|,	�$NE�T&Ep%�������T0 k� ����(%2't �1"t'%  ��    � ; t.R_�A�EA��[�|,	�$OE�T'Ex$���B����T0 k� ����(%2't �1"t'%  ��    � ; t.R[�A�EA��[�|,	�$OE�P)E��#���B����T0 k� ����(%2't �1"t'%  ��    � ; t/RS�A�EA��[�|,	�$PE�P*E��"���B����T0 k� ����(%2't �1"t'%  ��    � ; t/RK�A�EA��[�|,	�$PB�L+E��!���B����T0 k� ����(%2't �1"t'%  ��    � ; t/RC�A�FA��[�|,	t$QB�L,E�� ���B��ӼT0 k� ����(%2't �1"t'%  ��    � ; t0R?�A�FA��[�|,	t$QB�L.E�� ���B��ӼT0 k� ����(%2't �1"t'%  ��    � ; t0R7�A�FA��[�|,	t$QB�L/E�����B��ӼT0 k� ����(%2't �1"t'%  ��    � ; t0R/�A�FA��[�|,	t$RB�L0E�����B��ӸT0 k� ����(%2't �1"t'%  ��    � ; t0R+�A�GA��[�|,	t$RB�L1E�����B��ӸT0 k� ����(%2't �1"t'%  ��    � ; t1R#�A�GA��W�|,	�$RB�L2E�����B��ӸT0 k� ����(%2't �1"t'%  ��    � ; t 1R�A�GA��W�|,	�$RB�L3D�����B��ӸT0 k� ����(%2't �1"t'%  ��    � ; t 1R�A�GA��W�|,	�$SB�L4D�����B��ӸT0 k� ����(%2't �1"t'%  ��   � ; t 2R�A�HA��W�|,	�$SB�L6D�����R��ӸT0 k� ����(%2't �1"t'%  ��    � ; t 2R�A�HA��W�|,	�$SB�L7D�����R��ӸT0 k� ����(%2't �1"t'%  ��    � ; t 2Q��A�HA��W�|,	t$SB�P8D�����R��ӸT0 k� ����(%2't �1"t'%  ��    � ; t 2Q��A�HA��W�|,	t$SB�P9D�����R��ӸT0 k� ����(%2't �1"t'%  ��    � ; t 3Q��A�HA��W�|,	t$SB�T:D�����R��ӸT0 k� ����(%2't �1"t'%  ��    � ; t 3Q��A�IA��W�|,	t$SB�T;D�����R��ӸT0 k� ����(%2't �1"t'%  ��    � ; t$3Q��A�IA��W�|,	t$SB�T<D����R��ӸT0 k� ����(%2't �1"t'%  ��    � ; t$4Q��A�IA��W�|,$SB�X=D����R��ӸT0 k� ����(%2't �1"t'%  ��    � ; t$4Q��A�IA��W�|,$SK�X>D����R��ӸT0 k� ����(%2't �1"t'%  ��    � ; t$4Q��A�IA��W�|,$SK�\?D� ���R��ӸT0 k� ����(%2't �1"t'%  ��    � ; t$4Q��A�JA��W�|,$SK�\@D�(���RæӸT0 k� ����(%2't �1"t'%  ��    � ; t$5Q��A�JA��W�|,$SK�\@D�0���bçӸT0 k� ����(%2't �1"t'%  ��    � ; t$5Q��A�JA��W�|,$SK�`AD�8���béӸT0 k� ����(%2't �1"t'%  ��    � ; t$5Q��A�JA��W�|,$SK�`BD�@���bêӸT0 k� ����(%2't �1"t'%  ��    � ; t(5Q��A�JA��W�|,T$SK�dCD�H���bǬӸT0 k� ����(%2't �1"t'%  ��    � ; t(5Q��A�KA��W�|,T$SK�dDE�T���bǮӸT0 k� ����(%2't �1"t'%  ��    � ; t(6Q��A�KA��W�|,T$SK�dEE�\���"ǯӸT0 k� ����(%2't �1"t'%  ��    � ; t(6Q��A�KA��W�|,T$SK�hFE�d���"˱ӸT0 k� ����(%2't �1"t'%  ��    � ; �(6Q��A�KA��W�|,T$SK�hFE�l���"˳ӸT0 k� ����(%2't �1"t'%  ��    � ; �(6Q��A�KA��W�|,T$SK�hGE�t ���"˴ӸT0 k� ����(%2't �1"t'%  ��    � ; �(7Q��A�KA��W�|,T$SK�lHE�| ���"϶ӸT0 k� ����(%2't �1"t'%  ��    � ; �(7Q��A�LA��W�|,T$SK�lIE��!���"ϸӸT0 k� ����(%2't �1"t'%  ��    � ; �(7Q�A�LA��W�|,T$SK�lJE��!���"ӹӸT0 k� ����(%2't �1"t'%  ��    � ; �(7Qw�A�LA��W�|,T$SK�pJE��"���"ӻӸT0 k� ����(%2't �1"t'%  ��    � ; �,7Qo�A�LA��W�|,T$SK�pKEs�"����׽ӸT0 k� ����(%2't �1"t'%  ��    � ; �,8Qk�A�LA��W�|,T$SK�pLEs�#����ۿӸT0 k� ����(%2't �1"t'%  ��    � ; �,8Qc�A�LA��S�|,�$SK�tMEs�#������ӸT0 k� ����(%2't �1"t'%  ��    � ; �,8Q_�A�LA��S�|,�$SK�tMEs�$������ӸT0 k� ����(%2't �1"t'%  ��    � ; �,8QW�A�MA��S�|,�$SK�tNEs�$������ӸT0 k� ����(%2't �1"t'%  ��    � ; �,8QO�A�MA��S�|,�$SK�tOLS�%������ӸT0 k� ����(%2't �1"t'%  ��   � ; �,9QK�A�MA��S�|,�$SK�xOLS�&������ӸT0 k� ����(%2't �1"t'%  ��    � ; �,9QC�A�MA��S�!�,�$SK�xPLS�'������ӸT0 k� ����(%2't �1"t'%  ��    � ; �,9Q?�A�MA �S�!�,�$SK�xQLS�(������ӸT0 k� ����(%2't �1"t'%  ��    � ; �,9Q7�A�MA �S�!�,�$SK�|QLS�)������ӸT0 k� ����(%2't �1"t'%  ��    � ; �,9Q/�A�MA�S�!�,�$SK�|RLS�)s�����ӸT0 k� ����(%2't �1"t'%  ��    � ; �09Q+�A�NA�S�!�,�$SK�|SLS�*s�����ӸT0 k� ����(%2't �1"t'%  ��    � ; �0:Q#�A�NA�S�!�,�$SK�|SLS�+s����ӸT0 k� ����(%2't �1"t'%  ��    � ; �0:Q�A�NA�S�!�,�$SK��TLS�,s����ӸT0 k� ����(%2't �1"t'%  ��    � ; �0:Q�A�NA�S�!�,�$SK��ULS�,s����ӸT0 k� ����(%2't �1"t'%  ��    � ; �0:Q�A�NA�S�!�,�$SK��ULc�-s���ӸT0 k� ����(%2't �1"t'%  ��    � ; �0:Q�A�NA�S�!�,�$SK��VLc�.s���ӸT0 k� ����(%2't �1"t'%  ��    � ; �0:Q�A�NA�S�!�,�$SK��VLc�.s���ӸT0 k� ����(%2't �1"t'%  ��    � ; �0:P��A�NA�S�|,�$SK��WLc�/s���ӸT0 k� ����(%2't �1"t'%  ��    � ; �0;P��A�OA�S�|,�$SK��WLc�0s���ӸT0 k� ����(%2't �1"t'%  ��    � ; �0;P�A�OA�S�|,�$SK��XLc�0s���ӸT0 k� ����(%2't �1"t'%  ��    � ; �0;P�A�OA�S�|,�$SK��YLc�0s���ӸT0 k� ����(%2't �1"t'%  ��    � ; �4;P�A�OA�S�|,�$SK��YLd 0s���ӸT0 k� ����(%2't �1"t'%  ��    � ; �4<P߳A�OA�S�|,�$SK��ZLd 1s���ӸT0 k� ����(%2't �1"t'%  ��    � ; �4<P۳A�OA �S�|,�$SK��ZLd1C���ӸT0 k� ����(%2't �1"t'%  ��    � ; �8=PӲA�OA �S�|,�$SK��[Ld1C��#�ӸT0 k� ����(%2't �1"t'%  ��    � ; �8=PϲA�OA �S�|,4$SK��[Ld2C��'�ӸT0 k� ����(%2't �1"t'%  ��    � ; �<=PǲA�OA$�S�|,4$SK��\Ld2C��+�ӸT0 k� ����(%2't �1"t'%  ��    � ; �<>PñA�PA$�S�|,4$SK��\Ld2C���/�ӸT0 k� ����(%2't �1"t'%  ��    � ; �<>P��A�PA$�S�!�,4$SK��]Ld2C���3�ӸT0 k� ����(%2't �1"t'%  ��    � ; �@?P��A�PA(�S�!�,4$SK��]Ld3 ���3�ӸT0 k� ����(%2't �1"t'%  ��    � ; �@?P��A�PA(�S�!�,4$SK��]Ld3 ���7�ӸT0 k� ����(%2't �1"t'%  ��    � ; �@?P��A�PA(�S�!�,4$SK��^Ld3 ���;�ӸT0 k� ����(%2't �1"t'%  ��    � ; �D@P��A�PA,�S�!�,4$SK��^Ld4 ���?�ӸT0 k� ����(%2't �1"t'%  ��    � ; �D@P��A�PA,�S�!�,4$SK��_Ld4 ���C�ӸT0 k� ����(%2't �1"t'%  ��    � ; �D@P��A�PA,�S�!�,4$SK��_Ld4 c���C�ӸT0 k� ����(%2't �1"t'%  ��    � ; �HAP��A�PA0�S�!�,4$SK��`Ld4 c���G�ӸT0 k� ����(%2't �1"t'%  ��    � ; �HAP��A�PA0�S�!�,4$SK��`Ld5 c���K�ӸT0 k� ����(%2't �1"t'%  ��    � ; �HAP��A�QA0 �S�!�,4$SK��aLd5 c���K�ӸT0 k� ����(%2't �1"t'%  ��    � ; �LBP�A�QA0 �S�!�,4$SK��aLd5 c���O�ӸT0 k� ����(%2't �1"t'%  ��    � ; �LBP{�A�QA0 �S�|,D$SK��aLd 5 ����S�ӸT0 k� ����(%2't �1"t'%  ��    � ; �LBPs�A�QA4 �S�|,D$SB��bLd 6 ����T ӸT0 k� ����(%2't �1"t'%  ��    � ; �PCPo�A�QA4!�S�|,D$SB��bLd 6 ����TӸT0 k� ����(%2't �1"t'%  ��    � ; �PCPg�A�QA4!�S�|,D$SB��cLd$6 ����XӸT0 k� ����(%2't �1"t'%  ��    � ; �PCPc�A�QA4!�S�|,D$SB��cLd$6 ����\ӸT0 k� ����(%2't �1"t'%  ��    � ; �PDP[�A�QA4"�S�|,D$SB��cLd$6C���\ӸT0 k� ����(%2't �1"t'%  ��    � ; �TDPW�A�QA8"�S�|,D$SB��dLd(7C���`ӸT0 k� ����(%2't �1"t'%  ��    � ; �TDPO�A�QA8"�S�|,D$SB��dLd(7C���`ӸT0 k� ����(%2't �1"t'%  ��   � ; �TDPK�A�QA8"�S�|,D$SB��dLd(7C���dӸT0 k� ����(%2't �1"t'%  ��    � ; �XEPG�A�QA8#�S�|,D$SB��eLd,7C���h
ӸT0 k� ����(%2't �1"t'%  ��    � ; �XEP?�A�RA8#�S�|,D$SB��eLd,8C���hӸT0 k� ����(%2't �1"t'%  ��    � ; �XEP;�A�RA8#�S�|,D$SB��eLd,8C���lӸT0 k� ����(%2't �1"t'%  ��    � ; �XEP3�A�RA8$�S�|,D$SB��fLd08C���lӸT0 k� ����(%2't �1"t'%  ��    � ; �\FP/�A�RA8$�S�|,D$SB��fLd08S���pӸT0 k� ����(%2't �1"t'%  ��    � ; �\FP'�A�RA<$�S�|,D$SB��fLd08S���tӸT0 k� ����(%2't �1"t'%  ��    � ; �\FP#�A�RA<$�S�|,D$SB��gLd49S���tӸT0 k� ����(%2't �1"t'%  ��    � ; �\GP�A�RA<%�S�|,D$SB��gLT49S���xӸT0 k� ����(%2't �1"t'%  ��    � ; �`GP�A�RA<%�S�|,D$SB��gLT49S���xӸT0 k� ����(%2't �1"t'%  ��    � ; �`GP�A�RA<%�S�|,D$SB��hLT49S���xӸT0 k� ����(%2't �1"t'%  ��   � ; �`GP�A�RA<%�S�|,D$SB��hLT89S���xӸT0 k� ����(%2't �1"t'%  ��    � ; �`GP�A�RA<&�S�|,D$SB��hLT89S���|ӸT0 k� ����(%2't �1"t'%  ��    � ; �dH_��A�RA<&�S�|,D$SB��iLT8:S���|ӸT0 k� ����(%2't �1"t'%  ��    � ; �dH_��A�RA<&�S�|,D$SK��iD�<:S���|ӸT0 k� ����(%2't �1"t'%  ��    � ; �dH_�A�RA<'�S�|,D$SK��iD�<:S��ÀӸT0 k� ����(%2't �1"t'%  ��    � ; �dI_�A�SA<'�S�|,D$SK��jD�<;c��ÄӸT0 k� ����(%2't �1"t'%  ��   � ; �hI_�A�SA<'�S�|,D$SK��jD�@;c��ÄӸT0 k� ����(%2't �1"t'%  ��    � ; �hI_ߥA�SA@'�S�|,D$SK��jEt@<c��ÄӸT0 k� ����(%2't �1"t'%  ��    � ; �hI_פA�SA@(�S�|,D$SK��jEt@<c��ÈӸT0 k� ����(%2't �1"t'%  ��    � ; �hI_ӤA�SA@(�S�|,D$SK� kEt@<c��ÈӸT0 k� ����(%2't �1"t'%  ��    � ; �lJ_ϤA�SA@(�S�|,D$SK�kEt@=���ÈӸT0 k� ����(%2't �1"t'%  ��    � ; �lJ_ǤA�SA@(�S�|,D$SK�kEt@=���ÌӸT0 k� ����(%2't �1"t'%  ��    � ; �lJ_ãA�SA@)�S�|,D$SK�kEd@>���ÌӸT0 k� ����(%2't �1"t'%  ��    � ; �lK_��A�SA@)�S�|,D$SK�lEd@>���Ì ӸT0 k� ����(%2't �1"t'%  ��    � ; �pK_��A�SA@)�S�|,D$SK�lEd@?���Ð ӸT0 k� ����(%2't �1"t'%  ��    � ; �pK_��A�SA@)�S�|,D$SK�lEd@@���Ð!ӸT0 k� ����(%2't �1"t'%  ��    � ; �pL_��A�SA@*�S�|,D$SK� lEd@@���Ð"ӸT0 k� ����(%2't �1"t'%  ��    � ; �pL_��A�SA@*�S�|,D$SK�$mD4<A���Ô#ӴT0 k� ����(%2't �1"t'%  ��    � ; �tL_��A�SA@*�S�|,D$SK�(mD4<B�� Ô#ӴT0 k� ����(%2't �1"t'%  ��    � ; �tL_��A�SA@*�S�|,D$SK�,mD4<C��Ô$ӴT0 k� ����(%2't �1"t'%  ��    � ; �tM_��A�SA@+�S�|,D$SK�0mD4<C����%ӴT0 k� ����(%2't �1"t'%  ��    � ; �tM_��A�SA@+�S�|,4$SK�4nD4<C����&ӴT0 k� ����(%2't �1"t'%  ��    � ; �xM_��A�TA@+�S�|,4$TK�8nD4<C3���&ӴT0 k� ����(%2't �1"t'%  ��    � ; �xN_��A�TA@+�S�|,4 TK�<nD4<D3���'ӴT0 k� ����(%2't �1"t'%  ��    � ; �xN_�A�TA@,�S�|,4 TK�@nD48D3���(ӴT0 k� ����(%2't �1"t'%  ��    � ; �xN_{�A�TA@,�S�|,4 UK�DnD48E3���(ӴT0 k� ����(%2't �1"t'%  ��    � ; �|N_w�A�TA@,�S�|,4 UK�HoDD8E3��)ӴT0 k� ����(%2't �1"t'%  ��    � ; �|O_o�A�TA@,�S�|,4 VK�LoDD8E���*ӴT0 k� ����(%2't �1"t'%  ��    � ; �|O_k�A�TA@,�S�|,4 VK�PoDD8E���+ӴT0 k� ����(%2't �1"t'%  ��    � ; �|O_g�A�TA@-�S�|,4 VK�ToDD8F���+ӴT0 k� �� �� (%2't �1"t'%  ��    � ; �O__�A�TA@-�S�|,4 WK�ToDD4F���,ӴT0 k� �� �� (%2't �1"t'%  ��    � ; �O_[�A�TA@-�S�|,4 WK�XpDD4F��	�-ӴT0 k� �� �� (%2't �1"t'%  ��    � ; �P_W�A�TA@-�S�|,4 WK�\pDD4F��	�.ӴT0 k� ��!��!(%2't �1"t'%  ��    � ; �P_O�A�TA@.�S�|,4 WK�`pDD4F��	�/ӰT0 k� ��!��!(%2't �1"t'%  ��    � ; �P_K�A�TA@.�S�|,4 XK�dpDD4F��
�0ӰT0 k� ��!��!(%2't �1"t'%  ��    � ; �P_G�A�TA@.�S�|,4 XK�dpDD4F���1ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �Q_?�A�TA@.�S�|,4 XK�hpDD4F���2ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �Q_;�A�TA@/�S�|,4 XK�lqDT4F���3ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �Q_7�A�TA@/�S�|,4 XK�pqDT4F���4ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �Q_/�A�TA@/�S�|,4 XK�tqDT4G���5ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �Q_+�A�TA@/�S�|,4 XK�tqDT4G���6ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �R_'�A�TA@/�S�|,4 XK�xqDT4G���7ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �R_�A�TA@0�S�|,4 XK�|qD40G���8ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �R_�A�TA@0�S�|,4 XK�|rD40G����:ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �R_�A�TA@0�S�|,4 XK��rD40G����;ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �R_�A�UA@0�S�|,4 XK��rD40H����<ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �S_�A�UA@0�S�|,4 XK��rD4,H����>ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �S_�A�UA@1�S�|,4 XK��rD4,H����?ӰT0 k� ��"��"(%2't �1"t'%  ��   � ; �S_�A�UA@1�S�|,4 XK��rD4,H����@ӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �S^��A�UA@1�S�|,4 XK��sD4(H��C�BӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �S^��A�UA@1�S�|,4 XK��sD4(H��C�CӰT0 k� ��"��"(%2't �1"t'%  ��   � ; �S^�A�UA@1�S�|,4 XK��sE�$H��C�EӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^�A�UA@2�S�|,4 YK��sE�$I��C�FӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^�A�UA@2�S�|,D YK��sE�$I��C�HӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^�A�UA@2�S�|,D YK��sE�$I��	S�IӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^ߗA�UAD2�S�|,D YK��sE�$I��	S�JӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^חA�UAD2�S�|,DZK��sE�$I��	S�KӰT0 k� ��"��"(%2't �1"t'%  ��   � ; �T^ӖA�UAD2�S�|,DZK��tE�$I��	S�LӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^ϖA�UAD3�S�|,DZK��tE�$I��	S�MӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^˖A�UAD3�S�|,D[K��tE�$J��	c�NӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^ÖA�UAD3�S�|,D[K��tE�$K��	c�OӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^��A�UAD3�S�|,D[K��tD�$K��	c�OӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^��A�UAD3�S�|,D[K��tD�$K��	c�OӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^��A�UAD3�S�|,D\B��tD�$K��	c�OӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^��A�UAD4�S�|,D\B��tD�$L��	S�OӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^��A�UAD4�S�|,D]B��uD�$L��	S�PӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^��A�UAD4�S�|,D]B��uLT$M��	S�QӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �T^��A�UAD4�S�|,D^B��uLT$M��	S�QӰT0 k� ��"��"(%2't �1"t'%  ��   � ; �T^��A�VAD4�S�|,D^B��uLT$N��	S�QӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �|T^��A�VAD4�S�|,D^B��uLT$N��	c�RӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �|T^��A�VAD4�S�|,D_B��uLT$N��	c�RӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �|T^��A�VAD5�S�|,D_B��uLT$O��	c�SӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �|T^��A�VAD5�S�|,D`B��uLT$O��	c�SӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �|T^��A�VAD5�S�|,D`B��uLT$P��	c�SӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �xT^�A�VAD5�S�|,D`B��vLT$P��	S�SӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �xT^{�A�VAD5�S�|,DaB��vLT$P��	S�TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �xT^w�A�VAD5�S�|,DaB��vLd$Q� 	S�TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �xT^o�A�VAD5�S�|,DaB��vLd$Q� 	S�TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �xT^k�A�VAD5�S�|,DbB��vLd(Q� 	S�TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �tT^g�A�VAD6�S�|,DbB��vLd(R� 	c�TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �tT^c�A�VAD6�S�|,DcE��vLd(R� 	c�TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �tT^_�A�VAD6�S�|,DcE��vLd(S� 	c�TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �tT^W�A�VAD6�S�|,DcE�vLd(S�	c�TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �tT^S�A�VAD6�S�|,DdE�vLd(S�	c�TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �tT^O�A�WAD6�S�|,DdE�vLd(T���TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �pT^K�A�WAD6�S�|,DdE�wLd(T���TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �pT^G�A�WAD6�S�|,DdE�wLd(TD��T"�T0 k� ��"��"(%2't �1"t'%  ��    � ; �pT^?�A�WAD6�S�|,DeE�$wLd(UD��T"�T0 k� ��"��"(%2't �1"t'%  ��    � ; �pT^;�A�WAD7�S�|,DeE�,vLd(UD��T"�T0 k� ��"��"(%2't �1"t'%  ��   � ; �pT^7�A�WAD7�S�|,DeE�0vLd(UD��T"�T0 k� ��"��"(%2't �1"t'%  ��    � ; �pT^3�A�WAD7�S�|,DfE�8vLd(UD��T"�T0 k� ��"��"(%2't �1"t'%  ��    � ; �lT^/�A�WAD7�S�|,DfE�@vLd(VD��T"�T0 k� ��"��"(%2't �1"t'%  ��    � ; �lT^'�A�WAD7�S�|,DfE�HvLd(VD��T"�T0 k� ��"��"(%2't �1"t'%  ��    � ; �lT^#�A�WAD7�S�|,DgE�LvLd(VD��T"�T0 k� ��"��"(%2't �1"t'%  ��    � ; �lT^�A�WAD7�S�|,4gE�TuLd(WD��T"�T0 k� ��"��"(%2't �1"t'%  ��    � ; �lT^�A�WAD7�S�|,4gE�\uLd(WD ��T"�T0 k� ��"��"(%2't �1"t'%  ��    � ; �lT^�A�WAD7�S�|,4gB�dtLd(WD!��T"�T0 k� ��"��"(%2't �1"t'%  ��    � ; �lT^�A�WAD7�S�|,4hB�ltLd(WD"��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hT^�A�WAD8�S�|,4hB�tsLd(XT"��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hT^�A�WAD8�S�|,4hB�|sLd(XT#��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hT^�A�WAD8�S�|,�hB�sLd(XT$��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�WAD8�S�|,�iK��rLd(XT&��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�WAD8�S�|,�iK��rLd(YT'��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�WAD8�S�|,�iK��qLd(YT(��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]�A�XAD8�S�|,�iK��qLd(YT)��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]�A�XAD8�S�|,�iK��pLd(YT*��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]�A�XAD8�S�|,�iK��pLd(YT,��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]�A�XAD8�S�|,�iK��oLd(YT-��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]ߊA�XAD8�S�|,�iK��oLd(YT.��T"#�T0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]ۉA�XAD8�S�|,�iK��oLd(Yd.��T"#�T0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]׉A�XAD9�S�|,�hK��nLd(Yd/��T"#�T0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]ӉA�XAD9�S�|,�hK��nLd(Yd/��T"#�T0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]ˉA�XAH9�S�|,�hK��nLd(Yd0��T"#�T0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]ǈA�XAH:�S�|,�hK��nLd(Yd1��T"#�T0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]ÈA�XAH:�S�|,�hK��nLd(Yd3��T"#�T0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAL:�S�|,�hK��nLd(Yd4��T"#�T0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAL:�S�|,�hK��nLd(Yd5��T"#�T0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAL;�S�|,�hK��nLT(Yd7��T"#�T0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAP;�S�|,�hK��nLT(Yd8��T"#�T0 k� ��"��"(%2't �1"t'%  ��   � ; �hU]��A�XAP;�S�|,�hK��nLT(Yd:��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAP<�S�|,�hK��nLT(Xt;��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAT<�S�|,�hK��nLT(Xt=��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAT<�S�|,�hK��nLT(Xt>��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAT<�S�|,�hK��nD�(Xt@��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAX=�S�|,�hK��nD�(XtA��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAX=�S�|,�hK��nD�(XtC��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XAX=�S�|,�hK��nD�(Xt E��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XA\=�S�|,�hK��nD�(Xt E��TӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XA\>�S�|,�hK��nA�(X	T F��UӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]��A�XA\>�S�|,4hK��nA�(X	TF��VӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]{�A�XA\>�S�|,4hK��nA�(X	TG��VӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]w�A�YA`>�S�|,4hK��nA�(X	TH��WӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]s�A�YA`>�S�|,4hK��nA�(X	TI��WӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]o�A�YA`?�S�|,4hK��nLT(X�J��XӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]k�A�YA`?�S�|,4hK��nLT(X�J��YӰT0 k� ��"��"(%2't �1"t'%  ��    � ; �hU]g�A�YAd?�S�|,4hK��nLT(X�J��YӰT0 k� ��"��"(%2't �1"t'%  ��    � ;                                                                                                                                                                             � � �  �  �  c A�  �J����   �      � \��� ]� � � � �� T�P          �s&     T�U�    ���                � �          ]�  �  ���   8	(
         ��}z       ��Erq    ��;x�F{�    ��c   	              ?
         Ϡ      ���   @
	"           Y��          �I�     Y� �Qn     b��   
             
�� �         ��     ���    		'

           C$�         e     B�q3�    l�   	              �$          O     ���   8	
          ��           . ��    ��V ��     8     
                �q          O�     ���   X
          h  ��    B�(�     h�(�           	                ���/         ?    A  ���    0 0             h��  � �
   V�     h���                       ?	 Z �        ��     ��`   H		          o�� � �
    j �\�     o�V �_]    7��               U Z �        ��    ��` @0
            YQQ � �	    ~�&     Y:y��    X0                K	 Z �        �0�     ��`   (
"
           N��  � �	   � ��     N| �H    ��S                
	 Z          	 ���    ��`  H
w           _��       � ��     _�� ��    ��               P Z         
  ��b  �  ��@ (
          �� ��    � ���     �� ���                               �             �  ��H    0

 2                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          "�/  ��        � �?�  <� "�/ �?�  <�                      x                j  �       �                          "    ��        � �       "   �                                                               �                         �E � �� �  � ��� � �        	  
       
  0   E� ���B       �D `m@ �  u� �� l  �� l  �  l@ �� 0o� �D  p  ̄ 0p` �� p� � 0p� �$ @p� ˤ q` �� q� ބ �`� )D  k� H� d� .�  \� Ä }@ � p� -� �j� .� k� .�  k� �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ 
�\ U� 
�� V  
�| V ���� � 
�\ W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����    ;���   ������  
�fD
��L���"����D" � j  "  B   J jF�"     "�j  " ��
��
��"     
�j
�� 
  
 �
� �  �  
�     ��     � �       T    ��     �          ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  � 2( 2      �� �  ���        �; �  ���        �        ��        �        ��        �      ��     ��	��        ��                         I:  �� ��                                     �                ����              ����%��   ;  2�� �            91 Sergei Fedorov      0:01                                                                        5  5     � �KK � � � � � � � c� � �c� � � c� � �c� �		kj  � 
kr6 � ks& �kt& � kv. � kw1 �c� �c� � c� �c� �c� �cV% �c^ � c` � ca* �cb �k~ �k� �k�! � k� �k�# �	� � �	� � � � � �!� � �"B� � #B� �$K � �%K" �&"� � '"� � �(� � �)
� � �*"� � +"� �,"�	 �-*�."� � /"� � �0� � �1
� � �2"0 � �3"$ � � 4"? � � 5*M � 6*K= �7*6m � 8*Oe 9*<uH  *&mH  *&m � <*H= �  *Ce �>*4 � �  *Nl 
� �                                                                                                                                                                                                                 �� R         �    @ 
        �     Q P E a  ��                     �������������������������������������� ���������	�
��������                                                                                          ��    �1'�� ��������������������������������������������������������   �4, 6� 6 ���  I��� Q g���@w��@���@��                                                                                                                                                                                                                                                                                                                   @����                                                                                                                                                                                                                                              :    /    ��  4�J      U  	                           ������������������������������������������������������                                                                                                                                         p  ��             �          ��              	 
     ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� �������            x                 L    ,     ��  .�J      �  	                           ������������������������������������������������������                                                                                                                                         �  ��                �        � �              	     ��  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���                                                                                                                                                                                                                                                  	                                                              
        �             


             �  }�  �      ��������      v[����������������������������  R���������������������   	  '�����������������������������        '                                                                       ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" R > / 	                                � K� �t�                                                                                                                                                                                                                                                                                   
��                      e            c                  `                                                                                                                                                                                                                                                                                                                                                                                                      @ �  	(�  2�  2�  (�  F_e�  ��������E��� E�����������B����d������ށ         <  ���A :�� m          �   & AG� �  �   
              �                                                                                                                                                                                                                                                                                                                                        N K   �     
   	             !��                                                                                                                                                                                                                            Y��   �� �� �      �� :      ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� ���������  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    ;      7      "                       8     �   ���������J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p��  � ��� ��  � ��� �$ ^$     �  ��j��      1   �    >�����������J����   �    �   ����  ��   � � �N ^$  �   �                  #     �  t� ބ �� t� ބ � ��  4��4  �      �       W�������2���� g���  �     f ^�         ��  ;      W      ��F���2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                          �      �  a r!   f�"""""*��**"*�"�""�""v""*f   "  ""- ��"�"*"-""z"""""����            n   �  "  q  ��                          �  �                                 � gv"!g�vg�vggfvv|�b��r""gb"�vr�rgb��v���g���v���***�*q!q�"!a�!vwfqqr~� qw��q�~~q�����~~~�w~~w�w            �   ~   ��  ~~  �w      v    �                ggj�vvggvvgg!vg�g֪vvg�r�r��⢪rq**gjb�v�q*gjj*vv��gg�z�/�"!�"�*�""*z����qw�~q~ww��q~qwvq�w�`� ��� �w �~p w�p  ��                    �                        lggz�v��g        �       ggbvvrgggavvvqggav� �      ���w!z�w"""�!""*�"! ��        q� q�        `               �        �                      wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  " ! " ""  "!  "" "  """                                                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ "! ""! " ""  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  " ! " ""  "!  "" "  """                                                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                       �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ���� ��� ����                            �   O   T     ��                                 � ���� ��   � � �                                                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                        �          �   � � �  ��� ��  �                       �   �                      �������  ���    �        � ��                    ���� �                                                                                                                                                                                                      �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �            �  ��  �  �  ��  �                                          ���� ��� ����        ���� �                                              "  "  "                                                                                                                                                                               �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �     ��  ʘ ̪ "+�"" "" / ���                �                        ���� ��� ����                            ��  ��  ��� "  "/�����                                                                                                                                                                                  �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                � ��                    ���� �                                                                                                                                                                                                        �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �    ���                              �������  �                     �  �   �  �  ��  �  ��  �                                                                                                                                                                                                    �w
���̩ۚ,���+��   �   �   �   �  �  9  D3  D2 T2 DB DB �@ ��  ��  ��  �  "" ""�"!��" ��       �                w�  ��� ��� ��� ˼����ɀ�؊�˽ـ��˰��̰�̻@"���"+H�"$X�"$�@"E� U� E� D� ,˸  ��  ��  ,� "" �"" """�"!���� � �              �         �           �       �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                    ��   �  ��  �  �  �         � �������������  �                                                                                                                                       "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� �����                                                                                                                                                                                             ۻ� ۽� ��� H�DH�D�DP�E X�T H�P H�@ Ȥ� ̻� ˘ �� "*� �/�""/""/���                       ��  ۼ� ݻ� w�� b}ذgvz�w������ɨ�ͨ���ڋ��٭���ۻݻ� �   �          �   �   .   ."  ""  ""  ,   �   
            "  "  ""  "�   �           �   ��  �      �                                     �  �  �  ��  �  �  �  ��  �             �   �   �             � � "            � "�",�"+� ",                       "  .���"    �     �                                       �   ���                            �   �                                                                                                                 � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �                          � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                          �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �             �� ����  �       �   �   �                          �                                                                            �               �  �  ��  �   �   �       ���                                                                                                                                                                                                             �  ��� ܽи�؀  � ˚ �̹�̹�˹�˻ܻ��ܘ��܉���D���U�D�J�N T�� D�  T�  �  ��  �� �� ,ث"���"��� ���۝� {�� ��  ��� ��(�������� ˸� ɀ  ��  ��� �̀ �̈ �� ���虎�(���"��� ��� � �/�����              �   �   �   �   �        �� ��� ��           �� �   �   �   �   �   �        ��           �  �  ��  (� "�  �       � ����� ��     �  �  �          �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""����������D��M��M""""����������""""�����ADMA����""""����DD�M�""""��������AD�DM�""""�����������A�A�""""������AD�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��M��M�������D����3333DDDD�DD�M�D�������3333DDDDD�������M�DM�D����3333DDDD��A�M�M���M�����3333DDDDMM������D��D����3333DDDDA�A�A�D��M�D�����3333DDDD�������������D������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��           	 
          
        ((((((( 
	(((( """"��������AA�A             ! " # $ % & '   ( $ % ) ! " # * ('(&(%($(#("(! (((ADA�LL��L�D����3333DDDD + , -   . / 0 1  	 2         3       4 (((((((2	10/(.(-(,(+LL����������D����3333DDDD 5 6   7   8 9 1 :   $ % ) ! " #   ; ) ! " # $ % ) (#("(!()(%($ :198(((7(6(5""""����������A������    <     = 8 0 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>108(=((( (<""""�������I�I������ L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L""""�������I��D���I�������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7�D�M�D���M������3333DDDD  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`D�M�A�����MD�����3333DDDD 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
""""�����AMAD������ w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw""""������������������ w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xwwfFfFDfFFfFffdFffff3333DDDD + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+DDFFDfFFfdFffff3333DDDD � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(�""""wwwwwwwGGD � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(�""""wwwwwwqwAqwAwA �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(�""""wwwwqwqAwAqAqAq = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=A�A�A�A��LD�����3333DDDD    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( �A�LDL�L�D�L�����3333DDDD x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx""""wwwwwwDGAD w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww""""wwwwqqDAAq  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(""""wwwwwwwGGwGGwGwGw �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((�UQUUQUUQUUQUUUDUUUUU3333DDDD ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`DEQQUUDUTEUUUU3333DDDD M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M""""������������������������ � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(�""""�������DAADAI � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(��A�AM�M�DM��M334CDDDD 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5DD����M��DM�����3333DDDD x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x""""wwwwwwDGqGq w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwwGwwDGwwwwwwww + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+ADAH�DJ�H�H�����3333DDDD � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(��H��J�AD�DH�D����3333DDDD333333333333333333333333333333333333333333333333333333333333����  
�fD
��L���"���""""�������DD������D" � j  "  B   J jF� ����
��� �����
���� ����
��� �����
��� 0 q""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �KK � � � � � � � c� � �c� � � c� � �c� �	kj. � 
kr6 � ks& �kt& � kv. � kw1 �c� �c� � c� �c� �c� �cV% �c^ � c` � ca* �cb �k~ �k� �k�! � k� �k�# �	� � �	� � � � � �!� � �"B� � #B� �$K � �%K" �&"� � '"� � �(� � �)
� � �*"� � +"� �,"�	 �-*�."� � /"� � �0� � �1
� � �2"0 � �3"$ � � 4"? � � 5*M � 6*K= �7*6m � 8*Oe 9*<uH  *&mH  *&m � <*H= �  *Ce �>*4 � �  *Nl 
� ����L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������.�O�T�U��-�O�I�I�G�X�K�R�R�O� � � � � �.�/�=�����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3����������������������������������������$���<�K�X�M�K�O��0�K�J�U�X�U�\� � � � � � �.�/�=�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������.�/�=� �� �������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�2�3� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            