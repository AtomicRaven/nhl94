GST@�                                                            \     �                                               )  �   ��                    ����e j 
 J���������������z���        �h     #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    $�j� � �$  ��
  Y                                                                               ����������������������������������       ��    =b? 0Q0 45 118  4              	 

    
               ��� �4 �  ��                 nY 
)         8:�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             $F  "1          == �����������������������������������������������������������������������������                                ��  �   �  M�   @  #   �   �                                                                                '     
)nY  "$1F    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    C�|@Lÿ�df��T��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�x@Lþ�df��T��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�t@Lþ�df��T��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�pALþ�dfΈT��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�hALþ�dfΌT��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�dALþ�dfΌS��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�`BLþ�dfΌS��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��E�XBL���dfΐS��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��E�TCL���dfΐS��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��E�LCL��NdfΐS��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��   � )��E�HCL��NdfΔS��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��E�DDL��NdfΔS��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��E�<DL��NdfΔS��e|3�@�3� o�.A���3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��E�8EL��NdfΔS>�e|3�@�3� o�.A���3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��E�0EL��NdfΘS>�e|3�@�3� o�.A���3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��E�,FL���dfΘS>�e|3�@�3� o�.A���3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��E�$GK����dfΘS>�e|3�@�3� o�.A���3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��D? GK����dfΜS>�e|3�@�3� o�.A���3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��D?HK����dfΜS>�e|3�@�3� o�.A���3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��D?IK����dfΜS>�e|3�@�3� o�.A��3��SX? ��T0 k� �h	�l	U2d  �TT2q'  ��    � )��D?IK����dfΜS>�e|3�@�3� o�.A��3��SX? ��T0 k� �h
�l
U2d  �TT2q'  ��    � )��D?JK����dfΠS>�e|3�@�3� o�.A��3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I� JA���dfΠS>�e|3�@�3� o�.A��3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��KA���dfΠS>�e|3�@�3� o�.A��3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��KA���dfΠS>�e|3�@�3� o�.A��3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��KA���dfΤS>�e|3�@�3� o�/A��3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA���deΤR>�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA���deΤRN�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��   � )��I��LA���deΤRN�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA���deΨRN�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA���ddΤSN�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA���hdΤSN�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA���hdΤSN�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA���hdΤSN�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA���hdΤSN�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA��~hdΤSN�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA��~hdΠSN�e|3�@�3� o|/A��"���SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA��~hdΠSN�e|3�@�3� o|/A��3��SX? ��T0 k� �h�lU2d  �TT2q'  ��    � )��I��LA��~hdΠTN�e|3�@�3� o|/A��3��SX? ��T0 k� �h�lU2d  �TT2q'  ��   � )��I��LA��~hdΠTN�e|3�@�3� o|/A��3��SX? ��T0 k� �h �l U2d  �TT2q'  ��    � )��I��LA��~hdΠTN�e|3�@�3� o|/A��3��SX? ��T0 k� �h!�l!U2d  �TT2q'  ��   � )��I��LA��~hdΠTN�e|3�@�3� o|/A��3��SX? ��T0 k� �h#�l#U2d  �TT2q'  ��    � )��A��LA��~hcΜTN�e|3�@�3� o|/A��3��SX? ��T0 k� �h$�l$U2d  �TT2q'  ��    � )��A��LA��~hcΜTN�e|3�@�3� o|/A��3��SX? ��T0 k� �h%�l%U2d  �TT2q'  ��    � )��A��LA��~hc��TN�e|3�@�3� o|/A��3��SX? ��T0 k� �h&�l&U2d  �TT2q'  ��    � )��A��MA���hc��TN�e|3�@�3� o|/A��3��SX? ��T0 k� �h'�l'U2d  �TT2q'  ��    � )��A��MA���hc��UN�e|3�@�3� o|/A��3��SX? ��T0 k� �h(�l(U2d  �TT2q'  ��    � )��D>�MA���hc��UN�e|3�@�/� o|/A��3��SX? ��T0 k� �h)�l)U2d  �TT2q'  ��    � )��D>�MA���hc��UN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h*�l*U2d  �TT2q'  ��    � )��D>�MA���hc��UN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h,�l,U2d  �TT2q'  ��    � )��D>�NA���hc��UN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h-�l-U2d  �TT2q'  ��    � )��D>�NA���hc��UN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h.�l.U2d  �TT2q'  ��    � )��D>�NA���hc��UN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h/�l/U2d  �TT2q'  ��    � )��D>�OA���hc��VN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h0�l0U2d  �TT2q'  ��    � )��D>�OA��~hc��VN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h1�l1U2d  �TT2q'  ��    � )��DN�OA��~hc��VN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h2�l2U2d  �TT2q'  ��    � )��DN�OA��~hc��VN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h3�l3U2d  �TT2q'  ��    � )��DN�OA��~hc��VN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h5�l5U2d  �TT2q'  ��    � )��DN�OA��~hc��VN�e|3�@�/� o|/A��"s��SX? ��T0 k� �h6�l6U2d  �TT2q'  ��    � )��DN�OA��~hc��VN�e|3�@�/� o|/A��3��SX? ��T0 k� �h7�l7U2d  �TT2q'  ��    � )��DN�OA��~hc��VN�e|3�@�/� o|/A��3��SX? ��T0 k� �h8�l8U2d  �TT2q'  ��    � )��DN�OA��~hc��VN�e|3�@�/� o|/A��3��SX? ��T0 k� �h9�l9U2d  �TT2q'  ��    � )��DN�OA��~hc��VN�e|3�@�/� o|/A��3��SX? ��T0 k� �h:�l:U2d  �TT2q'  ��    � )��A��OA��~hc��WN�e|3�@�/� o|/A��3��SX? ��T0 k� �h;�l;U2d  �TT2q'  ��    � )��A��OA��Nhc��WN�e|3�@�/� o|/A��3��SX? ��T0 k� �h<�l<U2d  �TT2q'  ��    � )��A��OA��Nhc��WN�e|3�@�/� o|/A��3��SX? ��T0 k� �h=�l=U2d  �TT2q'  ��    � )��A��OA��Nhc��WN�e|3�@�/� o|/A��3��SX? ��T0 k� �h>�l>U2d  �TT2q'  ��    � )��A��OA��Nhc��WN�e|3�@�/� o|/A��3��SX? ��T0 k� �h@�l@U2d  �TT2q'  ��    � )��D>�OA��Nhc��W>�e|3�@�/� o|/A��3��SX? ��T0 k� �hA�lAU2d  �TT2q'  ��    � )��D>�PA���hc��W>�e|3�@�/� o|0A��3��SX? ��T0 k� �hB�lBU2d  �TT2q'  ��    � )��D>�PA���hc��W>�e|3�@�/� o|0A��3��SX? ��T0 k� �hC�lCU2d  �TT2q'  ��    � )��D>�PA���hc��W>�e|3�@�/� o|0A��3��SX? ��T0 k� �hD�lDU2d  �TT2q'  ��    � )��D>�PA���hcΔW>�e|3�@�/� o|0A��3��SX? ��T0 k� �hE�lEU2d  �TT2q'  ��    � )��L>�PA���hcΔW>�e|3�@�/� o|0A��3��SX? ��T0 k� �hF�lFU2d  �TT2q'  ��    � )��L>�PA���hcΔW>�e|3�@�/� o|0A��3��SX? ��T0 k� �hG�lGU2d  �TT2q'  ��    � )��L>�QA���hcΔW>�e|3�@�/� o|0A��3��SX? ��T0 k� �hH�lHU2d  �TT2q'  ��    � )��L>�QA���hcΔW>�e|3�@�/� o|0A��3��SX? ��T0 k� �hI�lIU2d  �TT2q'  ��    � )��L>�QA���hcΔW^�e|3�@�/� o|0A��3��SX? ��T0 k� �hJ�lJU2d  �TT2q'  ��    � )��L>�QA���hcΔW^�e|3�@�/� o|0A��3��SX? ��T0 k� �lK�pKU2d  �TT2q'  ��    � )��L>�QA���hcΔW^�e|3�@�/� o|0A��3��SX? ��T0 k� �lL�pLU2d  �TT2q'  ��    � )��L>�QA���hcΔW^�e|3�@�/� o|0A��3��SX? ��T0 k� �lM�pMU2d  �TT2q'  ��    � )��L>�QA���hcΔW^�e|3�@�/� o|0A��3��SX? ��T0 k� �lM�pMU2d  �TT2q'  ��    � )��L>�QA���lcΔW^�e|3�@�/� o|0A��3��SX? ��T0 k� �lN�pNU2d  �TT2q'  ��    � )��L>�QA���lcΔW^�e!�3�@�/� o|0A��3��SX? ��T0 k� �lO�pOU2d  �TT2q'  ��    � )��L>�QA���lcΔW^�e!�3�@�/� o|0A��3��SX? ��T0 k� �lP�pPU2d  �TT2q'  ��    � )��L>�RA��NlcΔV^�e!�3�@�/� o|0A��3��SX? ��T0 k� �pQ�tQU2d  �TT2q'  ��    � )��LN�RA��NlcΔV^�e!�3�@�/� o|0A��3��SX? ��T0 k� �pR�tRU2d  �TT2q'  ��    � )��LN�RA��NlcΔV^�e!�3�@�/� o|0A��3��SX? ��T0 k� �pS�tSU2d  �TT2q'  ��    � )��LN�RA��NlcΔV^�e!�3�@�/� o|0A��3��SX? ��T0 k� �pT�tTU2d  �TT2q'  ��    � )��LN�RA��NlcΔV^�e!�3�@�/� o|0A��3��SX? ��T0 k� �pT�tTU2d  �TT2q'  ��    � )��LN�RA��NlcΔV^�e!�3�@�/� o|0A��3��SX? ��T0 k� �tU�xUU2d  �TT2q'  ��    � )��LN�RA���lcΔV^�e!�3�@�/� o|0A��3��SX? ��T0 k� �tV�xVU2d  �TT2q'  ��    � )��LN�RA���lcΔV^�e!�3�@�/� o|0A��3��SX? ��T0 k� �tW�xWU2d  �TT2q'  ��    � )��LN�RA���lcΔV^�e!�3�@�/� o|0A��3��SX? ��T0 k� �tW�xWU2d  �TT2q'  ��    � )��LN�RA���lcΔV^�e|3�@�/� o|0A��3��SX? ��T0 k� �xX�|XU2d  �TT2q'  ��    � )��LN�RA���lcΔV^�e|3�@�/� o|0A��3��SX? ��T0 k� �xY�|YU2d  �TT2q'  ��    � )��B�`Er�3���C� |3�Id0	#?�E�#��<ÈT0 k� è:��:U2d  �TT2q' ��    �  �B�`Er�4���K�|3�Il0	C�E�$��D	ÌT0 k� ä:��:U2d  �TT2q' ��    �  �B��`Er�5���S�|3�Ix0	G�E�$��L	ÐT0 k� Ü;��;U2d  �TT2q' ��    �  �B��_Er�5r��[�|3�E��0	G�E�%��T
ÔT0 k� Ә;��;U2d  �TT2q' ��    �  �B��_Er�7r��k�(|3�E��1	O�F�&��dØT0 k� Ӕ>��>U2d  �TT2q' ��    �  �B��^Er�9r��s�0!�3�E��1	#S�F�'lÜT0 k� Ӥ@��@U2d  �TT2q' ��    �  �B��^Er�:r��{�8!�3�E��1	#W�F�'tӠT0 k� ӰA��AU2d  �TT2q' ��    �  B��]Er�;�����@!�3�E��1	#W�F�( |ӠT0 k� �B��BU2d  �TT2q' ��    �  B��\Er�=��	���P!�3�E��2	#[�F�) �Ӥ T0 k� ��D��DU2d  �TT2q' ��    �  E�\Er�?������X!�3�E��2	_�F�)� �Ӥ!T0 k� ��E��EU2d  �TT2q' ��    �  E�[Er�@������`!�3�E��2	c�F�*� �Ө#T0 k� ��E��EU2d  �TT2q' ��    �  E�ZEr�Ar�����h!�3�Es�2	c�F�*� �Ө$T0 k� ��G��GU2d  �TT2q' ��    �  E�ZEr�Cr�����p!�3�Es�3	c�F�*� �Ө&T0 k� ��H��HU2d  �TT2q' ��    �  E�,XEr�Fr������!�3�Es�4	#g�F�+� �Ө(T0 k� � I�IU2d  �TT2q' ��    �  E�4XD��Gr������|3�Es�4	#k�F�+� �Ө*T0 k� �J�JU2d  �TT2q' ��    �  E�<WD��Ir�����|3�Et 5	#k�F�+� �Ө+T0 k� J�JU2d  �TT2q' ��    �  E�DVD��Jr�����|3�Et5	#k�F�+� �Ө,T0 k� K�KU2d  �TT2q' ��    �  E�LUD��Lr� ����|3�Et6	#o�F�+� ��.T0 k�  L�$LU2d  �TT2q' ��    �  E�\TEb�Os�����|3�Et8	o�F�,� ���0T0 k� ,M�0MU2d  �TT2q' ��    �  E�`SEb�Qs�����|3�Et$9	o�F�,� ���1T0 k� �4N�8NU2d  �TT2q' ��    �  E�hREb�Rc�����|3�Et,9	o�F�,� ���2T0 k� �<O�@OU2d  �TT2q'  ��    �  E�pQEb�Tc����|3�Ed4:	o�@�,� ���3T0 k� �4N�8NU2d  �TT2q'  ��    �  E�xPEb�Vc����|3�Ed<;	o�@�,� ��4T0 k� �,N�0NU2d  �TT2q'  .�    �  E��NEb�Yc����|3�EdH=	#o�@�,� ��6T0 k� �4O�8OU2d  �TT2q'  ��    �  E��LEb�[c�#���|3�EdL?	#o�@�,� ��6T0 k� 0O�4OU2d  �TT2q'  ��    �  E��KEb�]c�+���|3�EdT@	#o�@�,� �$�7T0 k� 4P�8PU2d  �TT2q'  ��    �  E��JEb�_c�3�� |3�EdXA	#o�@b�,� �( �8T0 k� 4Q�8QU2d  �TT2q'  ��    �  E��IEb�`c�;��|3�Ed`B	#o�@b�,� �0!�8T0 k� 8R�<RU2d  �TT2q'  ��    �  E��IER�bc�C��|3�EddC co�@b�,� �8"�8T0 k� 8S�<SU2d  �TT2q'  ��    �  E��HER�fc#�S�� |3�EdlF co�@b�,� �H$��8T0 k� �@U�DUU2d  �TT2q'  ��    �  EøHER�gS#�W��(|3�EdpG co�@b�,� �P%��8T0 k� �DV�HVU2d  �TT2q'  ��    �  E��GER�iS#�_��0|3�EdtH co�@��,� �T&��8T0 k� �HX�LXU2d  �TT2q'  ��    �  E��FER�kS#�g��8|3�EdxI �o�@��,� �\'��7T0 k� �LY�PYU2d  �TT2q'  ��    �  E��DER�lS#�o��@|3�Ed|K �o�@��,� �d(��7T0 k� �PZ�TZU2d  �TT2q'  ��    �  E��BER�nS#�/w��H|3�A��L �o�@��,� �h)��7T0 k� �T[�X[U2d  �TT2q'  ��    �  C��@ER�oS#�/��T|3�A��N �o�@��,� �h)��7T0 k� �X[�\[U2d  �TT2q'  ��    �   C��=ER�sS�/���d|3�A��Po�@��,� �l(��7T0 k� �\]�`]U2d  �TT2q'  ��    � ! C��;P��tS�/���l|3�A��Ro�A�,� �l(��7T0 k� �`_�d_U2d  �TT2q'  ��    � " C��9P��vS�/���t|3�A��So�A�,� �l(��7T0 k� �d`�h`U2d  �TT2q'  ��    � # �C��7P��wS�/���||3�A��Uo�A�+� �l(��7T0 k� �`a�daU2d  �TT2q'  ��    � $ �C��6P��yS�/����|3�A��Vo�A�+� �l(��8T0 k� �\c�`cU2d  �TT2q'  ��    � % �C��4P��zC�/����|3�A��W�o�A�+� �l(��8T0 k� �\d�`dU2d  �TT2q'  ��    � & �C��2P��{C�/��Д|3�A��X�o�C��+� 3l(��8T0 k� �Xe�\eU2d  �TT2q'  ��    � ' �C��1P��}C�/��М|3�A��Y�o�C��+� 3p(��8T0 k� �Tf�XfU2d  �TT2q'  ��    � ( �C��.P�̀C����Ь|3�A�x\�k�C��*� 3p(��9T0 k� �Li�PiU2d  �TT2q'  �� 
   � ) �C��,P��C����д|3�A�x]�k�C��*� 3p(��8T0 k� �Hj�LjU2d  �TT2q'  �� 
   � * �C��*P���������|3�A�t^�k�C��*� 3p(��8T0 k� �Dk�HkU2d  �TT2q'  �� 
   � + �C��)P���������|3�A�p`�g�C��)� Cp'��8T0 k� �@m�DmU2d  �TT2q'  �� 
   � , �C��'P��~�������|3�A�la�g�C��)� Cp(��8T0 k� �<n�@nU2d  �TT2q'  �� 
   � - �C��&P��~��������|3�A�hb�c�C��(� Cp(��8T0 k� �8o�<oU2d  �TT2q'  �� 
   � . �C��&P��~��������|3�ETdd�_�C��(�Cp(��8T0 k� �8k�<kU2d  �TT2q'  �� 
   � / �NC�&P��}��������|3�ET\e�_�C��'�Cp(��8T0 k� �4h�8hU2d  �TT2q'  �� 
   � 0 �NC�$P��}�������|3�ETTh�W�C��&�Cp(��8T0 k� �0h�4hU2d  �TT2q'  �� 
   � 1 �NC�#P��|������ |3�ETPi�S�C��&�Cp(��8T0 k� �,f�0fU2d  �TT2q'  �� 
   � 2 �NC�"P��|�����q|3�ETLj�O�C��%�Cp(��8T0 k� �(e�,eU2d  �TT2q'  �� 
   � 3 �NC�"EҸ|�����q|3�ETDk�O�C��%�Cp'��8T0 k� �$e�(eU2d  �TT2q'  �� 
   � 4 �NC�!EҸ|����'�q|3�ET@l�K�C��$�Cp'��8T0 k� � f�$fU2d  �TT2q'  �� 
   � 5 �NC�!EҴ{����/�q|3�Ad8n�C�C��#�Cp(��8T0 k� �h�hU2d  �TT2q'  �� 
   � 6 �NC�EҰ{����;�q,|3�Ad,p�;�C��"�Sp(��7T0 k� ��k��kU2d  �TT2q'  �� 
   � 7 �NC�E�{����C�q4|3�Ad(q�7�C��!�Sp(��7T0 k� ��m��mU2d  �TT2q'  �� 
   � 8 �NC�E�{����K�q8|3�Ad r�3�C�� �Sp(��7T0 k� ��n��nU2d  �TT2q'  �� 
   � 9 �NC�E�z����O�q@|3�ETs/�C���Sp(��7T0 k� ��m��mU2d  �TT2q'  �� 
   � : �NC�E�z����_�qP|3�ETu#�C���Sp(��7T0 k� ��o��oU2d  �TT2q'  �� 	   � ; �NC�D2�z����g�qT|3�ETw�C�|�Sp(��7T0 k� ��o��oU2d  �TT2q'  �� 	   � < �NC�D2�y����k�a\|3�ET x�C�x�Sp(��7T0 k� ��o��oU2d  �TT2q'  �� 	   � < �NC�D2�y����s�ad|3�ES�y�C�t�Sp(��7T0 k� ��p��pU2d  �TT2q'  �� 	   � < �NC�D2�y����w�ah|3�ES�z�C�p�Sp(��7T0 k� ��q��qU2d  �TT2q'  �� 	   � < �NC�D2�y�����al
|3�ES�{�C�l�cl(��7T0 k� ��r��rU2d  �TT2q'  �� 	   � < �NC�D2�y����� ax|3�EC�}��C�d�cl)��6T0 k� ��q��qU2d  �TT2q'  �� 	   � < �NC�D2�y�����a||3�EC�}�C�`�cl)��6T0 k� ��p��pU2d  �TT2q'  �� 	   � < �NC�D2�y�����a�|3�EC�~�C�\�ch)��5T0 k� ��o��oU2d  �TT2q'  �� 	   � < �NC�D2�y�����a�|3�EC��C�X�ch)��5T0 k� ��n��nU2d  �TT2q'  �� 	   � < �NC�D2xy�w���a�|3�EC��ӯC�L�cd)��4T0 k� ��o��oU2d  �TT2q'  �� 	   � < �NC�DBty�o���a�|3�EC��˯C�H�cd*��3T0 k� ��n��nU2d  �TT2q'  �� 	   � < �E��DBpy�k���	a� |3�EC��ïC�D�cd*��3T0 k� �|m��mU2d  �TT2q'  �� 	   � < �E��DBlz�c���
Q��|3�A����C�@�c`+��2T0 k� �lm�pmU2d  �TT2q'  �� 	   � < �E��DB`z�W���Q��|3�A���C�4�s`,��1T0 k� �Tm�XmU2d  �TT2q'  �� 	   � < �E��ER\{�O���Q��|3�A|��C�0	�s\,��0T0 k� �Hl�LlU2d  �TT2q'  �� 	   � < �E��ERX{�K���Q��|3�At��C�(�s\-��/T0 k� �<l�@lU2d  �TT2q'  �� 	   � < �EӼERP{�C�����|3�Al~⓯C�$�s\.��.T0 k� �4l�8lU2d  �TT2q'  �� 	   � < �EӸERH|�3�����|3�A\~⃯C��sX/��,T0 k� �$k�(kU2d  �TT2q'  �� 	   � < �EӸER@|�/�����|3�AP}�w�C��sX0s�*T0 k� �k�kU2d  �TT2q'  �� 	   � < �EӴER<|�'�����|3�AH}�o�C�sX0s�'T0 k� �j�jU2d  �TT2q'  �� 	   � < �EӰER4}������|3�A@}�g�C� sX1s�$T0 k� �j�jU2d  �TT2q'  ��    � < �E�ER0}������|3�A8|�_�C��sX1s�"T0 k� � i�iU2d  �TT2q'  ��    � < �E�ER$}������|3�A#({�K�C��� sX2s�T0 k� ��h��hU2d  �TT2q'  ��    � < �E�
C�~�������|3�A# {�C�C��� sX2s�T0 k� ��h��hU2d  �TT2q'  ��    � < �E�
C�~�����!��|3�A#z�;�C��� sX3s�T0 k� ��g��gU2d  �TT2q'  �    � < }RS�	C�~�����"��|3�A#z�3�C����sX3s�T0 k� ��g��gU2d  �TT2q'  ��    � < zRS�C� �����%��|3�A"�y��C����sX3s�T0 k� ��f��fU2d  �TT2q'  ��    � < wRS�AQ������'��|3�A"�x��C����sX4s�T0 k� ��e��eU2d  �TT2q'  ��    � < tRS�AQ������(��|3�A"�w��C����sX4s�T0 k� ��e��eU2d  �TT2q'  ��    � < qRS�AQ������)��|3�A"�w��C����sX4s�T0 k� ��d��dU2d  �TT2q'  ��    � < oRS�AQ������+��|3�A"�v���C����sX4s�T0 k� ��c��cU2d  �TT2q'  ��    � < mRS�AQ������,��|3�A2�u��C����sX4s�T0 k� ��b��bU2d  �TT2q'  ��    � < jRc| AQ������/��|3�A2�t��C����sX4s�T0 k� ��`��`U2d  �TT2q'  ��    � < gRc{�AQ������0��|3�A2�s�ۯC���� �X4s�T0 k� ��`��`U2d  �TT2q'  ��    � < dRcw�EQ�~�����1��|3�A2�s�ϯC���� �X4s�
T0 k� ��_��_U2d  �TT2q'  ��    � < bRcs�EQ�~�����2w�|3�A2�rǯC���� �X4s�	T0 k� �x^�|^U2d  �TT2q'  ��    � < `Rco�EQ�~�����4o�|3�A2�q��C���� �X4s�T0 k� �p]�t]U2d  �TT2q'  ��    � < ^Rcg�EQ�}�����6c�|3�A2�p��C����CX4s�T0 k� �\\�`\U2d  �TT2q'  ��    � < [Rsc�EQ�}�����7[�|3�A2�o��C����CX5s�T0 k� �T[�X[U2d  �TT2q'  ��    � < YRsc�EQ�}�����8S�|3�EB�n��C����CX5s�T0 k� �PZ�TZU2d  �TT2q'  ��    � < WRs_�EQ�}�����:K�|3�EBxm��C����CX5s�T0 k� �LZ�PZU2d  �TT2q'  ��    � < URsW�EQ�|�����<;�|3�EBhl��C����CX6s� T0 k� �@X�DXU2d  �TT2q'  ��    � < RRsS�EQ||��� �=3�|3�EB`kw�C����CX7s��T0 k� �<W�@WU2d  �TT2q'  ��    � < PRsS�EQt|��� �>+�|3�EBXjo�C����CX7s��T0 k� �4V�8VU2d  �TT2q'  ��    � < NRsO�EAl|��� �?#�|3�EBPig�C����CX8s��T0 k� �,U�0UU2d  �TT2q'  ��    � < LRsG�EA\{�� �A�|3�EB@hS�C�w��CX9s��T0 k� �T� TU2d  �TT2q'  ��    � < JRsG�EAT{�{� �B�|3�EB8gK�C�o��SX:���T0 k� �S�SU2d  �TT2q'  ��    � < GRsC�EALz�s� �C�|3�EB0fC�E1o��SX:���T0 k� �R�RU2d  �TT2q'  ��    � < ERs?�EADz�s� �D��|3�E2(e;�E1g��SX;���T0 k� �Q�QU2d  �TT2q'  ��    � < CRs;�EA8y�g� �F��|3�E2c'�E1[��SX<���T0 k� � O�OU2d  �TT2q'  ��    � < ARs7�EA0y�_� �G��|3�E2b�E1W��SX<���T0 k� ��N� NU2d  �TT2q'  ��    � < ?Rs3�EA(y�[��H��|3�E2a�E1O��SX=c��T0 k� ��M��MU2d  �TT2q'  ��    � < =Rs3�EA x�S��I��|3�E2`�E1K��SX=c��T0 k� ��L��LU2d  �TT2q'  ��    � < ;Rs/�EAx�O��JP��|3�E1�_��E1K��SX=c��T0 k� ��K��KU2d  �TT2q'  ��    � < 9Rs+�EAw�?��LP��|3�E1�\��CAK��SX>c��T0 k� ��H��HU2d  �TT2q'  ��    � < 7Rs'�E1 v�;��xMP��|3�@��[��CAG�"C�cX>c��T0 k� ��F��FU2d  �TT2q'  ��    � < 5Rs#�E0�u�3��pNP��|3�@��Y��CA?�"C�cX>c��T0 k� ��D��DU2d  �TT2q'  ��    � < 3Rs#�E0�u�/��lOP��|3�@��X�ׯCA;�"C�cX>c��T0 k� ��C��CU2d  �TT2q'  ��    � < 1Rs�E0�t�'��dPP��|3�@��W�ϯCA7�"C�cX>c��T0 k� ��A��AU2d  �TT2q'  ��    � < /Rs�E0�s���`PP��|3�@��U�ǯCA7�"C�cX?c��T0 k� 1�@��@U2d  �TT2q' �    � < ,Rs�E0�s���XQP��|3�G�T@��CA3�"C�cX?c��T0 k� 1�?��?U2d  �TT2q' ��    � < )Rs�E0�r���PRP�|3�G�S@��CA/�"C�cX?c��T0 k� 1�=��=U2d  �TT2q' ��    � < &Rs�E0�p���DTPk�|3�G�P@��CA#�"s� �X?S��T0 k� 1�;��;U2d  �TT2q' ��    � < #Rs�E0�o����<U@c�|3�G�O@��CA�"s� �X?S��T0 k� ��9��9U2d  �TT2q'
 ��    � <  Rs�E0�n����4U@[�|3�G�M@��CA�"s� �X?S��T0 k� ��8��8U2d  �TT2q' ��    � < Rs�E0�m����,V@S�|3�G�L@��E1�"s� �X?S��T0 k� �|7��7U2d  �TT2q' ��    � < Rs�E0�l����(W@K�|3�G�K@�E1�"s� �X?S��T0 k� �t5�x5U2d  �TT2q' ��    � < Rs�E0�k���� X@C�|3�G�J@w�E1�3�X?S��T0 k� �h4�l4U2d  �TT2q' ��    � < Rs�C@�i����X@;�|3�G�H@o�E1�3�X?S��T0 k� !`3�d3U2d  �TT2q' ��    � < Rs�C@�h����Y@3�|3�G�G@g�E1�3�X?S��T0 k� !X1�\1U2d  �TT2q' ��    � < Rs�C@�g����Z@+�|3�G!�F@[�E0��3�X?S��T0 k� !P0�T0U2d  �TT2q' ��    � < Rr��C@�f����[@#�|3�G!�E0S�E0��3�X?S��T0 k� !D/�H/U2d  �TT2q' ��    � < Rr��C@�d�����[@�|3�G!xD0K�E0��3�X?C��T0 k� !<-�@-U2d  �TT2q' ��    � < Rr��C@�c�����\0�|3�G!tC0C�E0��3�X?C��T0 k� A4,�8,U2d  �TT2q' ��    � < Rr��C@|b�����]0�|3�G!pB0;�E0��3�X?C��T0 k� A(+�,+U2d  �TT2q' ��    � <��Rr��C@t`�����]0�|3�G!lA03�E ��3�X?C��T0 k� A )�$)U2d  �TT2q' ��    � <��Rr��C@p_�����^?��|3�G!d?0+�E ��"��X?C��T0 k� A(�(U2d  �TT2q' ��    � <��Rr��C@l]���o�_?��|3�G!`>0#�E ��"��X?C��T0 k� A'�'U2d  �TT2q' ��    � <��Rr��C@d\���o�`?��|3�G!\=0�E ��"��SX?C��T0 k� !%�%U2d  �TT2q' ��    � <��Rr��C@\Y�w�o�b?��|3�G!T;0�E���"��
SX?���T0 k�  �#��#U2d  �TT2q'! ��    � <��Rr��CPXW�o�o�c?��|3�G!L:0�E���"��
SX?���T0 k�  �!��!U2d  �TT2q'" ��    � <��Rr��CPPV�g�o�c?��|3�G!H9?��E���"��	SX?���T0 k�  � �� U2d  �TT2q'# ��    � <��Rr��CPLT�_�o�d?��|3�G!D8/��E���"��	SX?���T0 k� ����U2d  �TT2q'$ ��    � <��Rr��CPHS�W��e?��|3�G!@8/�E���"��	SX?��T0 k� ����U2d  �TT2q'% ��    � <��Rr��CPDQ�O��g/��|3�G!<7/�E���"��	SX?C{�T0 k� ����U2d  �TT2q'& ��    � <��Rr��CP<O�G��h/��|3�G!86/�E���"��	SX?Cw�T0 k� ����U2d  �TT2q'' ��    � <��Rr��CP8N�?��i/��|3�G!45/۾E���3�	SX?Cs�T0 k� ����U2d  �TT2q'( ��    � <��Rr��CP4L�7��j/��|3�G!04/׿E���3�SX?Ck�T0 k� ����U2d  �TT2q') ��    � <��Rr��E�0J�/��k/��|3�G!,3/��E���3�SX?Cg�T0 k� ����U2d  �TT2q'* ��    � <��Rr��E�,I�'��l/��|3�G!(2���E���3�SX?Cc�T0 k�  ���U2d  �TT2q'+ ��    � <��Rr��E�(G���n/��|3�@�$1���E���3�SX?C_�T0 k�  ���U2d  �TT2q'+ ��    � <��Rr��E�$E���o/��|3�@� 0���E���3�SX?CW�T0 k�  ���U2d  �TT2q', ��    � ;��Rr��E� D���p/��|3�@�0���E���3�SX?CS�T0 k�  |��U2d  �TT2q'- ��    � :��Rr��E�@�����s/��|3�@�.���E���3�SX?CG�T0 k� �l�pU2d  �TT2q'/ ��    � 9��Rr��E�?�����u/�|3�@�-���E���3�SX?3C�T0 k� �`�dU2d  �TT2q'/ ��    � 8��Rr��E�=����|v{�|3�@�,���E���3�SX?3?�T0 k� �X�\U2d  �TT2q'0 ��    � 7��Rr��E�;����xxw�|3�@�,���E���3�SX?37�T0 k� �P�TU2d  �TT2q'1 ��    � 6��Rr��E�:����tys�|3�@�+���E���3�SX?33�T0 k� �D	�H	U2d  �TT2q'1 ��    � 5��Rr��E� 8����p{s�|3�@� *���E���3�SX?3/�T0 k� �<�@U2d  �TT2q'2 ��    � 4��Rr��E��6����h|o�|3�@��)���EЋ�3�SX?3+�T0 k� �4�8U2d  �TT2q'2 ��    � 3��Rr��E��5����d~�k�|3�@��)��EЃ�3�SX?3#�T0 k�  ,�0U2d  �TT2q'3 ��    � 2��Rr��E��3����`�k�|3�@��(��E��3�SX?3�T0 k�   �$U2d  �TT2q'4 ��    � 1��Rr��E��1����\��g�|3�@��'��E�{�3�SX?3�T0 k�  �U2d  �TT2q'4 ��    � 0��Rr��E��0����T��d |3�@��'��E�w�3�SX?3�T0 k�  �U2d  �TT2q'5 ��    � /��Rr��E��.���P��`|3�@��&��E�o�3�SX?C�T0 k�   � U2d  �TT2q'5 ��    � .��Rr��E��,���L�`|3�@��%��E�k�3�SX?C�T0 k� �����U2d  �TT2q'5 ��    � -��Rr��E��+ߣ�H\|3�@��%��E�g�3�SX?C�T0 k� ������U2d  �TT2q'6 ��    � ,��Rr��E��)ߟ�@X|3�@��$/��E�_�3�SX?C�T0 k� ������U2d  �TT2q'6 ��    � +��Rr��E��(ߛ�<X|3�@��#/��E�[�3�SX?B��T0 k� ������U2d  �TT2q'7 ��    � *��Rr��E��&ߓ�4~T|3�@��#/��E�W�3�SX?B��T0 k� ������U2d  �TT2q'7 ��    � )��Rr��E��$ߏ�0~�P|3�@��"/��E�O�3�SX?B��T0 k� ������U2d  �TT2q'7 �    � )��Rr��C��#_���(~�P|3�@��!/��E�K�3�SX? ���T0 k� ������U2d  �TT2q'7 �    � )��Rr��C�!_���$}�L	|3�@��!/��E�C�3�SX? ���T0 k� /�����U2d  �TT2q'8 ��    � )��Rr��C� _�� }�L
|3�@�� /��E�?�3�SX? ���T0 k� /�����U2d  �TT2q'8 ��    � )��Rr��C�_{��|�H|3�@�� /��E�7�3�SX? ���T0 k� /�����U2d  �TT2q'8 ��   � )��Rr��C�_s��|�H|3�@��/��A�3�3�SX? ���T0 k� /�����U2d  �TT2q'8 ��    � )��Rr��EO�Os��{�D|3�@��/��A�/�3�SX? ���T0 k� /�����U2d  �TT2q'8 ��    � )��Rr��EO�Ok��{�D|3�@�� o��A�+�3�SX? ���T0 k� ������U2d  �TT2q'9 ��    � )��Rr��EO�Od �z�@|3�@�� o��A�#�3�SX? ���T0 k� ������U2d  �TT2q'9 ��    � )��Rr��EO�O`�y�@|3�@�� o��A��3�SX? ���T0 k� �����U2d  �TT2q'9 ��    � )��Rr��EO�OX� y�@|3�@�� o��A��3�SX? ���T0 k� �w��{�U2d  �TT2q'9 ��    � )��Rr��EO�OT x�<|3�@�� o��A��3�SX? ���T0 k� �o��s�U2d  �TT2q'9 ��    � )��Rr��EO�OL~�w�<|3�@�� o��A��3�SX? ���T0 k� �c��g�U2d  �TT2q'9 ��    � )��Rr��EO|?H~�v�<|3�@�� o��A��3�SX? ���T0 k� �[��_�U2d  �TT2q'9 ��    � )��Rr��EOx?@~�v�<|3�@�� o��A��3�SX? ���T0 k� /S��W�U2d  �TT2q'9 ��    � )��Rr��EOp?<~�u�8|3�@�� o��A��3�SX? ���T0 k� /G��K�U2d  �TT2q'8 ��    � )��Rr��C�p?4~�t�8|3�@�� o��A���3�SX? ���T0 k� /?��C�U2d  �TT2q'8 ��    � )��Rr��C�l?,~�s�8|3�@�� o��A���3�SX? ���T0 k� /7��;�U2d  �TT2q'8 ��    � )��Rr��C�h?(~�r�8|3�@�� o��A���3�SX? ���T0 k� //��3�U2d  �TT2q'8 ��    � )��Rr��C�d? ~�q�4 |3�@�� o��A��3� SX? ���T0 k� �#��'�U2d  �TT2q'8 ��    � )��Rr��C�`�~�p�4!|3�@�� o��A��3� SX? ���T0 k� ����U2d  �TT2q'8 ��    � )��Rr��C�\�	~�n�4#|3�@�� o��A��3� SX? ���T0 k� ����U2d  �TT2q'7 ��    � )��R���C�X
�
n�m�4$|3�@�� o��A��3� SX? ���T0 k� ����U2d  �TT2q'7 ��    � )��R���C�T	�
n�l�0&|3�@�� o��A�ߙ3� SX? ���T0 k� �����U2d  �TT2q'7 ��    � )��R���C�L��n�k�0(|3�@�� o� A�ۘ3� SX? ���T0 k� ������U2d  �TT2q'6 ��    � )��R���C�H��n�j�0)|3�@�� o�A�ח3� SX? ���T0 k� ������U2d  �TT2q'6 ��    � )��R���C�D��n�i�0+|3�@�� o�A�ӗ3��SX? ���T0 k� .�����U2d  �TT2q'6 ��    � )��R���C�@��	��h�,-|3�@�� o�A�Ӗ3��SX? ���T0 k� .�����U2d  �TT2q'5 ��    � )��R���C�8��	��g�,.|3�@�� o�A�ϕ3��SX? ���T0 k� .�����U2d  �TT2q'5 ��    � )��R���C�4��	��f�(0|3�@�� o�A�˔3��SX? ���T0 k� .�����U2d  �TT2q'4 ��    � )��R���C�0��	��e�(2|3�@�� o�A�Ǔ3��SX? ���T0 k� .�����U2d  �TT2q'4 ��    � )��Ub�C�(��	��d�$4|3�@�� o�A�Ó3��SX? ���T0 k� ������U2d  �TT2q'3 ��    � )��Ub�C�$��	��c�$5|3�@�� o�A���3��SX? ���T0 k� ������U2d  �TT2q'3 ��    � )��Ub{�C�  ��	��b� 7|3�@�� o�A���3��SX? ���T0 k� ������U2d  �TT2q'2 ��    � )��Ub{�C����	��b� 9|3�@�� o�A���3��SX? ���T0 k� ������U2d  �TT2q'2 ��    � )��Ubw�C���	μa�;|3�@�� o�A���3��SX? ���T0 k� ������U2d  �TT2q'1 ��    � )��Ubw�C���	μa�<|3�@�� o�	A���3��SX? ���T0 k� ������U2d  �TT2q'0 ��    � )��Ubw�A��	��`�>|3�@�� o�	A���3��SX? ���T0 k� �����U2d  �TT2q'0 ��    � )��Ubs�A��	��`�@|3�@�� o�
A���3��SX? ���T0 k� .w��{�U2d  �TT2q'/ ��    � )��Ubs�A��ޤ	��_�B|3�@�� o�A���3��SX? ���T0 k� .o��s�U2d  �TT2q'. ��    � )��D2o�A��ޠ	��_�D|3�@�� o�A���3��SX? ���T0 k� .c��g�U2d  �TT2q'- ��    � )��D2o�A��ޜ	��^�F|3�@�� o�A���3��SX? ���T0 k� .[��_�U2d  �TT2q'- ��    � )��D2o�A��ޘ	θ^�G|3�@�� o�A���3��SX? ���T0 k� .S��W�U2d  �TT2q', ��    � )��D2k�A��ސ	θ^�I|3�@�� o�A���3��SX? ���T0 k� �K��O�U2d  �TT2q'+ ��    � )��D2g�A��ތ	θ^� K|3�@�� o�A���3��SX? ���T0 k� �?��C�U2d  �TT2q'* ��    � )��D2g�A��ވ	θ]��M|3�@�� o�A���3��SX? ���T0 k� �7��;�U2d  �TT2q') ��    � )��D2c�A��ބ	θ]��O|3�@�| o�A���3��SX? ���T0 k� �/��3�U2d  �TT2q'( ��    � )��D2c�A��ހ	��]��Q|3�@�| o�A���3��SX? ���T0 k� �#��'�U2d  �TT2q'' ��    � )��D2_�A��N|	��]��S|3�@�| o�A���3��SX? ���T0 k� ����U2d  �TT2q'& ��    � )��D2[�A��Nt	��]��S|3�@�x o�A���3��SX? ���T0 k� ����U2d  �TT2q'% ��    � )��D2[�A��Np	��^��U|3�@�x o�A���3��SX? ���T0 k� .���U2d  �TT2q'$ ��    � )��D2W�A��Nl	��^��V|3�@�x o�A���3��SX? ���T0 k� -����U2d  �TT2q'# ��    � )��DBS�A��Nh	ΰ_��W|3�@�t o�A���3��SX? ���T0 k� -�����U2d  �TT2q'" ��    � )��DBO�A��>d	ΰ_��X|3�@�t o�A���3��SX? ���T0 k� -���U2d  �TT2q'! ��    � )��DBO�A��>`	ά_��Y|3�@�t o�A��3��SX? ���T0 k� -���U2d  �TT2q'  ��    � )��DBK�A��>\	Ψ`��[|3�@�p o�A�{�3��SX? ���T0 k� �ۯ�߯U2d  �TT2q' ��    � )��DBG�A��>X	Ψ`��[|3�@�p o�A�{�3��SX? ���T0 k� �ӭ�׭U2d  �TT2q' ��    � )��DBC�A��>T	��`��\|3�@�p o�A�w�3��SX? ���T0 k� �ˬ�ϬU2d  �TT2q' ��    � )��DB?�A��>P 	��a��]|3�@�p o�A�w�3��SX? ���T0 k� ����ëU2d  �TT2q' ��    � )��DB;�A��>L!	��a��^!�3�@�l o�A�s�3��SX? ���T0 k� ������U2d  �TT2q' ��    � )��DB7�A��>H"	��a��^!�3�@�l o�A�s�3��SX? ���T0 k� ������U2d  �TT2q' ��    � )��DB3�A��>D#	��a��_!�3�@�l
 o�A�o�3��SX? ���T0 k� ������U2d  �TT2q' ��    � )��DB/�A��.D$	Μa��`!�3�@�h
 o�A�k�3��SX? ���T0 k� -�����U2d  �TT2q' ��    � )��DR+�A��.@%	Θa��`!�3�@�h
 o�A�k�3��SX? ���T0 k� -�����U2d  �TT2q' ��    � )��DR'�A��.<&	Θa��`!�3�@�h
 o�A�g�3��SX? ���T0 k� -�����U2d  �TT2q' ��    � )��DR#�A��.8(	Δa��a!�3�@�h	 o�A�g�3��SX? ���T0 k� -����U2d  �TT2q' ��   � )��DR�A��.8)	Δa��a!�3�@�d	 o�A�c�3��SX? ���T0 k� -w��{�U2d  �TT2q' ��    � )��DR�A���4*	��a>�b!�3�@�d	 o�A�c�3��SX? ���T0 k� �o��s�U2d  �TT2q' ��    � )��DR�A��4+	��a>�b!�3�@�d	 o�A�_�3��SX? ���T0 k� �c��g�U2d  �TT2q' ��    � )��DR�A{��0-	��a>�c!�3�@�d	 o�A�_�3��SX? ���T0 k� �[��_�U2d  �TT2q' ��    � )��DR�Aw��0.	��a>�c|3�@�` o�A�[�3��SX? ���T0 k� �S��W�U2d  �TT2q'
 ��    � )��DR�As��,/	��a>�d|3�@�` o�A�[�3��SX? ���T0 k� �K��O�U2d  �TT2q'	 ��    � )��DR�As��,1	Όa>�d|3�@�` o�A�[�3��SX? ���T0 k� �?��C�U2d  �TT2q' ��    � )��DQ��Ao��,2	Έa��d|3�@�` o�A�W�3��SX? ���T0 k� �7��;�U2d  �TT2q' ��    � )��Da��Ak��(3	Έa��d|3�@�` o�A�W�3��SX? ���T0 k� -/��3�U2d  �TT2q' ��    � )��Da��Ag�(5	Έa��d|3�@�\ o�A�S�3��SX? ���T0 k� -#��'�U2d  �TT2q' ��    � )��Da��Ac�(6	΄a��e|3�@�\ o�A�S�3��SX? ���T0 k� -���U2d  �TT2q'  ��    � )��Da��Ac�(8>�a��e|3�@�\ o�A�O�3��SX? ���T0 k� -���U2d  �TT2q'  ,�    � )��Da��A_�(9>�a��e|3�@�\ o�A�O�3��SX? ���T0 k� -���U2d  �TT2q'  ��    � )��Ea��A[�(;>�a��e|3�@�\ o�A�K�3��SX? ���T0 k� �����U2d  �TT2q' ��    � )��Ea��AW��(<>�a��e|3�@�X o�A�K�3��SX? ���T0 k� ������U2d  �TT2q' ��    � )��Ea��AW��(>>|a��e!�3�@�X o�A�K�3��SX? ���T0 k� ����U2d  �TT2q' ��    � )��Ea��AS��(?>|a��e!�3�@�X o�A�G�3��SX? ���T0 k� ����U2d  �TT2q' ��    � )��Ea��AO��$@>xa^�e!�3�@�X o�A�G�3��SX? ���T0 k� �ۉ�߉U2d  �TT2q' ��    � )��EQ��AO��$B>xa^�e!�3�@�X o�A�G�3��SX? ���T0 k� �ӈ�׈U2d  �TT2q' ��    � )��EQ��AK��$C>xa^�e!�3�@�T o�A�C�3��SX? ���T0 k� �ˇ�χU2d  �TT2q' ��    � )��EQ��K�G��$D>ta^�e!�3�@�T o�A�C�3��SX? ���T0 k� ,���ÅU2d  �TT2q' ��    � )��EQ��K�G��$F>ta^�e!�3�@�T o�A�?�3��SX? ���T0 k� ,�����U2d  �TT2q' ��    � )��EQ��K�C��$GNpa^�e!�3�@�T o� A�?�3��SX? ���T0 k� ,�����U2d  �TT2q' ��    � )��C��K�?��$HNpa^�e!�3�@�T o� A�?�3��SX? ���T0 k� ,�����U2d  �TT2q' ��    � )��C��K�?��$INpa^�e!�3�@�P o� A�;�3��SX? ���T0 k� ,�����U2d  �TT2q' ��    � )��C��K�;��$KNla^�e!�3�@�P o�!A�;�3��SX? ���T0 k� ����U2d  �TT2q'	 ��    � )��C��K�;��$LNla^�e|3�@�P o�!A�;�3��SX? ���T0 k� ��}��}U2d  �TT2q'	 *�    � )��C��K�7��$MNh`^�d|3�@�P o�!A�7�3��SX? ���T0 k� ��~��~U2d  �TT2q'	 ��    � )��C��K�3��$NNh`n�d|3�@�P o�!A�7�3��SX? ���T0 k� �w~�{~U2d  �TT2q'	 ��    � )��C��K�3��$ONh`n�d|3�@�P o�"A�7�3��SX? ���T0 k� �o~�s~U2d  �TT2q'	 ��    � )��C�t K�/��$PNd`n�d|3�@�P o�"A�3�3��SX? ���T0 k� <g�kU2d  �TT2q'	 ��    � )��C�lK�/��$QNd`n�d|3�@�L o�"A�3�3��SX? ���T0 k� <_�cU2d  �TT2q'	 ��    � )��C�dK�+��$RNd`n�d|3�@�L o�"A�3�3��SX? ���T0 k� <W�[U2d  �TT2q'	 ��    � )��C�\K�+��$TN``n�d|3�@�L o�#A�3�3��SX? ���T0 k� <K��O�U2d  �TT2q' ��    � )��C�XL'�� UN``n�d|3�@�L o�#A�/�3��SX? ���T0 k� <C��G�U2d  �TT2q' ��    � )��C�PL'�� VN``n�d|3�@�L o�#A�/�3��SX? ���T0 k� ,;��?�U2d  �TT2q' ��    � )��C�HL#�� WN\`n�d|3�@�L o�#A�/�3��SX? ���T0 k� ,3��7�U2d  �TT2q' ��    � )��E�@L#�� XN\`n�d|3�@�L o�$A�+�3��SX? ���T0 k� ,'��+�U2d  �TT2q' ��    � )��E�8L�� YN\`n�d|3�@�H o�$A�+�3��SX? ���T0 k� ,��#�U2d  �TT2q' ��    � )��E�0	L�� ZN\`n�d|3�@�H o�$A�+�3��SX? ���T0 k� ,���U2d  �TT2q' ��    � )��E�(
L�� ZN\`n�d|3�@�H o�$A�+�3��SX? ���T0 k� L���U2d  �TT2q' ��    � )��E� L�. ZN\`n�d|3�@�H o�$A�'�3��SX? ���T0 k� L���U2d  �TT2q' ��    � )��E�L�. ZN\`n�d|3�@�H o�%A�'�3��SX? ���T0 k� K����U2d  �TT2q' ��    � )��E�L�.[N\`n�d|3�@�H o�%A�'�3��SX? ���T0 k� K�����U2d  �TT2q' ��    � )��D1L�.\N\`n�d|3�@�H o�%A�'�3��SX? ���T0 k� K���U2d  �TT2q' ��   � )��D1L�.]N\`n�d|3�@�H o�%A�#�3��SX? ���T0 k� ����U2d  �TT2q' ��    � )��D0�L�^N\an�d|3�@�D o�&A�#�3��SX? ���T0 k� �߈��U2d  �TT2q' ��    � )��D0�L�_N\an�e|3�@�D o�&A�#�3��SX? ���T0 k� �ۉ�߉U2d  �TT2q' ��    � )��D0�L�`N\an�e|3�@�D o�&A�#�3��SX? ���T0 k� �ӊ�׊U2d  �TT2q' ��    � )��EP�L�`N\an�e|3�@�D o�&A��3��SX? ���T0 k� �ˋ�ϋU2d  �TT2q' ��    � )��EP�L�`N\an�e|3�@�D o�&A��3��SX? ���T0 k� �Ǎ�ˍU2d  �TT2q'  ��    � )��EP�L�aN\an�e|3�@�D o�&A��3��SX? ���T0 k� ����ÎU2d  �TT2q'  ��    � )��EP�L�bN\an�e|3�@�D o�'A��3��SX? ���T0 k� ������U2d  �TT2q'  ,�    � )��EP�L�cN\an�e|3�@�D o�'A��3��SX? ���T0 k� ������U2d  �TT2q'  ��   � )��L�L�cN\an�e|3�@�D o�'A��3��SX? ���T0 k� ������U2d  �TT2q'  ��    � )��L�L�dN\an�e|3�@�@ o�'A��3��SX? ���T0 k� ������U2d  �TT2q'  ��    � )��L�L�eN\an�e|3�@�@ o�'A��3��SX? ���T0 k� ������U2d  �TT2q'  ��   � )��L�L���fN\an�e|3�@�@ o�(A��3��SX? ���T0 k� ������U2d  �TT2q'  ��    � )��L�L���fN\an�e|3�@�@ o�(A��3��SX? ���T0 k� ������U2d  �TT2q'  ��    � )��L�L��� gN\an�e|3�@�@ o�(A��3��SX? ���T0 k� ������U2d  �TT2q'  ��    � )��L�L��� hN\an�e|3�@�@ o�(A��3��SX? ���T0 k� ������U2d  �TT2q'  ��   � )��L�L��� hN\an�e|3�@�@ o�(A��3��SX? ���T0 k� ������U2d  �TT2q'  ��    � )��L�L��� iN\an�e|3�@�@ o�(A��3��SX? ���T0 k� ������U2d  �TT2q'  ��    � )��L� L��� i>\an�e|3�@�@ o�)A��3��SX? ���T0 k� ������U2d  �TT2q'  ��    � )��L| L���$i>\an�e|3�@�@ o�)A��3��SX? ���T0 k� ������U2d  �TT2q'  ��    � )��Lx!L���$j>\an�e|3�@�< o�)A��3��SX? ���T0 k� ������U2d  �TT2q'  ��   � )��L p"L���$j>\an�e|3�@�< o�)A��3��SX? ���T0 k� �����U2d  �TT2q'  ��    � )��L l#L���$j>\an�e|3�@�< o�)A��3��SX? ���T0 k� �����U2d  �TT2q'  ��    � )��L d$L���(k>\an�e|3�@�< o�)A��3��SX? ���T0 k� �{���U2d  �TT2q'  ��    � )��L `$L���(k>\a^�f|3�@�< o�)A��3��SX? ���T0 k� �{���U2d  �TT2q'  ��    � )��L \%L���(k>\a^�f|3�@�< o�*A��3��SX? ���T0 k� �w��{�U2d  �TT2q'  ��   � )��L T&L���(k>\a^�f|3�@�<  o�*A��3��SX? ���T0 k� �w��{�U2d  �TT2q'  ��    � )��L P&L���(k>\a^�f|3�@�<  o�*A��3��SX? ���T0 k� �s��w�U2d  �TT2q'  ��    � )��L H'L���(l>\a^�f|3�@�<  o�*A��3��SX? ���T0 k� �s��w�U2d  �TT2q'  ��    � )��L D(L���(l>\a^�f|3�@�<  o�*A��3��SX? ���T0 k� �o��s�U2d  �TT2q'  ��    � )��L @(K����,l>\a��f|3�@�<  o�*A��3��SX? ���T0 k� �o��s�U2d  �TT2q'  ��    � )��L <)K����,l>\a��f|3�@�<  o�*A��3��SX? ���T0 k� �o��s�U2d  �TT2q'  ��    � )��L 4*K����,l�\a��f|3�@�<  o�*A��3��SX? ���T0 k� �o��s�U2d  �TT2q'  ��    � )��L 0*K����,l�\a��f|3�@�<  o�+A��3��SX? ���T0 k� �o��s�U2d  �TT2q'  ��    � )��L ,+K����,l�\`��e|3�@�8  o�+A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L  ,K����,l�\`��e|3�@�8  o�+A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L -A���0l�\`��e|3�@�8  o�+A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L .A���0l�`_��e|3�@�8  o�+A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L .A���4l�`_��e|3�@�8  o�+A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L /A���4l�`_��e|3�@�8  o�+A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L /A���8l�`^��e|3�@�8  o�,A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L 0K����<l`^��e|3�@�8  o�,A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L 0K����<l`]��e|3�@�8  o�,A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�1K����@kd\��e|3�@�8  o�,A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�1K����Dkd\��e|3�@�;� o�,A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�2K����Dkd[��e|3�@�;� o�,A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�3K����HjdZ��e|3�@�;� o�,A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�3K����LjhZ��e|3�@�;� o�,A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�4K����PjhY��e|3�@�;� o�,A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�4K���TihY��e|3�@�;� o�-A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��   � )��L/�5K���TihX��e|3�@�7� o�-A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�5K���XhhX��e|3�@�7� o�-A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�5K���\hhX��e|3�@�7� o�-A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�6L��\hhW��e|3�@�7� o�-A��3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�6L��~\hhW��e|3�@�7� o�-A���3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�7L��~\hhW��e|3�@�7� o�-A���3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�7L��~\hhV��e|3�@�7� o�-A���3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�8L��~\ghV��e|3�@�7� o�-A���3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�8L��~`g hV��e|3�@�7� o�-A���3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�9L��~`g hV��e|3�@�7� o�-A���3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L/�9L���`g hV��e|3�@�7� o�.A���3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L�9L���`g lU��e|3�@�7� o�.A���3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L�:L���`g lU��e|3�@�7� o�.A���3��SX? ���T0 k� �k��o�U2d  �TT2q'  ��    � )��L�:L���`g�lU��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��   � )��L�;L���`g�pU��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��L�;L���`g�pU��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��L�;L���`g�pU��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�<L���`g�tT��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�<L˿�`g�tT��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�=Lǿ~`f�xT��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�=Lǿ~`f�xT��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�=Lǿ~`f�|T��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�>Lǿ~df�|T��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�>Lǿ~df�|T��e|3�@�7� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�>Lǿ~df��T��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�?Lǿ~df��T��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�?Lǿ~df��T��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��C�?Lÿ~df��T��e|3�@�3� o�.A���3��SX? ��T0 k� �k��o�U2d  �TT2q'  ��    � )��                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��$^ ]�.�.� � �% R�R  � �	   ����     R������    3 ?           [ Z���         �p�    ���   8

          ���.    	   ��k�    �����k&    ����            !  Z���        �     ���   0
%           cG�           ��     cG���                    =	 Z��         �`     ���   0
 
          V#T   � �
	   ��)�     V6���2[    ���}          	 Z��          ��    ���   8          e�     
    .��K�     e���K�                    9	 Z��          �      ���   P
	         ���a  ��
      B�,'    ���a�,'                              ���z                ���   P             ��~       V ƹ    ��~ ƹ                        �         �     ��J   8	            0[         j��[�     0Xv��[�     (��                 <         �p     ��@   (
I          ���=   	     ~��$2    ������&�     3��              @         ��     ��@   P	
          ���� ��
     � ���    ���� ���                              ���b       	       �  ��@     5           ?
�   5	     � �e8     ?
� �e8                       	   �        
 �`     ��@    2         ��Y   �	   � �{    ��X� �{                        �          �      ��@   P
w

                ��      �                                                                           �                               ��        ���          ��                                                                 �                          Y|�  ��        ���a�     X�����    7                   x        ���    j  �   �   �                          Y    ��        ���       X  ��           "                                                �                         ���k������� ���� � � �������        
 	        
    ?: ��y        � �`� � a� �d  \� ɤ  ]  �� ]` �� d� )D  \� �� g` �D [� � �[� �  \����. ����< ����J ����X � A _� A$ _� 
�\ W  
�\ W� 
� W� 
�\ W� �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }`���� ����� � 
�| W����� � 
�| W����� � �� u� � @[� ʄ  \@ �� 0\� �$ @\� ˤ ]` �� ]� �� �c@ �� d@ � d` �$ d� �D d� �d d� = �`� >  a����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������� )�� Y  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    $�j � ��$  �
� �  �  
�  U    ��     � s  �   ��    ��     ��k      ��    ��     �           � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �%      ��!T ���        � � �  ��        �        ��        �        ��        �    ��    X� � i        ��                         T�) , �� �                                    �                  ���� 	           W u���%��   )����                8 Cam Neely k son v    1:13                                                                        3  2     � �
� �J� �,J� y �C1 � C) �C# � C"# � C#3 �	C$3 � 
C&+ � C'( �C.4 � C6< �J� � J�! �J�. �J�& � J� �cj  �cr tkV � � k^ �7"� �7 "� �'"� �'*� � �"� � � "� � �� � �
� �*:w? )�w? )�w? )�w#*8w/  *Gw/ %*Kw?  *Bw/  *Gw? )�wR  *JxM**8d] +*Gd]  *Et_ -*Gd_  *Et }/*<d �0*2t �1*:d � 2*Pt �3)�d � 4*&| �5**|=  *Pt � 7*Et �8"|9)�tG  *Et �;"|<)�tJ  *Et x  "R z |  "R z                                                                                                                                                                                                                         �� R         �    @ 
        �     b P E d  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��    ��3�� ��������������������������������������������������������   �4, w� 6@#��@A�@T�@� A� �0��l ������                                                                                                                                                                                                                                                                                                                    �"@]�@��A,�                                                                                                                                                                                                                                     /    #    ��  D�J    	  I!  	                           ������������������������������������������������������                                                                    	                                                                   �      �      �                �  �          	  
 	 
 	 	 ������ ���� ������ ����� ���� ������������������  ���� � ���������������������������������������������������������������� ����������������������� ������������� ��������� ��������������������� �������� ����� ������������� ������� ���������������            �            	     ,    %    ��  	f�J                                  �������������������������������������������������������                                                                                                                              	       �  �      �                 V � 0            	   	 	 ������������� �������������������������������� ������  ��� ����������������������������� ����� ��� ������������������ � �� ������������������������������������ ����������� �����  ����   � ���������� �����������������            x                                                                                                                                                                                                                                                                                                              �             


            �   }�    �                                                              N�     'w               ��������   ������������  R�����������������    ��������������������  'q  N�����������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 2 G :               	                  � ���� �\                                                                                                                                                                                                                                                                                     
)nY  "$1F                    a      a            m                                                                                                                                                                                                                                                                                                                                                                                                                      @ �  >�  <�  9#�  H#�  EZm� ��� Q��0�A �N (�0f���˖�{�˦��������������                ���B :�� H	         	 �   & AG� �   �   
              �                                                                                                                                                                                                                                                                                                                                        B L   �                        !��                                                                                                                                                                                                                            Y   �� �� ����      �� B 	     ������ ���� ������ ����� ���� ������������������  ���� � ���������������������������������������������������������������� ����������������������� ������������� ��������� ��������������������� �������� ����� ������������� ������� ���������������������������� �������������������������������� ������  ��� ����������������������������� ����� ��� ������������������ � �� ������������������������������������ ����������� �����  ����   � ���������� �����������������             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    4      6   �  X                       B     �  �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f        p���� ��  p�� 5� �� ��   �@���6 ��  �@���6 �$ ^$ �r@  �@  �r@   2   K 
�|   �    ���   ����� ��   ����� �$ ^$      z 
o� ��  z 
o� �$���  � ��� �� � ��� �$ ) �  ��)  �      �   d   .���� e����J  g���         f ^�         ��  )      .      ��$��������J���J��@  ��      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                               s   D   O   w   w   v   u   f   T   �   �              3@  DDp ��4 ��tp��wpO�tpdfwGfeTwfeWwfUFwdUFweTfp�DDp���p���@�w�p   C   D   O   D   w   u   U   U  F  d  f   f   D   �   �   �DD ���7���uP��e`O�V ffg ffG Ufw UU� FUN dFw ffp DDp ��p ��@ w�p  C4 4D@O�C���O�Dt�GVfeVfdFfdFfdUfffUfffwFff�DDD���� ���                    0   G   W   W   U   E   E   w   �   �   @    fg D� O�� �� w�}�w��}����������M���M���M��������y�                    �   �   �   �   �   �   �   �   ~   w       ���w���w���~���~�DMw�������������y�                        w���w}��wt��wt��w}M�����������   M   M   ~�  p�  p   p   p      �   �   �   �               vd  eVp ffpw�Op���w���G���M�}�                                     v   ub  ub  f   `   P               "  f  U` wfP        p   p   p   p   p   p   p   p                               C4 �y�                              f  vU`vf`D�O������p}�w�  ?�  ?�  ?�  33  3#                                      f  Ug	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  "!  "" "  """           """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """""" "!   " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  "!  "" "  """           """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                          �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                                      "  "  "           �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                       �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �                           � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                                                                                                                                                                �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���            /�      �                           �   �   �   �   �   �    �      �  �  �   �     �  � � ̂" ɭ" ��� ��� ̰  �                           �            �     �                                                                                                                                                                                   "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��                     �  �� �                         ����     �   �  �  �  ��  �   �                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��      �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                    �     �                                                                                                                                                                                               �  ��� ��� ��� �ݪ�                       �   �    �z� 
�� ������������ ˍ� ��� ���������ˉ����� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��                    ˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                                         �  ��  �� ��  ��                 �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                                  �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                    �   ��   ���  ��            �           �   �                           �                        ���� ��� ����                            �    � �  ��                  ���          ��� ���  �"  " ��"�""��"! � �  �   �   �   �                                                                                                                                  	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                                   ��                  �                        ���� ��� ����                      �  �� ��  �    � ���                                                �   ���                            �   �                                                                                                   �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                �   �   �   D   E�  U�  UO                         "  "  "           �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                          �� ̻ ��˛��  �� �˚̻���ۚ����I���䘼�^���^�٘�:�^�� ^�� D�( �) �) �) ��) ˹� ț�+��,��,����  �𫝝 ��� �ɍ ��ݨ��ډ�݊�� ��D@ �D�  J�� ݩ� ��� �ۻ �ک �ڹ�ɻ��̸���������� ����������            �   ��  ��  ��  ��  ��                                          �� ��� ��� ��  �                         �   �   �"!�����                            �  �� Ș ��  ��  �                �   �                     �                             �   �   �   �   �   �                                                                                                                                                 �   �  �  �  ��  ��  C�  U=  UJ  DZ  D  E  �4 
�: ���+��"��""� """ ""   �   �                        ɪ��ɪw̚�p�������������˻��۽��ݸ�̲-ۻ"""�""�2"�@  �C  �D  �T  D@  �   �   �   "�  "     �� �  �                                        ܰ ˻ �ݚ��w{`  g`  w                      �  �  ��"� ��� "                                  �   �                      �������  ���    �                    �   ���                       ���              �   ��  ���  � �    �                                                                                                                                      ��̻������̹�̸�ݸ�����U�X�U�U�U D�T �K ̸  �� *� "� �"�����������������                �   �   �   T   T0  C3  C3  33� 3;� ;̸ ̚  �� �
˰  �" ""�""� !���������    �             �   ��      �                    �� ������}����zvw� w
�  
�        ��� �����݋���ݻ�̻۩�̽                 �   ��   ��                            ����    
�  ��  ��  ��  �����  �   �          ��                           � ��                    ���� �                                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwwDwwAwwA""""wwwwwwqADDGG""""wwwwwwqAqwAwG""""wwwwDDtwwwww""""wwwwwqGDADGqGGqw""""wwwwwwDqGqG""""wwwwwwwwwwwwqwwqww""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUEUUEUUUUUUTDUUUU3333DDDDAEQQDUDEUTUUUU3333DDDDUETQEUADQDEUDUUUU3333DDDDUQUUDUDEUTUUUU3333DDDDEQUEQUEUEUQEUUDUUUU3333DDDDQEEDEEEDUTEUUUU3333DDDDQUUQUUQUUQUUUDUUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
� �J� �,J� y �C1 � C) �C# � C"# � C#3 �	C$3 � 
C&+ � C'( �C.4 � C6< �J� � J�! �J�. �J�& � J� �cj  �cr tkV � � k^ �7"� �7 "� �'"� �'*� � �"� � � "� � �� � �
� �*:w? )�w? )�w? )�w#*8w/  *Gw/ %*Kw?  *Bw/  *Gw? )�wR  *JxM**8d] +*Gd]  *Et_ -*Gd_  *Et }/*<d �0*2t �1*:d � 2*Pt �3)�d � 4*&| �5**|=  *Pt � 7*Et �8"|9)�tG  *Et �;"|<)�tJ  *Et x  "R z |  "R z3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.�����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�����������������������������������������#��-�G�S��8�K�K�R�_� � � � � � � � � � � �,��<�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,��<� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� ��!������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 