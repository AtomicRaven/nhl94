GST@�                                                            \     �                                               L  �   ��                    ����e ��	 J���������������z���        �h     #    z���                                d8<n    �  ?     X�����  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"     "�j��   * ��
  ��                                                                              ����������������������������������       ��    =b? 0Q0 45 118  4             	 

    
               ��� �4 �  ��                 �nY 	)         8:�����������������������������������������������������������������������������������������������������������������������������=  0b  4  11                                         �  �  �  �                  n  
)          = �����������������������������������������������������������������������������                                �   3       �   @  &   �   �                                                                                 '    	�)nY  
)n    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E 3 �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������        J�@m7�^ϴY|+�=c�^d1B�c�E��P�13� T0 k� �ߠ�㠉?�D#B(%2't   ��D   0�����    J�@m7�^׳Y|+�=c�^h2B�g�J��P�13� T0 k� ���롉?�D#B(%2't   ��D   0�����    J�@m7�^߳Y|+�=c�^l4B�o�J��P�03� T0 k� ����?�D#B(%2't   ��D   0�����    J�@m7���Y|+�=c�.l6B�s�J�#�P�03� T0 k� �������?�D#B(%2't   ��D   0�����    J�@m7���Y|+�=c�.p8B�{�J�'�P�/3� T0 k� ������?�D#B(%2't   ��D   0�����    I��@m7����Y|+�=c�.t9B��J�+�P�.3� T0 k� �����?�D#B(%2't   ��D   0�����    I��@m7����Y|+�=g�.t;Bχ�EQ/�P�.3� T0 k� �����?�D#B(%2't   ��D   0�����    I��@m7���Y|+� �g�.x=BϏ�EQ/�P�-3� T0 k� �����?�D#B(%2't   ��D   0�����    I�� @m7���Y|+� �g�.|?Bϓ�EQ3�
� -3� T0 k� �#��'��?�D#B(%2't   ��D   0���      I��!@m7���Y|+� �g�.�ABϛ�EQ7�
�,3� T0 k� �+��/��?�D#B(%2't   ��D   0���     F�"@m7���Y|+� �g���CBϣ�EQ7�
�,3� T0 k� �3��7��?�D#B(%2't   ��D   0���     F�#@m7��'�Y|+� �g���DBϫ�EQ;�
�+3� T0 k� �;��?��?�D#B(%2't   ��D   0���     F�$@m7��/�Y|+� �g���FBϳ�EA;�
�$*3� T0 k� �C��G��?�D#B(%2't   ��D   0���     F�%@m7��7�Y|+� �g���HBϷ�EA?�
�,*3� T0 k� �O��S��?�D#B(%2't   ��D   0��� 
    F&@m7��?�Y|+� �g���JBϿ�EA?�
�4)3� T0 k� �W��[��?�D#B(%2't   ��D   0���     E�'@m7��G�Y|+� �g�.�LB���EAC�
�<)3� T0 k� �_��c��?�D#B(%2't   ��D   0���     E�(@m7��O�Y|+� �g�.�NB���EAC�
�D(3� T0 k� �g��k��?�D#B(%2't   ��D   0���     E�)@m7��W�Y|+� �g�.�PB���E�C�
�L(3� T0 k� �o��s��?�D#B(%2't   ��D   0���     E�*@m7��_�Y|+� �k�.�RB���E�C�
�X'3� T0 k� �w��{��?�D#B(%2't   ��D  0���     E� +@m7��g�Y|+� �k�.�TB���E�G�
�`'3� T0 k� ������?�D#B(%2't   ��D   0���     E�$,@m7��o�Y|+� �k�.�VB���E�G�
�h&3� T0 k� �������?�D#B(%2't   ��D   0���     E�,-@m7��w�Y|+� �k�.�WB���E�G�
�p&3� T0 k� �������?�D#B(%2't   ��D   0���     E�4-@m7� �Y|+� �k��YB��E�G�
�x&3� T0 k� �������?�D#B(%2't   ��D   0���     E�8.@m7� ��Y|+� �k��[B��E�G�
�%3� T0 k� �������?�D#B(%2't   ��D   0���     E�@/@m7� ��Y|+� �k��]B��E�C�
�%3� T0 k� �������?�D#B(%2't   ��D   0���      E�H0@m7� ��Y|/� �k��_B��E�C�
�$3� T0 k� �������?�D#B(%2't   ��D   0��� "    E�P1@7� ��Y|/� �k��aB�'�E�C�
�$3� T0 k� �������?�D#B(%2't   ��D   0��� $    E�T2@7����Y|/� �k��bB�3�EAC�
�#3� T0 k� �˿�Ͽ�?�D#B(%2't   ��D   0��� &    E�\2@7����Y|/� �k��dB�;�EA?�
�#3� T0 k� �Ӿ�׾�?�D#B(%2't   ��D   0��� (    E�d3@7����Y|/� �k��fB�C�EA?�
�"3� T0 k� �۽�߽�?�D#B(%2't   ��D   0��� *    E�l4@7����Y|3� �k��gB�O�EA?�
��"3� T0 k� ���罉?�D#B(%2't   ��D   0��� ,    E�t4@7��ǮY|3� �k��iB�W�EA;�
��"3� T0 k� ���）?�D#B(%2't   ��D   0��� .    B�|5@7��ϮY|7� �o���kE�c�EA;�
��!3� T0 k� ������?�D#B(%2't   ��D   0��� 0    B��5@7��ׯY|7� �o���lE�k�EA7�
��!3� T0 k� �������?�D#B(%2't   ��D   0��� 2    B��5@7��߯Y|7� �o���nE�s�EA7�
��!3� T0 k� �����?�D#B(%2't   ��D   0��� 4    B��6@7���Y|;� �o���oE��EA3�
�� 3� T0 k� �����?�D#B(%2't   ��D   0��� 6    B��6@7���Y|;� �o�� qE���E�/�
�� 3��T0 k� �����?�D#B(%2't   ��D   0��� 8    B��6@7���Y|;� �o�rE���E�/�
��3��T0 k� �����?�D#B(%2't   ��D   0��� :    B��7@7����Y|;� �o�tE���E�+�
�3��T0 k� ���#��?�D#B(%2't   ��D   0��� ;    B��7@7����Y|;� �o�uE���E�'�
�3��T0 k� �'��+��?�D#B(%2't   ��D   0��� <    C�7@7���Y|;� �o�wDЯ�E�#�
�3��T0 k� �/��3��?�D#B(%2't   ��D   0��� =    C�7@7���Y|;� �o�$xDз�E�#�
� 3��T0 k� �3��7��?�D#B(%2't   ��D   0��� >    C�7@7���Y|;� �o�(zDп�E��
�(3��T0 k� �;��?��?�D#B(%2't   ��D   0��� ?    C�7@7���Y|;� �o�0{D���E��
�03��T0 k� �?��C��?�D#B(%2't   ��D   0��� @    C�7@7���Y|;� �o�8|D���E��
�83��T0 k� �G��K��?�D#B(%2't   ��D   0��� A    C�7@7��'�Y|;� �o��@~E���E��
�D3��T0 k� �O��S��?�D#B(%2't   ��D   0��� B    C�6@7��+�Y|;� �o��DE���EQ�
�L3��T0 k� �S��W��?�D#B(%2't   ��D   0��� C    C�6@7��3�Y|;� �o��L�E���EQ��T3��T0 k� �[��_��?�D#B(%2't   ��D   0��� D    C�6@7��7�Y|;� �o��T�E���EQ��\3��T0 k� �_��c��?�D#B(%2't   ��D   0��� E    C 6@7��?�Y|;� �o��\E���EQ��d3��T0 k� �g��k��?�D#B(%2't   ��D   0��� F    C 5@7��C�Y|;� �s��`E���EQ��l3��T0 k� �k��o��?�D#B(%2't   ��D   0��� G    C5@7��K�Y|;� �s��hEp��E@���x3��T0 k� �o��s��?�D#B(%2't   ��D   0��� H    C 4@7��O�Y|;� �s��p~Ep��E@��3��T0 k� �w��{��?�D#B(%2't   ��D   0��� I    C(4@7��S�Y|;� �s��x~Eq�E@��3��T0 k� �{����?�D#B(%2't   ��D   0��� J    C03@7��[�Y|;� �s�߀}Eq�E@��
��3��T0 k� �������?�D#B(%2't   ��D   0��� K    C83@7��_�Y|;� �s�߈}Eq�E@��
��3��T0 k� �������?�D#B(%2't   ��D   0��� L    E�@2@7��c�Y|;� �s�ߐ|Eq�C@��
��3��T0 k� �������?�D#B(%2't   ��D   0��� M    E�L2@7��g�Y|;� �s�ߔ|Eq�C@��
��3��T0 k� �������?�D#B(%2't  �D   0��� S    E�T1@7��o�Y|;� �s��{Eq�C@��
��3��T0 k� �������?�D#B(%2't  ��O   0��� Y    E�\1@7��s�Y|;� �s��zEq�C@��
��3��T0 k� �������?�D#B(%2't  �O    ��� Y    E�d0@7��w�Y|;� �s��zEq�C@����3��T0 k� �����?�D#B(%2't  �O    ��� Y    E�l0@7��{�Y|;� �s��yEq#�E0����3��T0 k� �����É?�D#B(%2't  ��O    ��� Y    E�t/@7����Y|;� �s��xEq'�E0����3��T0 k� �����ĉ?�D#B(%2't  ��O    ��� Y    E�|/@7����Y|;� �s���xEq'�E0����3��T0 k� �����ŉ?�D#B(%2't  ��O    ��� Y    @`�.@7����Y|;� �s���wEq+�E0����3��T0 k� �����Ɖ?�D#B(%2't  ��O    ��� Y    @`�.@7����Y|;� �s���vEq/�E0����3��T0 k� ���ǉ?�D#B(%2't  ��O    ��� Y    @`�-@7����Y|;� �s���uEq/�E ����3��T0 k� ���ȉ?�D#B(%2't 	 ��O    ��� Y    @`�-@7����Y|;� �s���tEq3�E ����3��T0 k� �'��+ɉ?�D#B(%2't 
 ��O    ��� Y    @`�,@7����Y|;� �s���sEq7�E ����3��T0 k� �3��7ɉ?�D#B(%2't  ��O    ��� Y    @`�,@7����Y|;� �s���sEq7�E ��� 3��T0 k� �C��Gʉ?�D#B(%2't  ��O    ��� Y    @`�+@7����Y|;� �s��rEq7�E ���3��T0 k� �O��Sˉ?�D#B(%2't  ��O    ��� Y    @`�+@7����Y|;� �s�pqEq;�B����3��T0 k� �_��c̉?�D#B(%2't  ��O    ��� Y    @`�*@7����Y|;� �s�ppEq;�B����3��T0 k� �k��o͉?�D#B(%2't  ��O    ��� Y    @`�*@7����Y|;� �s�pnEq?�B����3��T0 k� �{��Ή?�D#B(%2't  ��O    ��� Y    @`�)@7����Y|;� �w�pmEq?�B����3��T0 k� �����ω?�D#B(%2't  ��O    ��� Y    @`�)@7����Y|;� �w�p lEq?�B����3��T0 k� �����Љ?�D#B(%2't  ��O    ��� Y    @`�(@7����Y|;� �w�p(kEq?�B����
3��T0 k� �����щ?�D#B(%2't  ��O    ��� Y    @`�(@7����Y|;� �w�p0jEq?�B���� 	3��T0 k� �����҉?�D#B(%2't  ��O    ��� Y    @`�(@7��óY|;� �w�p4iEq?�B����$3��T0 k� �����҉?�D#B(%2't  ��O    ��� Y    @`�'@7��ǳY|;� �w�p<gEqC�B����(3��T0 k� �����Ӊ?�D#B(%2't  ��O    ��� Y    @`�'@7��˳Y|;� �w��DfEqC�B���3,3��T0 k� �����ԉ?�D#B(%2't  ��O    ��� Y    @`�&@7��ϳY|;� �w��LeEqC�B���3,3��T0 k� �����Չ?�D#B(%2't  ��O    ��� Y    @a &@7��ϳY|;� �w��PcBAC�C ��303��T0 k� �����։?�D#B(%2't  ��O    ��� Y    @a&@7��ӳY|;� �w��XbBAC�C ��343��T0 k� ���׉?�D#B(%2't  ��O    ��� Y    @a%@7��׳Y|;� �w��\aBAC�C ��343��T0 k� ���؉?�D#B(%2't  ��O    ��� Y    @a%@7��۳Y|;� �w�Pd_BAC�C ��383��T0 k� �#��'ى?�D#B(%2't  ��O    ��� Y    @a$@7��ߴY|;� �w�Ph^BAC�C ��3<3��T0 k� �3��7ډ?�D#B(%2't  ��O    ��� Y    @a$@7���a�;� �w�Pp]BAC�C ��3@"���T0 k� �?��Cۉ?�D#B(%2't  ��O    ��� Y    @a $@7���a�;� �w�Pt\@C�C ��3@ "���T0 k� �O��Sۉ?�D#B(%2't  ��O    ��� Y    @a$#@7���a�;� �w�P|Z@C�C ��3G�"���T0 k� �[��_܉?�D#B(%2't  ��O    ��� Y    @a,#@7���a�;� �w�P�Y@C�C ��3G�"���T0 k� �k��o݉?�D#B(%2't  ��O    ��� Y    @a0#@7���a�;� �w�P�X@C�C ��3K�"���T0 k� �w��{މ?�D#B(%2't  ��O    ��� Y    @a4"@7����a�;� �w�P�W@C�C ��3O�"���T0 k� �����߉?�D#B(%2't  ��O    ��� Y    @a<"@7����a�;� �w�P�V@aC�C��3O�"���T0 k� �������?�D#B(%2't  ��O    ��� Y    @a@"@7����a�;� �w�P�U@aC�C��3S�"���T0 k� ������?�D#B(%2't  ��O    ��� Y    @aD!@7���a�;� �w�P�T@aC�C��CS�"���T0 k� ������?�D#B(%2't  ��O    ��� Y    @aH!@7��a�;� �w�`�R@aC�C��CW�"���T0 k� ������?�D#B(%2't  ��O    ��� Y    @aL!@7��a�;� �w�`�Q@aC�C��C[�"���T0 k� ������?�D#B(%2't  ��O    ��� Y    @aT!@7��Y|;� �w�`�P@�C�C��C[�3��T0 k� ������?�D#B(%2't  ��O    ��� Y    @aX @7��Y|;� �w�`�O@�C�C��C_�3��T0 k� ������?�D#B(%2't  ��O    ��� Y    @a\ @7��Y|;� �w�`�N@�C�C��C_�3��T0 k� ������?�D#B(%2't  ��O   ��� Y    @a` @7��Y|;� �w�`�M@�C�C��Cc�3��T0 k� ����?�D#B(%2't  ��O    ��� Y    @ad@7�#�Y|;� �w�`�L@�C�C��Cc�3��T0 k� ����?�D#B(%2't  ��O    ��� Y    @ah@7�+�Y|;� �w�`�KCAC�C��Cg�3��T0 k� �#��'�?�D#B(%2't  ��O    ��� Y    @al@7�3�Y|;� �w�`�JCAC�C ��Cg�3��T0 k� �/��3�?�D#B(%2't  ��O    ��� Y    @ap@7�7�Y|;� �w�`�ICAC�C ��Ck�3��T0 k� �?��C�?�D#B(%2't  ��O    ��� Y    @at@7�?�Y|;� �{�`�ICAC�C ��Ck�3��T0 k� �K��O�?�D#B(%2't  ��O    ��� Y    @ax@7�C�Y|;� �{�`�HCAC�C!�Co�3��T0 k� �[��_�?�D#B(%2't  ��O    ��� Y    @a|@7�K�Y|;� �{�`�GCAC�C!�Co�3��T0 k� �g��k�?�D#B(%2't  ��O    ��� Y    @a�@7�O�a�;� �{�`�FCAC�C!�Cs�"s��T0 k� �w��{�?�D#B(%2't  ��O    ��� Y    @a�@7�[�a�;� �{�`�ECAC�C!�Cs�"s��T0 k� ������?�D#B(%2't  ��O    ��� Y    @a�@7�g�a�8  �{�`�DCQC�C!�Cw�"s��T0 k� �������?�D#B(%2't  ��O    ��� Y    @a�@7��s�a�8 �{�`�CCQC�C!�Cw�"s��T0 k� ������?�D#B(%2't  ��O    ��� Y    @a�@7��{�a�8 �{�`�CCQC�C!�C{�"s��T0 k� ������?�D#B(%2't  ��O    ��� Y    @a�@7���a�8 �{�`�BCQC�C!�C{�"s��T0 k� ������?�D#B(%2't  ��O    ��� Y    @a�@7���a�8 �{�`�ACQC�K��C�"s��T0 k� ������?�D#B(%2't  ��O    ��� Y    @a�@7���a�8 �{�`�@CQC�K��C�"s��T0 k� �������?�D#B(%2't  ��O    ��� Y    @a�@7���a�8 �{�a ?CQC�K�#�C�"s��T0 k� �������?�D#B(%2't  ��O    ��� Y    @a�@7���a�8 �{�a?CQC�K�'�C��"s��T0 k� �������?�D#B(%2't  ��O    ��� Y    @a�@7���a�8 �{�a>CQC�K�+�C��"s��T0 k� �����?�D#B(%2't  ��O    ��� Y    @a�@7���Y|8 �{�a=E!C�K�+�C��3��T0 k� �����?�D#B(%2't  ��O    ��� Y    @a�@7����Y|8 �{�a<E!C�K�/�C��3��T0 k� ���#��?�D#B(%2't  ��O    ��� Y    @a�@7����Y|8 �{�a<E!C�K�3�C��3��T0 k� �+��/��?�D#B(%2't  ��O    ��� Y    @a�@7����Y|8 �{�a;E!C�K�7�C��3��T0 k� �+��/��?�D#B(%2't  ��O    ��� Y    @a�@7����Y|8 �{�a:E!C�K�7�C��3��T0 k� �;��?��?�D#B(%2't  ��O    ��� Y    @a�@7����Y|8 �{�a:E!G�K�;�C��3��T0 k� �G��K��?�D#B(%2't  ��O    ��� Y    @a�@7����Y|8 �{�a 9E!G�K�?�C��3��T0 k� �W��[��?�D#B(%2't  ��O    ��� Y    @a�@7����Y|8 �{�a 8E!K�K�?�C��3��T0 k� �c��g��?�D#B(%2't  ��O    ��� Y    @a�@7���Y|8 �{�a$8E!K�K�C�C��3��T0 k� �s��w��?�D#B(%2't  ��O    ��� Y    @a�@7���Y|8 �{�a(7E!O�K�C�C��3��T0 k� �| �� �?�D#B(%2't  ��O    ��� Y    @a�@7���Y|8 �{�a,6B�O�K�G�C��3��T0 k� �� �� �?�D#B(%2't  ��O    ��� Y    @a�@7���Y|8 �{�a,6B�O�K�K�C��3��T0 k� �����?�D#B(%2't  (�O    ��� Y    @a�@7��'�Y|8 �{�a05B�S�K�K�C��3��T0 k� 4����?�D#B(%2't  ��O    ��� Y    @a�@7��/�Y|8�{�a45B�S�K�O�C��3��T0 k� 4����?�D#B(%2't  ��O    ��� Y    @a�@7��7�Y|8�{�a84B�W�K�O�C��3��T0 k� 4����?�D#B(%2't  ��O    ��� Y    @a�@7��;�Y|8�{�a83I1W�K�S�C��3��T0 k� 4����?�D#B(%2't  ��O    ��� Y    @a�@7��C�Y|8�{�a<3I1W�K�S�3��3��T0 k� 4����?�D#B(%2't  ��O    ��� Y    @a�@7��K�Y|8�{�Q@2I1[�K�W�3��3��T0 k� �����?�D#B(%2't  ��O    ��� Y    @a�@7��S�Y|8�{�Q@2I1[�K�[�3��3��T0 k� �����?�D#B(%2't  ��O    ��� Y    @a�@7��[�Y|8�{�QD1I1[�K�[�3��3��T0 k� �|���?�D#B(%2't  ��O    ��� Y    @a�@7��_�Y|8�{�QH1IA_�K�_�3��3��T0 k� �x	�|	�?�D#B(%2't  ��O    ��� Y    @a�@7��g�Y|8�{�QH0IA_�K�_�3��3��T0 k� �t
�x
�?�D#B(%2't  ��O    ��� Y    @a�@7��o�Y|8�{�QL0IA_�K�c�3��3��T0 k� �p�t�?�D#B(%2't  ��O    ��� Y    @a�@7��s�Y|8�{��P/IA_�K�c�3��3��T0 k� �p�t�?�D#B(%2't  ��O    ��� Y    @a�@7��{�Y|8�{��P.IA_�K�g�3��3��T0 k� �l�p�?�D#B(%2't  ��O    ��� Y    @a�@7���Y|8�{��T.I1_�K�g�3��3��T0 k� �h�l�?�D#B(%2't 
 ��O    ��� Y    @a�@7� b��Y|8�{��X-I1_�K�k�3��3��T0 k� �d�h�?�D#B(%2't 	 ��O    ��� Y    @a�@7� b��Y|8�{��X,I1_�K�k�S��3��T0 k� D`�d�?�D#B(%2't 	 ��O    ��� Y    @a�@7� b��Y|8�{��\+I1_�K�k�S��3��T0 k� D\�`�?�D#B(%2't  ��O    ��� Y    @a�@7� b��Y|8�{��\+I1_�K�o�S��3��T0 k� DX�\�?�D#B(%2't  ��O    ��� Y    @a�@7� b��Y|8�{��`*IA_�K�o�S��3��T0 k� DT�X�?�D#B(%2't  ��O    ��� Y    @a�@7� b��Y|8�{��`)IA_�K�s�S��3��T0 k� DT�X�?�D#B(%2't  ��O    ��� Y    @a�@7� b��Y|8�{��d(IA_�K�s�S��3��T0 k� $P�T�?�D#B(%2't  ��O    ��� Y    @a�@7� b��Y|8�{��d'IA_�K�w�S��3��T0 k� $P�T�?�D#B(%2't  ��O    ��� Y    @a�@7� b��Y|8�{��h&IA_�K�w�S��3��T0 k� $P�T�?�D#B(%2't  ��O    ��� Y    @b @7� b��Y|8�{��l%I1_�K�w���3��T0 k� $P�T�?�D#B(%2't  ��O    ��� Y    @b @7� b��Y|8�{��l$I1_�K�{���3��T0 k� $P�T�?�D#B(%2't   ��O    ��� Y    @b@7� b��Y|8���p"I1_�K�{���3��T0 k� 4T�X�?�D#B(%2't   ,�O    ��� Y    @b@7� b��Y|8���p!I1_�K����3��T0 k� 4T�X�?�D#B(%2't   ��O    ��� Y    @b@7� b��Y|8���t I1_�K����3��T0 k� 4T�X�?�D#B(%2't  ��O    ��� Y    @b@7� b��Y|8���t@a_�K����3��T0 k� 4T�X�?�D#B(%2't  ��O    ��� Y    @b@7� b��Y|8���t@a_�K�����3��T0 k� 4X�\�?�D#B(%2't  ��O    ��� Y    @b@7� b��Y|8���x@a_�K�����3��T0 k� �X�\�?�D#B(%2't  ��O    ��� Y    @b@7� b��Y|8���x@a_�K�����3��T0 k� �X�\�?�D#B(%2't  ��O    ��� Y    @b@7� b��Y|8���|@a_�K�����3��T0 k� �X�\�?�D#B(%2't  ��O    ��� Y    @b@7� b��Y|8���|@a_�K�����3��T0 k� �X�\�?�D#B(%2't  ��O    ��� Y    @b@7� b��Y|8����@a_�K�����3��T0 k� �\�`�?�D#B(%2't  ��O    ��� Y    @b@7� b��Y|8����@a_�K����{�3��T0 k� �\ �` �?�D#B(%2't  ��O    ��� Y    @b@7� b��Y|8����@_�K����{�3��T0 k� �\!�`!�?�D#B(%2't  ��O    ��� Y    @b@7� b��Y|8����@_�K����w�3��T0 k� �\!�`!�?�D#B(%2't  ��O    ��� Y    @b@7� c�Y|8����@_�K����s�3��T0 k� �`"�d"�?�D#B(%2't  ��O    ��� Y    @b@7� c�Y|8����@_�K����o�3��T0 k� �`#�d#�?�D#B(%2't  ��O    ��� Y    @b@7� c�Y|8����@_�K���k�3��T0 k� �`$�d$�?�D#B(%2't  ��O    ��� Y    @b@7� c�Y|8 ����K�_�K���g�3��T0 k� �`%�d%�?�D#B(%2't  ��O    ��� Y    @b @7� c�Y|8 ����	K�_�K���c�3��T0 k� �`&�d&�?�D#B(%2't  ��O    ��� Y    @b @7� c�Y|8 ����K�_�K���_�3��T0 k� $d'�h'�?�D#B(%2't  ��O    ��� Y    @b @7� c Y|8 ����K�_�B�[�3��T0 k� $d'�h'�?�D#B(%2't  ��O    ��� Y    @b$@7� c Y|8 ����K�_�B�W�3��T0 k� $d(�h(�?�D#B(%2't  ��O    ��� Y    @b$@7� c Y|8 ����K�_�B�S�3��T0 k� $d)�h)�?�D#B(%2't  ��O    ��� Y    @b$@7� c$Y|8 ���� K�_�B�S�3��T0 k� $h*�l*�?�D#B(%2't  ��O    ��� Y    @b(@7� c(Y|8 �����K�_�B�O�3��T0 k� �h+�l+�?�D#B(%2't  ��O    ��� Y    @b(@7� c,Y|8 �����K�_�@���K�3��T0 k� �h,�l,�?�D#B(%2't  ��O    ��� Y    @b(@7� c0Y|8 �����K�_�@���G�3��T0 k� �h-�l-�?�D#B(%2't  ��O   ��� Y    @b,@7� c0Y|8 �����K�_�@���C�3��T0 k� �h-�l-�?�D#B(%2't  ��O    ��� Y    @b,@7� c4Y|8 �����K�_�@���#C�3��T0 k� �l.�p.�?�D#B(%2't  ��O    ��� Y    @b,@7� c8Y|8 �����K�_�@���#?�3��T0 k� �l/�p/�?�D#B(%2't  ��O    ��� Y    @b,@7� c<Y|8 �����K�_�E���#;�3��T0 k� �l0�p0�?�D#B(%2't  ��O    ��� Y    @b0@7� c@Y|8 �����K�_�E���#7�3��T0 k� $l1�p1�?�D#B(%2't  ��O    ��� Y    @b0@7� cDY|8 �����K�_�E���#7�3��T0 k� $l2�p2�?�D#B(%2't  ��O    ��� Y    @b0@7� cDY|8 �����K�_�E���#3�3��T0 k� $p3�t3�?�D#B(%2't  ��O    ��� Y    @b4@7� cHY|8 �����K�_�E���#/�3��T0 k� $p3�t3�?�D#B(%2't  ��O    ��� Y    @b4@7� cLY|8 �����K�_�AQ��#+�3��T0 k� $p4�t4�?�D#B(%2't  ��O    ��� Y    @b4@7� cPY|8 �����K�_�AQ��#+�3��T0 k� �p5�t5�?�D#B(%2't  ��O    ��� Y    @b4@7� cPY|8 ��q��K�_�AQ��#'�3��T0 k� �t6�x6�?�D#B(%2't  ��O    ��� Y    @b8@7� cTY|8 ��q��K�_�AQ��##�3��T0 k� �t7�x7�?�D#B(%2't  ��O    ��� Y    @b8@7� cX	Y|8 ��q��K�_�AQ��##�3��T0 k� �t8�x8�?�D#B(%2't  ��O    ��� Y    @b8@7� c\	Y|8 ��q��K�_�A���#�3��T0 k� �t9�x9�?�D#B(%2't   ��O    ��� Y    @b8@7� c\
Y|8 ��q��K�_�A���#�3��T0 k� �t9�x9�?�D#B(%2't   ��O   ��� Y    @b<@7� c`
Y|8 ��q��K�_�A���#�3��T0 k� �x:�|:�?�D#B(%2't   -�O    ��� Y    @b<@7� cdY|8 ��q��K�_�A���#�3��T0 k� $x;�|;�?�D#B(%2't   ��O    ��� Y    @b<@7� cdY|8 ��q��K�_�A���#�3��T0 k� $x<�|<�?�D#B(%2't   ��O    ��� Y    @b<@7� chY|8 ��q��K�_�D1��#�3��T0 k� $x=�|=�?�D#B(%2't   ��O    ��� Y    @b@@7� clY|8 ��q��K�_�D1��#�3��T0 k� $|>��>�?�D#B(%2't   ��O    ��� Y    @b@@7� clY|8 ��a��K�_�D1��#�3��T0 k� $|?��?�?�D#B(%2't   ��O    ��� Y    @b@@7� cpY|8 ��a��K�_�D1��#�3��T0 k� �|?��?�?�D#B(%2't  ��O    ��� Y    @bD@7� ctY|8 ��a��K�_�EᏐ#�3��T0 k� �|A��A�?�D#B(%2't  ��O    ��� Y    @bD@7� cxY|8��a��K�_�EᏐ#�3��T0 k� ��B��B�?�D#B(%2't  ��O    ��� Y    @bD@7� cxY|8��a��K�_�Eዑ#�3��T0 k� ��C��C�?�D#B(%2't  ��O    ��� Y    @bD@7� c|Y|8��a��K�_�Eᇒ#�3��T0 k� ��D��D�?�D#B(%2't  ��O    ��� Y    @bD@7� c�Y|8��a��K�_�Eდ"��3��T0 k� ��D��D�?�D#B(%2't  ��O    ��� Y    @bH@7� c�Y|8��a��K�_�Eე"��3��T0 k� $�E��E�?�D#B(%2't  ��O    ��� Y    @bH@7� c�Y|8��a��K�_�E��"��3��T0 k� $�F��F�?�D#B(%2't   ��O    ��� Y    @bH@7� c�Y|8��a��K�_�E�{�"��3��T0 k� $�G��G�?�D#B(%2't   ��O    ��� Y    @bH@7� c�Y|8��a��K�_�E�w�"��3��T0 k� $�H��H�?�D#B(%2't   ��O    ��� Y    @bH@7� c�Y|8��Q��K�_�E�s�"��3��T0 k� $�I��I�?�D#B(%2't   ��O   ��� Y    @bL@7� c�Y|8��Q��K�_�E�s�"��3��T0 k� �J��J�?�D#B(%2't   ��O    ��� Y    @bL@7� c�Y|8��Q��K�_�E�o�"��3��T0 k� �J��J�?�D#B(%2't   ��O    ��� Y    @bL@7� c�Y|8��Q��K�_�I�k�"��3��T0 k� �K��K�?�D#B(%2't   ��O    ��� Y    @bL@7� c�Y|8��Q��K�_�I�k�"��3��T0 k� �L��L�?�D#B(%2't   ��O    ��� Y    @bL@7� c�Y|8��Q��K�_�I�g�"��3��T0 k� �M��M�?�D#B(%2't   ��O    ��� Y    @bL@7� c�Y|8��Q��K�_�I�g�"��3��T0 k� �N��N�?�D#B(%2't   ��O    ��� Y    @bP@7� c�Y|8��Q��K�_�I�c�"��3��T0 k� �O��O�?�D#B(%2't   ��O    ��� Y    @bP@7� c�Y|8��Q��K�_�I�c�"��3��T0 k� �O��O�?�D#B(%2't   ��O    ��� Y    @bP@7� c�Y|8��Q��K�_�I�c�"��3��T0 k� �P��P�?�D#B(%2't   ��O    ��� Y    @bP@7� c�Y|8��Q��K�_�I�c���3��T0 k� ��Q��Q�?�D#B(%2't   ��O    ��� Y    @bP@7� c�Y|8��Q��K�_�I�_���3��T0 k� �R��R�?�D#B(%2't   ��O    ��� Y    @bP@7� c�Y|8��A��K�_�I�_���3��T0 k� �R��R�?�D#B(%2't   ��O    ��� Y    @bT@7� c�Y|8��A��K�_�I�[���3��T0 k� �S��S�?�D#B(%2't   ��O    ��� Y    @bT@7� c�Y|8��A��K�_�I�[���3��T0 k� �T��T�?�D#B(%2't   ��O    ��� Y    @bT@7� c�Y|8��A��K�_�I�[���3��T0 k� �U��U�?�D#B(%2't   ��O    ��� Y    @bT@7� c�Y|8��A��K�_�I�W����3��T0 k� �U��U�?�D#B(%2't   ��O    ��� Y    @bT@7� c�Y|8��A��K�_�I�W����3��T0 k� �V��V�?�D#B(%2't   ��O    ��� Y    @bT@7� c�Y|8���K�_�I�W����3��T0 k� �W��W�?�D#B(%2't   ��O    ��� Y    @bX@7� c�Y|8���K�_�I�W����3��T0 k� �W��W�?�D#B(%2't   ��O    ��� Y    @bX@7� c�Y|8���K�_�I�S����3��T0 k� �X��X�?�D#B(%2't   ��O    ��� Y    @bX@7� c�Y|8���K�_�I�S����3��T0 k� �Y��Y�?�D#B(%2't   ��O    ��� Y  ��@{��  ��b���S��(@mO�A^C����3�T0 k� �������? t�B(%2't   ��"    ����8  ��@{��  ��b���S��(@mO�A^?����3�T0 k� ����ê�? t�B(%2't   ��"    ����8  ��E��  ��Y����S��(@mO�A^;����3�T0 k� ����ñ�? t�B(%2't   ��"    ����8  ��E��  ��Y����W��)@mO�A^7����"��T0 k� ����ö�? t�B(%2't   ��"    ����8  ��E��  ��Y����W��)@mO�A^3����"��T0 k� ����ú�? t�B(%2't   ��"    ����8  ��E��  ��Y����[��)@mO�A^3����"��T0 k� �þ�Ǿ�? t�B(%2't   ��"   ����8  ��E��  ��Y����[��)@mO�A^/����"��T0 k� �������? t�B(%2't   ��"    ����8  ��E��  ��Y����_��*@mO�A^+����"��T0 k� �����? t�B(%2't   ��"    ����8  ��E��  ��Y����_��*@mO�A^'����"��T0 k� �����É? t�B(%2't   ��"    ����9  ��E��  ��Y����c��*@mO�A^#����"��T0 k� �����ŉ? t�B(%2't   ��"    ����:  ��E��  ��Y����g��*@mO�A^#����"��T0 k� �����Ɖ? t�B(%2't   ��"    ����;  ��E��  ��Y����g��+@mO�A^����"��T0 k� �����Ɖ? t�B(%2't   ��"    ����<  ��E���  ��Y����k��+@mS�A^����"��T0 k� �����ˉ? t�B(%2't   ��"    ����=  ��E���  ��b+���o��+@mS�A^����"��T0 k� �����Ή? t�B(%2't   ��"    ����>  ��E���  ��b+���o��+@mS�A^����3�T0 k� �����щ? t�B(%2't   ��"    ����?  ��E���  ��b+���s��+@mS�A^����3�T0 k� �����ԉ? t�B(%2't   ��"    ����@  ��E���  ��b+���w�|,@mS�A^����3�T0 k� �����Չ? t�B(%2't   ��"    ����A  ��E���  ��b+���w�|,@mS�A^����3�T0 k� ����׉? t�B(%2't   ��"    ����B  ��E���  ��b+���{�|,@mS�A^����3�T0 k� ���؉? t�B(%2't   ��"    ����C  ��E���  ��b+����|,@mS�A^����3�T0 k� ���ډ? t�B(%2't   ��"    ����D  ��E���  ��b+����|,@mS�A^����3�T0 k� ���ډ? t�B(%2't   ��"    ����E  ��E��  ��b+��̃�|-@mS�A]�����3�T0 k� ���ۉ? t�B(%2't   ��"    ����F  ��B\�  ��b+��̃�x-@mS�A]�����3�T0 k� ���#ډ? t�B(%2't   ��"    ����G  ��B\�  ��b+��̇�x-@mS�A]�����3�T0 k� �'��+ى? t�B(%2't   ��"    ����H  ��B\�  ��Y���̇�x-@mS�A]�����3�T0 k� �+��/ى? t�B(%2't   ��"    ����I  ��B\�  ��Y���̋�x-@mS�A]�����3�T0 k� �3��7ډ? t�B(%2't   ��"    ����J  ��B\#�  ��Y���̋�x.@mS�A]�����3�T0 k� �7��;ډ? t�B(%2't   ��"    ����K  ��B\+�  ��Y���̋�x.@mS�A]�����3�T0 k� �?��Cۉ? t�B(%2't   ��"    ����L  ��B\/�  ��Y���̋�t.@mS�A]�����3�T0 k� �G��Kۉ? t�B(%2't   ��"    ����M  ��B\7�  ��Y������x.@mS�A]�����3�T0 k� �K��O܉? t�B(%2't   ��"    ����N  ��B\?�  �߂Y������x.@mS�A]�����3�T0 k� �S��W݉? t�B(%2't   ��"    ����O  ��B\C�  �߂Y������x.@mS�A]�����3�T0 k� �[��_މ? t�B(%2't   ��"    ����P  ��B\K�  �߂Y������x/@mS�A]�����3�T0 k� �c��g߉? t�B(%2't   ��"    ����Q  ��B\S�  �߁Y�����|/@mS�A]�����3�T0 k� �k��o��? t�B(%2't   ��"    ����S  ��Bl[�  �߁Y����{�|/@mW�A]�����3�T0 k� �o��s�? t�B(%2't   ��"    ����U  ��Blc�  �߂Y����w�|/@mW�A]�����3�T0 k� �w��{�? t�B(%2't   ��"    ����W  ��Blg�  �߂Y����s�|/@mW�A]�����3�T0 k� �����? t�B(%2't   ��"    ����Y  ��Blo�  �߂Y����o��/@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����[  ��Blw�  �߂Y����k��0@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����]  ��Bl�  �߃Y����k��0@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����_  ��Bl��  �߃Y����g��0@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����a  ��Bl��  �߃Y����c��0@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����c  ��Bl��  �ۃY����_��0@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����e  ��Bl��  �ۄY����[��0@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����g  ��Bl��  �ۄY����[��0@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����i  ��B|��  �ۄY����W��1@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����k  ��B|��  �ۄY����S��1@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����m  ��B|��  �ۄY����O��1@mW�A]�����3�T0 k� �������? t�B(%2't   ��"    ����o  ��B|��  �ۅY����O��1@mW�A]�����3�T0 k� ������? t�B(%2't   ��"    ����p    @��@��� ���Y�  �����A]�A]�����3� T0 k� �˺�Ϻ�?�D#B(%2't   ��/   0����n    @��@��� ���Y�  �����A]�A]�����3� T0 k� �˺�Ϻ�?�D#B(%2't   /�/   0����o    @��@��� ���Y�  �����A]�A]�����3� T0 k� �Ӵ�״�?�D#B(%2't   ��/ 
  0����p    @l��@��� ���Y�  �����A]�A]�����3� T0 k� �Ӳ�ײ�?�D#B(%2't   ��/ 
  0����q    @l��@��� ���Y��L����A]�A]�����3� T0 k� �װ�۰�?�D#B(%2't   ��O 
  0����r    @l��@�����Y��L����A]�A]�����3� T0 k� �ׯ�ۯ�?�D#B(%2't   ��O 
  0����s    @l��@�����Y��L����A]�A]�����3� T0 k� �ۭ�߭�?�D#B(%2't   ��O 
  0����t    @l��@�����Y��L����A]�A]�����3� T0 k� �۫�߫�?�D#B(%2't   ��O 
  0����t    @��@l����a��L� ��A]�A������"�� T0 k� �ߧ�㧉?�D#B(%2't   ��F 
  0����t    @��@l����a�� �� ��A]�A������"�� T0 k� �ߣ�㣉?�D#B(%2't   ��F 
  0����t    @��@l�����a�� �� ��A]�A������"�� T0 k� �ߠ�㠉?�D#B(%2't   ��F 
  0����t    @��@l�����a�� �� ��A]�A������"�� T0 k� �ߟ�㟉?�D#B(%2't   ��F 
  0����t    @��@l�����a�� �� ��A��A������"�� T0 k� �ߞ�㞉?�D#B(%2't   ��F 
  0����t    B���B������a�� �� l��A��A������"�� T0 k� �ߝ�㝉?�D#B(%2't   ��F 
  0����t    B���B������a�� �� l��A��A������"�� T0 k� �ߜ�㜉?�D#B(%2't   �F 
  0����s    B���B���\��a�� �� l��A��A���]��"�� T0 k� �ߜ�㜉?�D#B(%2't   ��F
  0����r    B���B���\��a�� �� l��A��A���]��"�� T0 k� �ߜ�㜉?�D#B(%2't   ��F 
  0����q    B���B���\��a�� �� l��A��A���]��"�� T0 k� �ߜ�㜉?�D#B(%2't   ��F 
  0����p    B���O��\��a�� ��]�A��A���]��"�� T0 k� �ߜ�㜉?�D#B(%2't   ��F 
  0����o    B���O��\��Y�� ��]�A��A���]��3� T0 k� �ߜ�㜉?�D#B(%2't   ��F 
  0����n    B���O����Y�� ��]�A��BM��M��3� T0 k� �ߜ�㜉?�D#B(%2't   ��F 
  0����m    B���O����Y�� ��]�A��BM��M��3� T0 k� �ߜ�㜉?�D#B(%2't   ��F 
  0����l    B���O����Y�� ��]�D��BM��M��3� T0 k� �ߜ�㜉?�D#B(%2't   ��F 
  0����k    B���O����Y�� ��m�D��BM��M��3� T0 k� �ߝ�㝉?�D#B(%2't   ��F   0����j    B���O����Y�� ��m�D��BM��M��3� T0 k� �ߝ�㝉?�D#B(%2't   ��F   0����i    E��O�� ���Y�� ��m�D��@��M��3� T0 k� �ߝ�㝉?�D#B(%2't   ��F   0����h    E��O�� ���Y�� ��m�D��@��M��3� T0 k� �ߝ�㝉?�D#B(%2't   ��F   0����g    EúO�� ���Y�� ��m�D��@��=��3� T0 k� �ߝ�㝉?�D#B(%2't   ��F   0����f    EúO�� ���Y�� ��m�D}�@��=��3� T0 k� �ߞ�㞉?�D#B(%2't   ��F   0����e    EúO�� ���Y�� ��}#�D}�@��=��3� T0 k� �ߞ�㞉?�D#B(%2't   ��F   0����c    eǺO�����Y�� ��}#�D}�B���=��3� T0 k� �ߞ�㞉?�D#B(%2't   ��F   0����a    e˻O�����Y�� ��}'�D}�B���=��3� T0 k� �ߞ�㞉?�D#B(%2't   ��F   0����_    e˻O�����Y�� ��}+�D}�B���=��3� T0 k� �ߞ�㞉?�D#B(%2't   ��F   0����]    eϻO�����Y�� ��}+�D}�B���=��3� T0 k� �ߟ�㟉?�D#B(%2't   ��F   0����[    eϻO�����Y�� ��}/�D}�B���-��3� T0 k� �ߟ�㟉?�D#B(%2't   ��F   0����Y    eӻO�����Y�� ��}/�D}�B���-��3� T0 k� �ߟ�㟉?�D#B(%2't   ��F   0����W    eӼO�����Y�� ��}3�D}�B���-��3� T0 k� �ߟ�㟉?�D#B(%2't   ��F   0����U    e׼O�����Y�� ��}3�D}�B���-��3� T0 k� �ߟ�㟉?�D#B(%2't   ��F   0����S    eۼO�����Y�� ��}7�D}#�B���-��3� T0 k� �ߠ�㠉?�D#B(%2't   ��F   0����Q    eۼO�����Y�� ��};�D}'�B������3� T0 k� �ߠ�㠉?�D#B(%2't   ��F   0����O    e,߼O�����Y�� ��};�D}'�B������3� T0 k� �ߠ�㠉?�D#B(%2't   ��F   0����M    e,߽E�����Y�� ��}?�D}+�B������3� T0 k� �ߠ�㠉?�D#B(%2't   ��F   0����K    e,�E����Y�� ��}?�D}+�B������3� T0 k� �ߠ�㠉?�D#B(%2't   ��F   0����I    e,�E����Y�� ��}C�D}/�B������3� T0 k� �ߠ�㠉?�D#B(%2't   ��F   0����G    e,�E����Y�� ��}C�D}/�B������3� T0 k� �ߡ�㡉?�D#B(%2't   ��F   0����F    e,�E����Y�� ��}G�D}3�B������3� T0 k� �ߡ�㡉?�D#B(%2't   ��F   0����E    e,�E�����Y����}G�D}3�B�é���3� T0 k� �ߡ�㡉?�D#B(%2't   ��O   0����D    e,�E��<��Y����}K�D}7�B�ǩ��3� T0 k� �۠�ߠ�?�D#B(%2't   ��D   0����C    e,�E��<��Y�����}K�D}7�B�˩��3� T0 k� �נ�۠�?�D#B(%2't   ��D   0����B    e,�E��<��Y�����}O�D}7�B�ө� 3� T0 k� �ן�۟�?�D#B(%2't   ��D   0����A    e�E��<��Y�����}O�D};�B�ש�3� T0 k� �ӟ�ן�?�D#B(%2't   ��D   0����@    e�E��<��Y�����}S�D};�B�۩�3� T0 k� �Ϡ�Ӡ�?�D#B(%2't   ��D   0����?    e�E��<��Y�����}S�D}?�B�ߩ-�3� T0 k� �Ϡ�Ӡ�?�D#B(%2't   ��D   0����>    e��E}�L��Y�����}W�D}?�B��-�3� T0 k� �ע�ۢ�?�D#B(%2't   ��D   0����=    e��E}�L��Y�����}[�D}C�B��-�3� T0 k� �ۢ�ߢ�?�D#B(%2't   ��D   0����=    e��E}�L��Y�����}[�D}C�B��-�3� T0 k� �ߢ�㢉?�D#B(%2't   ��D   0����=    e��E}�L��Y�����}_�D}C�B���-�3� T0 k� ���磉?�D#B(%2't   ��D   0����=    e��E}�L��Y�����}_�D}G�B����3� T0 k� ���磉?�D#B(%2't   ��D   0����=    e��E}�L��Y�����}c�D}G�B���	3� T0 k� ���뤉?�D#B(%2't   ��D   0����=    e��E}�L��Y�����}c�D}K�B���
3� T0 k� ���뤉?�D#B(%2't   ��D   0����=    e-�E}�L��Y����}g�D}K�B���3� T0 k� ���뤉?�D#B(%2't   ��D   0����=    e-�D�#�L��Y����}k�D}K�B���3� T0 k� ���륉?�D#B(%2't   ��D   0����=    e-�D�#�<��Y����}k�D}O�B����3� T0 k� ���礉?�D#B(%2't   ��D   0����=    e-�D�'�<��Y����}o�D}O�B�#���3� T0 k� ���礉?�D#B(%2't   ��D   0����=    e-�D�'�<��Y����}o�D}S�B�'���3� T0 k� �ߥ�㥉?�D#B(%2't   ��D   0����>    e-�D�+�<��Y����}s�D}S�B�/���3� T0 k� �ۥ�ߥ�?�D#B(%2't   ��D   0����?    e-�D�+�<��Y����}s�D}S�B�7���3� T0 k� �ۥ�ߥ�?�D#B(%2't   ��D   0����@    e-�D�/� |ÓY����}w�D}W�B�?���3� T0 k� �ߧ�㧉?�D#B(%2't   ��D   0����A    e-�D�/� |ÓY����}w�D}W�B�C���3� T0 k� ���秉?�D#B(%2't   ��D   0����B    e-�D�3� |ÓY����}{�D}W�B�K���3� T0 k� ���稉?�D#B(%2't   ��D   0����C    e-�D�3� |ǔY����}{�F[�B�S���3� T0 k� ���稉?�D#B(%2't   ��D   0����D    E�D�3� |ǔY����}�F[�B�[���3� T0 k� ���먉?�D#B(%2't   ��D   0����E    E�D�7� |ǕY����}�F_�B�c���3� T0 k� ���멉?�D#B(%2't   ��D   0����F    E�D�7� |˕Y����}�F_�B�k���3� T0 k� ���몉?�D#B(%2't   ��D   0����G    E�D�7� |˖Y����}��Fc�B�s���3� T0 k� ���憎?�D#B(%2't   ��D   0����H    E�D�7� |˖Y����}��Fc�B�{���3� T0 k� ���韛?�D#B(%2't   ��D   0����I    E��D�7� |˖Y����}��E�g�B�����3� T0 k� ����?�D#B(%2't   ��D   0����J    E��D�7� |˗Y����}��E�k�B�����3� T0 k� ����?�D#B(%2't   ��D   0����K    E�#�D�7� |ϗY����}��E�k�B�����3� T0 k� ����?�D#B(%2't   ��D   0����L    E�#�D�7� �ϘY����}��E�o�B�����3� T0 k� ����?�D#B(%2't   ��D  0����M    E�'�D�7� �ϙY����}��E�s�B�����3� T0 k� ����?�D#B(%2't   ��D   0����N    D�'�D�7� �ϙY����}��B�w�B�����3� T0 k� ����?�D#B(%2't   ��D   0����O    D�+�D�7� �ϚY����}��B�{�B�����3� T0 k� ����?�D#B(%2't   ��D  0����P    D�/�A�7� �ӛY����}��B��B�����3� T0 k� ����?�D#B(%2't   ��D   0����Q    D�/�A�7� �ӛY����}��B���B�ǩ��3� T0 k� ������?�D#B(%2't   ��D   0����R    D�3�A�7� �לY����}��B���B�ө�3� T0 k� ������?�D#B(%2't   ��D   0����S    F7�A�7� �םY����}��B���B�۩�3� T0 k� �������?�D#B(%2't   ��D   0����T    F7�A�7� �۞Y����}��B���B��� 3� T0 k� �������?�D#B(%2't   ��D   0����U    F;�A�7� �۟Y����}��B���B��� 3� T0 k� �������?�D#B(%2't   ��D   0����V    F?�A�7� �ߟY���#�}��B���B���!3� T0 k� ������?�D#B(%2't   ��D   0����W    FC�A�7� �ߠY���#�}��B���B���� "3� T0 k� ������?�D#B(%2't   ��D   0����X    FG�A�7� ��Y���#�}��B���B���$"3� T0 k� �����?�D#B(%2't   ��D   0����Y    FK�A�7� ��Y���'�}��B���B���,#3� T0 k� �����?�D#B(%2't   ��D  0����Z    D�O�A�7� ��Y���'�}��B���B���4#3� T0 k� �����?�D#B(%2't   ��D   0����[    D�S�A�7� ��Y���'�}��B���B�#��8$3� T0 k� �����?�D#B(%2't   ��D   0����\    D�W�A�7�,�Y���+�}��B���B�+��@$3� T0 k� �����?�D#B(%2't   ��D  0����]    D�[�A�7�,�Y���+�}��B���B�3��H%3� T0 k� �����?�D#B(%2't   ��D   0����^    D�_�A�7�,�Y���+�}��B���B�;��L%3� T0 k� �����?�D#B(%2't   ��D   0����_    D�c�A�7�,��Y���+�}��B���B�C��T&3� T0 k� �����?�D#B(%2't   ��D   0����`    D�g�A�7�,��Y���/�}��B���B�O��\'3� T0 k� �����?�D#B(%2't   ��D   0����b    D�k�A�7���Y���/�}��B���B�W��d'3� T0 k� �����?�D#B(%2't   ��D   0����d    D�s�A�7��Y���/�}��B���B�_��h(3� T0 k� �����?�D#B(%2't   ��D   0����f    D�w�A�7��Y���3�}��B���B�g��p(3� T0 k� �����?�D#B(%2't   ��D   0����h    D�{�A]7��Y���3�}��B���B�s��x)3� T0 k� ���#��?�D#B(%2't   ��D   0����j    D��A]7��Y���3�}��B���B�{���)3� T0 k� �#��'��?�D#B(%2't   ��D   0����l    D��A]7��Y���3�}��B��B߃���)3� T0 k� �'��+��?�D#B(%2't   ��D   0����n    D��A]7��Y���7�}��B��Bߋ���*3� T0 k� �+��/��?�D#B(%2't   ��D   0����p    D��A]7��Y���7�}��B��Bߓ���*3� T0 k� �/��3��?�D#B(%2't   ��D   0����r    D��A]7��Y���7�}��B��Bߟ���+3� T0 k� �3��7��?�D#B(%2't   ��D   0����t    D��A]7�#�Y���7�}��B�'�Bߧ���+3� T0 k� �7��;��?�D#B(%2't   ��D   0����v    D��A]7��'�Y���;�}��B�/�B߯���,3� T0 k� �;��?��?�D#B(%2't   ��D   0����w    D��A]7��/�Y���;�}��B�7�B߷���,3� T0 k� �C��G��?�D#B(%2't   ��D   0����y    D��A]7��3�Y���;�}��B�C�B߿���-3� T0 k� �G��K��?�D#B(%2't   ��D   0����{    D��A]7��7�Y���;�}��B�K�B�˩��-3� T0 k� �K��O��?�D#B(%2't   ��D   0����}    D��A]7��;�Y���?�}��B�S�B�ө��-3� T0 k� �O��S��?�D#B(%2't   ��D   0����~    D��A7�]?�Y���?�}��B�_�B�۩��.3� T0 k� �W��[��?�D#B(%2't   ��D   0�����    D���A7�]G�Y���?�}��B�g�B����.3� T0 k� �[��_��?�D#B(%2't   ��D   0�����    D���A7�]K�Y���?�}��B�o�B����/3� T0 k� �_��c��?�D#B(%2't   ��D   0�����    D���A7�]O�Y���C�}��B�{�B�����/3� T0 k� �g��k��?�D#B(%2't   ��D   0�����    D���A7�]W�Y���C�}��I��B�����/3� T0 k� �k��o��?�D#B(%2't   ��D   0�����    D���A7�][�Y���C�}��I��B���03� T0 k� �o��s��?�D#B(%2't   ��D   0�����    D���A7�]_�Y���C�}��I��J@��03� T0 k� �w��{��?�D#B(%2't   ��D   0�����    D���A7�]g�Y���C�}��I��J@��13� T0 k� �{����?�D#B(%2't   ��D   0�����    D���A7�mk�Y���G�}��I��J@�� 13� T0 k� ������?�D#B(%2't   ��D   0�����    D���A7�mo�Y���G�}��I.��J@'��(13� T0 k� �������?�D#B(%2't   ��D   0�����    D���A7�mw�Y���G�}��I.��J@/��023� T0 k� �������?�D#B(%2't   ��D   0�����    D���A7�m{�Y���G�}��I.��E 7��823� T0 k� �������?�D#B(%2't   ��D   0�����    E��@�7�m��Y���K�}��I.��E ?��@23� T0 k� �������?�D#B(%2't   ��D   0�����    E��@�7�m��Y���K�}��I.��E C��L33� T0 k� �������?�D#B(%2't   ��D   0�����    E��@�7�m��Y���K�}��I��E K��T33� T0 k� �������?�D#B(%2't   ��D   0�����    E��@�7�m��Y���K����I��E O��\33� T0 k� �������?�D#B(%2't   ��D   0�����    E��@�7�m��Y���K����I��E W��d43� T0 k� �������?�D#B(%2't   ��D  0�����    E��@�7�m��Y���K��� I��E0[��l43� T0 k� �������?�D#B(%2't   ��D   0�����    E��@�7�m��Y���O���I��E0c��x43� T0 k� �������?�D#B(%2't   ��D   0�����    E��@�7�}��Y���O�� I.��E0g�π43� T0 k� �ë�ǫ�?�D#B(%2't   ��D   0�����    E��@�7�}��Y���O��I.��E0o�ψ53� T0 k� �ǫ�˫�?�D#B(%2't   ��D   0�����    E��@�7�}��Y���O��I.��E0s�ϐ53� T0 k� �ϫ�ӫ�?�D#B(%2't   ��D   0�����    E��@�7�}��Y���O��I.��E0w�Ϙ53� T0 k� �ӫ�׫�?�D#B(%2't   ��D   0�����    D���@�7�}ûY���O��I.��E0{�ߤ63� T0 k� �۪�ߪ�?�D#B(%2't   ��D   0�����    D���@m7��˺Y���S�.I��E0��߬63� T0 k� �߮�㮉?�D#B(%2't   ��D   0�����    D��@m7��ϺY���S�.I��E0��ߴ63� T0 k� ���뱉?�D#B(%2't   ��D   0�����    D��@m7��׺Y�#��S�.I�E0��߼63� T0 k� ����?�D#B(%2't   ��D   0�����    D��@m7��ߺY�#��S�.	I�E@����73� T0 k� ������?�D#B(%2't   ��D   0�����    D��@m7���Y�#��S�.
I�E@����73� T0 k� �������?�D#B(%2't   ��D   0�����    D��@m7���Y�#��S�.I/�E@����73� T0 k� �����?�D#B(%2't   ��D   0�����    D��@m7���Y�#��W�.I/�E@����83� T0 k� �����?�D#B(%2't   ��D   0�����    D��@m7����Y�#��W�. I/�E@����83� T0 k� �����?�D#B(%2't   ��D   0�����    D��@m7����Y�#��W�.$I/�E@����83� T0 k� �����?�D#B(%2't   ��D   0�����    D��@m7���Y�#��W�.$I/�E@����83� T0 k� ���#��?�D#B(%2't   ��D   0�����    D�'�@m7���Y�#��W��(I�E@���93� T0 k� �'��+��?�D#B(%2't   ��D   0�����    D�+�@m7���Y�#��W��(I�E@���93� T0 k� �/��3��?�D#B(%2't   ��D   0�����    D�3�@m7���Y�#��W��,I�E@ü�93� T0 k� �7��;��?�D#B(%2't   ��D   0�����    D�8 @m7��'�Y�#��[��0I�E@Ǿ�93� T0 k� �?��C��?�D#B(%2't   ��D   0�����    D�<@m7��/�Y|'��[��4I�E�Ͽ�$93� T0 k� �G��K��?�D#B(%2't   ��D   0�����    D�D@m7��3�Y|'��[��4I/�E���0093� T0 k� �K��O?�D#B(%2't   ��D   0�����    D�H@m7�;�Y|'��[��8I/�E���0893� T0 k� �O��S��?�D#B(%2't   ��D   0�����    D�P@m7�C�Y|'��[��<I/#�E���0@93� T0 k� �W��[��?�D#B(%2't   ��D   0�����    D�X@m7�K�Y|'��[��<I/#�E���0D93� T0 k� �_��c��?�D#B(%2't   ��D   0�����    D�`@m7�S�Y|+��[��@I/'�E���0L93� T0 k� �g��k��?�D#B(%2't   ��D   0�����    D�d@m7�[�Y|+��[�NDB�+�E���0T83� T0 k� �o��s��?�D#B(%2't   ��D   0�����    D�l
@m7�c�Y|+��_�NDB�+�E���0\83� T0 k� �w��{��?�D#B(%2't   ��D   0�����    D�t@m7�k�Y|+��_�NHB�/�E���0d83� T0 k� ������?�D#B(%2't   ��D   0�����    D�|@m7��s�Y|+��_�NLB�3�E���@l73� T0 k� �������?�D#B(%2't   ��D   0�����    D��@m7��{�Y|+��_�NL B�7�E���@t73� T0 k� �������?�D#B(%2't   ��D   0�����    D��@m7����Y|+��_�NP"B�;�E���@|73� T0 k� �������?�D#B(%2't   ��D   0�����    D��@m7����Y|+��_�NT#B�?�E���@�63� T0 k� �������?�D#B(%2't   ��D   0�����    D��@m7����Y|+��_�NT%B�C�E���@�63� T0 k� �������?�D#B(%2't   ��D   0�����    I��@m7����Y|+��_�NX&B�G�E���@�53� T0 k� �������?�D#B(%2't   ��D   0�����    I��@m7����Y|+��_�NX(B�K�E��@�53� T0 k� �������?�D#B(%2't   ��D   0�����    I��@m7����Y|+��c�N\*B�O�E��@�43� T0 k� ����ß�?�D#B(%2't   ��D   0�����    I��@m7����Y|+��c�N`+B�S�E��@�33� T0 k� �Ǟ�˞�?�D#B(%2't   ��D   0�����    I��@m7�^��Y|+�=c�^`-B�W�E��@�33� T0 k� �ϟ�ӟ�?�D#B(%2't   ��D   0�����    I��@m7�^ǴY|+�=c�^d/B�_�E��@�23� T0 k� �נ�۠�?�D#B(%2't   ��D   0�����                                                                                                                                                                            � � �  �  �  c A�  �J����  �      � \��Y� ]�3�3� � �#�C�         �  �V    �C�  �V               ��  	 ����         T�       ���   8�         ���         �  ��    ���  ��               ��        
	 ���         �       ���   H
          ��         �VG     �  �2'    ��               4         n     ���   (	          ����         �M��    �����M��                        	  �$           �     ���   H
4
           ^.         . �rJ     #% �{    y�   	             ��$          3�  �  ���   P
	B          Nv ��     B��     L#��     #                      ���i               ?  ���    8		 1             ��Ƥ  �<	     V�_W�    ��Ƥ�_W�                    �� Y         	�    ��h   8
(
         ��j@  � �	   j bi�    ���g c�    �I��             �� Y�        � �   	  ��`  @

"          ��S� � �
    ~ W��    ��EQ W��     @             	�� Y�         0       ��@    

'          ��?� � �	    � Tݲ    ��?� T��      �            	�� Y         	 �@�     ��@  8
          ��7�  > > 
	  � �x�    ��O� ��    ���m            # )�� Y         
 ���     ��@   X
         ��sM ��
      � �_�    ��t� �_�    ��                         ���R              ?  ��@    0 0 	                 ��      �                                                                           �                               ��        ���          ��                                                                 �                          YE  ��        �!7�     X�!x�    
��-                x                j  �   �   �                          Y    ��        �"       X  "           "                                                �                              ��M ���_ b W T � ���!"   	        
      
    F�n [�C       �d �r@ �� s@ ��  s` �� s� �� �m@ �� n@ �� 0n` �D  n� �� o  #� `t� $d u� �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ���� � 
�\ U� 
�| V  
�| V ���� � � 0i@ �d  i� פ i� �$ �j� �$ k� �D k� �d l  Є l  Ф l@ �� 0m@ �D  m� ̄ 0m� �� n@ � 0n` �� �o� �� p� �� t� � �t� �  u����� � $d p� ?� �[� @� 0\� A ]  A$ ]@ 
�| U� 
� V  
�\ V  
�< V� 
�� V� 
�| W  
�| W� 
� W� 
�\ W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� Y ������  ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"     "�j��   * �
� �  �  
� ��    ��     �   �        ��     � �      ��    ��     ��_          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �OBB(      ��R �  ��        � �T ��        �        ��        �        ��        �    ��     � f�        ��                         ��  0  �����                                     �                 ����            �� ���%��  �� Y 2���2           �CHI my Roenick      0:00                                                                        6  6     � �
"�EC
� � �k� � � � � �k� � � k� � �	k~ � �k� � �	k� � �
cj � � cr � �cs � �cv � � cx � �KC �K3 �c� � c� �  "H � � ". | � "@ | � "P � � "& |	 "* |Y  "P � �"2 | � "@ | � "P � � "& |	 "* |Y  "P �Y  "J �Y  "P �	 ""* |Y  "P � � $"& |	 %"* |Y  "P � � '"& |	 ("* |Y  "P � � *"J � +"  |8,!� |`  "O �Z  "O �6/"2 |V 0"@ |V ": �T 2"@ |T ": �S "  |_  " �C6"* |[ "< �`  "D � �9!� �:"  |(;!� |P <"I �`  "P �X  *K=X  *K=                                                                                                                                                                                                                         L� P `            @ 
        �     e P E i  ������               �������������������������������������� ���������	�
��������                                                                                          ��    ���    ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, ;  B }�  ���� �� �� ���@���@A��W���������                                                                                                                                                                                                                                                                                                        2�����"                                                                                                                                                                                                                                          $ #    ��  L�J      #�                             ������������������������������������������������������*�                                                                                                                                     �    ��              7          ��   � 
           	 	 ���� ������������� ������ �����������   ������������� ������������������ ���� ��������������������� ��� ���  �������������� ����� �������������� �������  ���������� ������������������������������ ������������������ ������������ �                              X  	  (    ��  4�J      :  	                           ������������������������������������������������������                                                                                                                                          �  ��              �          ��               	 
     � ����� �����  � ��������������� ������ ����������� � ����������� ���� ����� ���  ����� ���  ������ � ������� ��������������������� �� ���������������� ��� ��������������������������� � ��������������������������� ���������           �                                                                                                                                                                                                                                                                                                  	         �             


           �   }�         ������������  z   ����������������������������    ������������������������  N�������������������������                                     vg                 'u  'u                     �ww�ww333wwwwwwww�ww�ww�ww�ww333wwww % K ?                                 � [ �\                                                                                                                                                                                                                                                                                     	�)nY  
)n        `      e                  k            m                                                                                                                                                                                                                                                                                                                                                                                                              0 '  � ��  � ��  � @��  � #��  � ��  ��(�������������������{�����������������8�����2          .         K          �   & AG� �   �   
           ���                                                                                                                                                                                                                                                                                                                                    p I N   �      ��               !��                                                                                                                                                                                                                            Y   �� �� Ѱ�      �� Z      ���� ������������� ������ �����������   ������������� ������������������ ���� ��������������������� ��� ���  �������������� ����� �������������� �������  ���������� ������������������������������ ������������������ ������������ �� ����� �����  � ��������������� ������ ����������� � ����������� ���� ����� ���  ����� ���  ������ � ������� ��������������������� �� ���������������� ��� ��������������������������� � ��������������������������� ���������      �     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    3      3    �  X                       4     �  �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$ ^h  ��     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@       �      �     ��    `d � � ��� �� � ��� �$ L �  ��L  �      �  ��   /���� e����J  g���        f ^�         �� q��      /      ��ZX�������J���J��~����      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 " ""   "" "!  "" "  """ !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                   " ""   "" "!  "" "  """ !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """ "! ""! " ""  !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r`��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �    �   "   "   "  �  �   �         +  "  "     �  �                        �   ���                            �   �                                                                                                   ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r`                         ����    
�  ��  ��  ��  �����  �   �          ��                           � ��                    ���� �                                                                                                                                                                                                              	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                       ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                            �������  ���    �    �   �   �   D   E�  U�  UO                         "  "  "                    �   ���                            �   �                                                                                                                         	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                       "   "  !�    ��                              �                        ���� ��� ����                            ��  ��  ���              �  �˰ ��� �wp ���                                                                                                                                                                                       	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                         �  �  �  �  �   �       �               �    �                    �   �   �                                   ��  ��  ���              �  �˰ ��� �wp ���                                                                                                                                                                                 �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �   ��  �  ��  ��  ��� �� /   �           �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                                           "" "" ""�/"  "  "  " "" �"/ �/� I� U� DU� 3EY CEZ 4T�"4U��4U���U�/DZ�"�J�+ʌ�+������ �   �   ��ɪ��ɪ��̚���ț��̋ ��P ��P���_��������������  �            �   �   ��  �"  "  �"  �/  ��  �   �   �" �""� �"���             � �� �  � �� �                         �  �  �� ���  � �� �   �   �      �                                � �� ���H���     ̰ �˻���ݹ��w���&ɧvvɪ�p              �  �� �� �� ��                         ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                     w 
�� ɚ� ���
�˻Ɋ�����������-� �"+ ". "$ "$ �U  Z�  Z�  J�  J�  �D  ��  ��  ɘ ˰ "  �"/�"" "  �  �            g���z��ȩ�����ة�� ���  ̰  ̰  ˰  ��  �  N�� T4�CD  CD0 C40 C30 3;� ܰ �� �� �  �  "  �""�"" �"/���  � �  �      �     �   �   ��  �"" �""  ""   "                 �   ��   �                            � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                                       "  "(��ȩ�ܚ��ۊ����� ��  �   �   �   �   �� ��� ̻� ˽� ��� �w� �������������������������� �̻ ���         �   �       �   �   "" �+� Ȼ� ɫ� ɨ� ��                �� �I��3 ��D 
UD 
UD TD  T�  ˸  ��  �� ̰ �+ ��"/ �"/  ����  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �   �   �                .                      ��  ��  ���  ��  �  �  �   �                                                                                                                                                                                           �   �   �   b   g   �  
�  �� �� �� �̻ ������ɨ�-�ݼ-ݍ�"Չ� X���DDX�TCZES3�T3�@ ��"��"�� ""� �"/��/��        �   ��  ��  ��  ��  wp  ��� ���������̻��̽��̽���ؚ��ڨ��؛˻��˸� ��  �C  D0  3   0   0   �   �   �    �  /   ���             0  #! 02�>0 1                     �    � �� �  �� 	  
  �  ",  ""  �"   "                      ��  ��  �               �������  ���    �                    ��� ���� ��  ���� �                                                                                                                                                                                         � 
��	�˽���w��{k��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            �  �  �  ��  �           / �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw  ��  �   ��  �                                        ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                                     �� ̻ ��˛��  �� �˚̻���ۚ����I���䘼�^���^�٘�:�^�� ^�� D�( �) �) �) ��) ˹� ț�+��,��,����  �𫝝 ��� �ɍ ��ݨ��ډ�݊�� ��D@ �D�  J�� ݩ� ��� �ۻ �ک �ڹ�ɻ��̸���������� ����������            �   ��  ��  ��  ��  ��                                          �� ��� ��� ��  �                         �   �   �" �!  �  �� �   �                �  �� Ș ��  ��  �    ��˰ɜ˰��˻�̻���������3���DDD�                                                                                                                                                                                                             �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
"�DC
� � �k� � � � � �k� � � k� � �	k~ � �k� � �	k� � �
cj � � cr � �cs � �cv � � cx � �KC �K3 �c� � c� �  "H � � ". | � "@ | � "P � � "& |	 "* |Y  "P � �"2 | � "@ | � "P � � "& |	 "* |Y  "P �Y  "J �Y  "P �	 ""* |Y  "P � � $"& |	 %"* |Y  "P � � '"& |	 ("* |Y  "P � � *"J � +"  |8,!� |`  "O �Z  "O �6/"2 |V 0"@ |V ": �T 2"@ |T ": �S "  |_  " �C6"* |[ "< �`  "D � �9!� �:"  |(;!� |P <"I �`  "P �X  *K=X  *K=3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0�������������������������������������������-�N�X�O�Y�Z�G�T��;�[�[�Z�Z�[� � � � � �-�2�3�����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������-�2�3� ��!�������������������������������������-�2�3�	�
�������������������� � � � � � �����������������������������������������%��������������������,�>�0� �� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                