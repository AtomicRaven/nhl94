GST@�                                                            \     �                                               � ��     �  >            ����e $�	 J�����������x�������        �g     	#    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"      �j* , . ���
��
�"   "D�j��
� " ��
  �                                                                               ����������������������������������       ��    =b 0Qb 4 114  4c  c  c        	 
      	   
       ��G �� � ( �(                 nn 
)1         88�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             �n  11          == �����������������������������������������������������������������������������                                �|  |      ��   @  #   �   �                                                                                '      
)n1n  1�1n    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E x �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    	�S7�M\�>[�nB�<L��B�i@��@lh[_�S��`Z3�T0 k� ��L��L2d qD�QC"3Q  ��"    � 3�;	�S3�M\�?[�nB�@L��B��h@��@ll[_�S��`Z3�T0 k� ��L��L2d qD�QC"3Q  ��"    � 3�;	�S3�M\�?[�nB�DL��B��h@��@ll[_�S��_Z3�T0 k� ��L��L2d qD�QC"3Q  ��"    � 3�;	�S3�M\�@[�nB�HL��B��g@��@lp[_�S��_Z3�T0 k� ��M��M2d qD�QC"3Q  ��"    � 3�;	�S/�M\�@�nB�LM��B��g@��@lp[_�S��^Z3�T0 k� ��M��M2d qD�QC"3Q  ��"    � 3�;	� S/�M\�@�nB�PM��B��f@��@lt[_�S��]Z3�T0 k� ��M��M2d qD�QC"3Q  ��"    � 3�;	� S+�M\�A�nB�TM��B��f@��@lx[_�S��]Z3�T0 k� ��N��N2d qD�QC"3Q  ��"    � 3�;	��S+�M\�A�nB�TM��B��e@��@lx\_�S��\Z3�T0 k� ��N��N2d qD�QC"3Q  ��"    � 3�;	��S'�E|�B�nB�XM��B��e@���@l|\_�S��\Z3�T0 k� ��Q��Q2d qD�QC"3Q  ��"    � 3�;	��S'�E|�B�nB�\M��B� d@���@l|\_�S��[Z3�T0 k� ��S��S2d qD�QC"3Q  ��"    � 3�;	��S'�E|�B�nB�`M��B�d@���@l�\_�S��[Z3�T0 k� ��T��T2d qD�QC"3Q  ��"    � 3�;	��S#�E|�C�nB�dM��B�c@���@l�\_�S��ZZ3�T0 k� ��V��V2d qD�QC"3Q  ��"    � 3�;	��S#�E|�C�nB�hM��B�c@���@l�\_�S��ZZ3�T0 k� ��W��W2d qD�QC"3Q  ��"    � 3�;	��S�E|�C�nB�hM��B�b@���@l�]_�S�|YZ3�T0 k� ��X��X2d qD�QC"3Q  ��"    � 3�;	��S�A��D�nB�lM��B� b@���@l�]_�S�|YZ3�T0 k� ��W��W2d qD�QC"3Q  ��"    � 3�;	��S�A��D�nB�lM��B�(b@���@l�]_�S�|XZ3�T0 k� ��U��U2d qD�QC"3Q  ��"    � 3�;�S�A��D�nB�lM��B�,a@���@l�]_�S�|WZ3�T0 k� ��T��T2d qD�QC"3Q  ��"    � 3�;�S�A��D�nE�pN��B�4a@���@l�^_�S�|WZ3�T0 k� ��S��S2d qD�QC"3Q  ��"    � 3�;�S�A��D+�nE�tN��B�<`@���@l�^_�S�|VZ3�T0 k� ��R��R2d qD�QC"3Q  ��"    � 3�;�S�F�D+�nE�tO��B�@`@���@l�^_�S�|VZ3�T0 k� ��R��R2d qD�QC"3Q  ��"    � 3�;�S�F�D+�nE�xO��B�H`@���@l�^_�S�|UZ3�T0 k� ��R��R2d qD�QC"3Q  ��"    � 3�;�S�F�D+�nE�xO��B�L_@���@l�__�S�|TZ3�T0 k� ��R��R2d qD�QC"3Q  ��"    � 3�;�S�F�D+�nE�|O��B�T_@���@l�__�S�|TZ3�T0 k� ��R��R2d qD�QC"3Q  ��"    � 3�;�S�F�E+�nE��O��B�X^@���@l�__�S�|SZ3�T0 k� ��S��S2d qD�QC"3Q  ��"    � 3�;�S�E��E+�nD܄P��B�\^@���@l�`_|S�|SZ3�T0 k� ��O��O2d qD�QC"3Q  ��"    � 3�;�S�E��E+�nD܈P��@md^@���@l�`_|S�|RZ3�T0 k� ��L��L2d qD�QC"3Q  ��"    � 3�;�S�E��E+�nD܈Q��@mh]@���@l�a_xS�|RZ3�T0 k� ��J��J2d qD�QC"3Q  ��"    � 3�;�S�E��E+�nD܌Q��@ml]@���@l�a_tS�|QZ3�T0 k� ��H��H2d qD�QC"3Q  ��"    � 3�;�S�E��E+�nDܐQ��@mt]@���@l�a_pS�|QZ3�T0 k� ��G��G2d qD�QC"3Q  ��"    � 3�;�T�E��E+�nDܔR��@mx\@���@l�b_lS�|PZ3�T0 k� ��B��B2d qD�QC"3Q  ��"    � 3�;,�T�E��D+�nDܔR��@m|\@���@l�b_hS�|PZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�;,�T��E��D+�nDܘR��@m�\@���@l�c_hS�|OZ3�T0 k� ��;��;2d qD�QC"3Q  ��"   � 3�;,�T��E��D+�nDܘR��@m�[@���@l�c_dS�|OZ3�T0 k� ��9��92d qD�QC"3Q  ��"    � 3�;,�T��E��C+�nDܜR��@m�[@���@l�c_`S�|NZ3�T0 k� ��7��72d qD�QC"3Q  ��"    � 3�;,�U��E��C+�nDܜS��@m�[@���@l�d_\S�|NZ3�T0 k� ��4��42d qD�QC"3Q  ��"    � 3�;,�U��E��C+�nDܠS��@m�Z@���@l�d_\S�|MZ3�T0 k� ��2��22d qD�QC"3Q  ��"    � 3�;,�U��E��B+�nD�S��@m�Z@���@l�d_XS�|MZ3�T0 k� ��/��/2d qD�QC"3Q  ��"    � 3�;,�U�E��B+�nD�S�� @m�Z@���@l�e_TS�|LZ3�T0 k� ��.��.2d qD�QC"3Q  ��"    � 3�;,�U�E��A+�nD�S�� @m�Z@���@l�e_PS�|LZ3�T0 k� ��,��,2d qD�QC"3Q  ��"   � 3�;,�V��E��@+�nD�S�� @m�Y@���@l�e_PS�|KZ3�T0 k� ��*��*2d qD�QC"3Q  ��"    � 3�;,�V��E��@+�nD�S�� @m�Y@���@l�f_LS�|KZ3�T0 k� ��*��*2d qD�QC"3Q  ��"    � 3�;,�V��E��?+�nB��S�� @m�Y@���@l�f_HS�|KZ3�T0 k� ��)��)2d qD�QC"3Q  ��"    � 3�;,�V<��E��>+�nB��S��!@m�X@���@l�f_HS�|JZ3�T0 k� ��(��(2d qD�QC"3Q  ��"    � 3�;,�V<��E��=+�nB��R��!@m�X@���@l�g_DS�|JZ3�T0 k� ��'��'2d qD�QC"3Q  ��"    � 3�;,�W<��E��=+�nB��R��!@m�X@���@l�g_@S�|IZ3�T0 k� ��&��&2d qD�QC"3Q  ��"   � 3�;,�W<��E��<+�nB��R��!@m�X@���@l�g_@S�|IZ3�T0 k� ��(��(2d qD�QC"3Q  ��"    � 3�;,�W<��E��;+�nB��R��!@m�W@���@l�g_<S�|IZ3�T0 k� ��(��(2d qD�QC"3Q  ��"    � 3�;,�W<��E� :+�nB��R��"@m�W@���@l�h_8S�|HZ3�T0 k� ��(��(2d qD�QC"3Q  ��"    � 3�;,�XL�E� 9+�nB��R��"@m�W@���@l�h_8S�|HZ3�T0 k� ��(��(2d qD�QC"3Q  ��"    � 3�;,�XL�E�8+�nB��R��"@m�W@���@l�h_4S�|HZ3�T0 k� ��'��'2d qD�QC"3Q  ��"    � 3�;,�XL�E�7+�nB��R��"@m�V@���@l�i_4S�|GZ3�T0 k� ��&��&2d qD�QC"3Q  ��"    � 3�;,�XL�E�6+�nB��R��"@m�V@���@l�i_0S�|GZ3�T0 k� ��%��%2d qD�QC"3Q  ��"    � 3�;,�XL�E�5+�nB��R��#@m�V@���@l�i_,S�|FZ3�T0 k� ��$��$2d qD�QC"3Q  ��"    � 3�;,�YL�E�4+�nB��R��#@m�V@���@l�i_,S�|FZ3�T0 k� ��#��#2d qD�QC"3Q  ��"    � 3�;,�YL�E�3+�nB��R��#@m�V@���@l�j_(S�|FZ3�T0 k� ��"��"2d qD�QC"3Q  ��"    � 3�;,�YL�E�2+�nB��R��#@m�U@���@l�j_(S�|EZ3�T0 k� ��!��!2d qD�QC"3Q  ��"    � 3�;,�YL�E�1+�nB��R��#@m�U@���@l�j_$S�|EZ3�T0 k� �� �� 2d qD�QC"3Q  ��"    � 3�;,�ZL�E�/+�nB��R��#@m�U@���@l�j_$S�|EZ3�T0 k� ����2d qD�QC"3Q  ��"    � 3�;,�ZL�E�.+�nB��R��$@m�U@���@l�k_ S�|DZ3�T0 k� ��"��"2d qD�QC"3Q  ��"    � 3�;,�ZL�E�-�nB��R��$@m�U@���@l�k_ S�|DZ3�T0 k� ��$��$2d qD�QC"3Q  ��"    � 3�;,�Z\�E�,�nB��R��$@m�T@���@l�k_S�|DZ3�T0 k� ��%��%2d qD�QC"3Q  ��"    � 3�;,�Z\�E�+�nB��R��$@m�T@���@l�k_S�|DZ3�T0 k� ��&��&2d qD�QC"3Q  ��"    � 3�;,�Z\�E�*�nBL�R��$@n T@���@l�l_S�|CZ3�T0 k� ��&��&2d qD�QC"3Q  ��"    � 3�;,�[\��E�)�nBL�R��$@n T@���@l�l_S�|CZ3�T0 k� ��&��&2d qD�QC"3Q  ��"    � 3�;,�[\��E�(�nBL�R��$@nT@���@l�l_S�|CZ3�T0 k� ��&��&2d qD�QC"3Q  ��"    � 3�;,�[\��E�'��nBL�R��%@nS@���@l�l_S�|BZ3�T0 k� ��&��&2d qD�QC"3Q  ��"    � 3�;,�[\��E�&��nBL�S��%@nS@���@l�m_S�|BZ3�T0 k� ��*��*2d qD�QC"3Q  ��"    � 3�;,�[\��E�%��nDܼS��%@nS@���@l�m_S�|BZ3�T0 k� ��-��-2d qD�QC"3Q  ��"    � 3�;,�\\��E�$��nDܼS��%@nS@���@l�m_S�|BZ3�T0 k� ��/��/2d qD�QC"3Q  ��"    � 3�;,�\\��E�#��nDܼS��%@nS@���@l�m_S�|AZ3�T0 k� ��0��02d qD�QC"3Q  ��"    � 3�;,�\\��E�#��nD��T��%@nR@���@l�m_S�|AZ3�T0 k� ��1��12d qD�QC"3Q  ��"    � 3�;�\l��A� "��nD��T��%@nR@���@l�n_S�|AZ3�T0 k� ��0��02d qD�QC"3Q  ��"    � 3�;�\l��A� !��nD��T��&@nR@���@l�n_S�|AZ3�T0 k� ��.��.2d qD�QC"3Q  ��"    � 3�;�\l��A��!��nD��T��&@nR@���@l�n_S�|@Z3�T0 k� ��-��-2d qD�QC"3Q  ��"    � 3�;�]l��A�� ��nD��T��&@n R@���@l�n_S�|@Z3�T0 k� ��-��-2d qD�QC"3Q  ��"    � 3�; ]l��A�� K�nD��T��&@n$R@���@l�n_S�|@Z3�T0 k� ��,��,2d qD�QC"3Q  ��"    � 3�; ]l��E\�K�nD��T��&@n$Q@���@l�o_ S�|@Z3�T0 k� ��&��&2d qD�QC"3Q  ��"    � 3�; ]l��E\�K�nD��U��&@n(Q@���@l�o_ S�|?Z3�T0 k� ��!��!2d qD�QC"3Q  ��"    � 3�; ]l��E\�K�nD��U��&@n,Q@���@l�o^�S�|?Z3�T0 k� ����2d qD�QC"3Q  ��"    � 3�;]l��E\�K�nD��U��&@n,Q@���@l�o^�S�|?Z3�T0 k� ����2d qD�QC"3Q  ��"    � 3�;]l��E\�{�nL|�U��'@n0Q@���@l�o^�S�|?Z3�T0 k� ����2d qD�QC"3Q  ��"    � 3�;]l��EL�{�nL|�U��'@n0Q@���@l�o^�S�|>Z3�T0 k� ����2d qD�QC"3Q  ��"    � 3�;]|��EL�{�nL|�U��'@n4Q@���@m p^�S�|>Z3�T0 k� ����2d qD�QC"3Q  ��"    � 3�;]|��EL�{�nL|�U��'@n4P@���@m p^�S�|>Z3�T0 k� ����2d qD�QC"3Q  ��"    � 3�;]]|��EL�{�nL|�U��'@n8P@���@m p^�S�|>Z3�T0 k� ����2d qD�QC"3Q  ��"    � 3�;]]|��EL�{�nL|�U��'@n<P@���@m p^�U;|>Z3�T0 k� ��	��	2d qD�QC"3Q  ��"    � 3�;]]|��A�{�nL|�U��'@n<P@���@mp^�U;|=Z3�T0 k� ��	��	2d qD�QC"3Q  �"    � 3�;]]|��A�{�nL|�U��'@n@P@���@mp^�U;|=Z3�T0 k� ��	��	2d qD�QC"3Q  ��/    � 3�;]] ���A�{�nL|�V��'@n@P@���@mq^�U;|=Z3�T0 k� ����2d qD�QC"3Q  ��/    � 3�;�] ���A�{�nL|�V��(@nDP@���@mq^�U;|=Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;�] ���A�{�nL|�V��(@nDP@���@mq^�U;|=Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;�] ���Gl�{�nL|�V��(@nHO@���@mq^�U;|<Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;�] ���Gl�{�nL|�V��(@nHO@���@mq^�U;|<Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;�]���Gl�{�nL|�V��(@nLO@���@mq^�U;|<Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;�]���Gl���nL��V��(@nLO@���@mq^�@�|<Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]���Gl���nL��V��(@nPO@���@mr^�@�|<Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]���G\���nL��V��(@nPO@���@mr^�@�|<Z3�T0 k� ��	��	2d qD�QC"3Q  ��    � 3�;=]���G\���nL��V��(@nPO@���@mr^�@�|;Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]���G\���nL��V��(@nTO@���@mr^�@�|;Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]��G\���nL��V��(@nTO@���@mr^�@�|;Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]�G\���nL��V��)@nXN@���@mr^�@�|;Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]�GL���nL��V��)@nXN@���@mr^�@�|;Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]�GL���nL��V��)@n\N@���@ms^�@�|;Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]�GL���nL��W��)@n\N@���@ms^�@�|:Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]�GL���nL��W��)@n\N@���@ms^�@�|:Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]�GL���nL��W��)@n`N@���@ms^�@�|:Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]�GL���nL��W��)@n`N@���@ms^�@�|:Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]�GL���nL��W��)@ndN@���@ms^�@�|:Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;=]�GL���nL��W��)@ndN@���@ms^�@�|:Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�GL���nL��W��)@ndN@���@ms^�@�|:Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�	GL|��nL��W��)@nhN@���@ms^�@�|9Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�
GLt��nL��W��*@nhM@���@mt^�@�|9Z3�T0 k� ����2d qD�QC"3Q  ��   � 3�;M]�GLp��nL��W��*@nlM@���@mt^�@�|9Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�GLl��nL��W��*@nlM@���@mt^�@�|9Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�GLh��nL��W��*@npM@���@mt^�@�|9Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�GLd��nL��W��*@npM@���@mt^�@�|9Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�GL`��nL��W��*@npM@���@mt^�@�|8Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�GL\��nL��W��*@ntM@���@mt^�@�|8Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�GL\��nL��W��*@ntM@���@mt^�@�|8Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�GLX��nL��W��*@ntM@���@mu^�@�|8Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�GLT��nL��W��*@nxM@���@mu^�@�|8Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]�GLT��nL��W��*@nxM@���@mu^�@�|8Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]��GLP��nL��W��*@nxL@���@mu^�@�|8Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]��GLL��nL��W��*@nxL@���@m u^�@�|8Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]��GLL��nL��W��*@n|L@���@m u^�@�|8Z3�T0 k� �� �� 2d qD�QC"3Q  ��    � 3�;M]��GLH��nL��W��*@n|L@���@m u^�@�|7Z3�T0 k� �� �� 2d qD�QC"3Q  ��    � 3�;M]��GLH��nL��W��+@n|L@���@m u^�@�|7Z3�T0 k� ��!��!2d qD�QC"3Q  ��    � 3�;M]��GLH��nL��W��+@n�L@���@m u^�@�|7Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]��GLD��nL��W��+@n�L@���@m u^�@�|7Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]��GLD��nL��W��+@n�L@���@m u^�@�|7Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]��GLD��nL��W��+@n�L@���@m v^�@�|7Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M]��GLD��nL��W��+@n�L@���@m$v^�@�|7Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M^l�GL@��nL��W��+@n�L@���@m$v^�@�|7Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M^l�GL@��nL��W��+@n�L@���@m$v^�@�|7Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M^l�GL@{�nL|�W��+@n�L@���@m$v^�@�|7Z3�T0 k� ����2d qD�QC"3Q  ��    � 3�;M^l�GL@{�nL|�W��+@n�L@���@m$v^�@�|7Z3�T0 k� �x�|2d qD�QC"3Q  ��    � 3�;M^l�GL@{�nL|�W��+@n�L@���@m$v^�@�|6Z3�T0 k� �t�x2d qD�QC"3Q  ��    � 3�;M^\�A\@{�nL|�W��+@n�L@���@m$v^�@�|6Z3�T0 k� �p�t2d qD�QC"3Q  ��    � 3�;M^\�A\@{�nL|�W��+@n�L@���@m$v^�@�|6Z3�T0 k� �p�t2d qD�QC"3Q  ��    � 3�;M^\�A\@{�nL|�W��+@n�K@���@m$v^�@�|6Z3�T0 k� �l�p2d qD�QC"3Q  ��    � 3�;M^\�A\@K�nL|�W��+@n�K@���@m(v^�@�|6Z3�T0 k� �h�l2d qD�QC"3Q  ��    � 3�;M^\�A\@K�nBL�W��+@n�K@���@m(v^�@�|6Z3�T0 k� �h�l2d qD�QC"3Q  ��    � 3�;M^\�A�@K�nBL�W��+@n�K@���@m(v^�@�|6Z3�T0 k� �d�h2d qD�QC"3Q  ��    � 3�;M^\�A�@K�nBL�W��+@n�K@���@m(w^�@�|6Z3�T0 k� �d�h2d qD�QC"3Q  ��    � 3�;M^\�A�@K�nBL�W��+@n�K@���@m(w^�@�|6Z3�T0 k� �`�d2d qD�QC"3Q  ��    � 3�;M^\�A�@��nBL�W��,@n�K@���@m(w^�@�|6Z3�T0 k� �X�\2d qD�QC"3Q  �    � 3�;M^̨A�@��n@�W��,@n�K@���@m(w^�@�|6Z3�T0 k� �D�H2d qD�QC"3Q  ��"    � 3�;M^̤ A�@��n@�W��,@n�K@���@m(w^�@�|6Z3�T0 k� �@�D2d qD�QC"3Q  ��"    � 3�;M^̤ A�@��n@�W��,@n�K@���@m(w^�@�|5Z3�T0 k� �<�@2d qD�QC"3Q  ��"    � 3�;=^̠!A�@��n@�W��,@n�K@���@m(w^�@�|5Z3�T0 k� �8�<2d qD�QC"3Q  ��"    � 3�;=^̠!A�@��n@�W��,@n�K@���@m,w^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=^̜"A�@��n@�W��,@n�K@���@m,w^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=^ܜ"A�@��n@�W��,@n�K@���@m,w^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=^ܘ"A�@��n@�W��,@n�K@���@m,w^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=^ܘ#A�@��n@�W��,@n�K@���@m,w^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=^ܔ#A�@� n@�W��,@n�K@���@m,w^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^ܔ$A�@� n@�W��,@n�K@���@m,w^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�$A�@�n@�W��,@n�K@���@m,w^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�%A�@�n@l�W��,@n�K@���@m,w^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�%A�@�n@l�W��,@n�K@���@m,x^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�%A�@�n@l�W��,@n�K@���@m,x^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�&A�@�n@l�W��,@n�K@���@m,x^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�&A�@�n@l�W��,@n�J@���@m0x^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�'A�@� n@l�W��,@n�J@���@m0x^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�'A�@�$n@l�W��,@n�J@���@m0x^�@�|5Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�'A�@�,n@l�W��,@n�J@���@m0x^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�(A�@�0n@l�W��,@n�J@���@m0x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�(A�@�8n@l�W��,@n�J@���@m0x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�(A�@�<n@l�W��,@n�J@���@m0x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�)A�@�Dn@l�W��-@n�J@���@m0x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�)A�@�Hn@��W��-@n�J@���@m0x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�|)A�@�Pn@��W��-@n�J@���@m0x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�|*A�@�Tn@��W��-@n�J@���@m0x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�|*A�@�\n@��W��-@n�J@���@m0x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�x*A�@�dn@��W��-@n�J@���@m0x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�x+A�@�hm@��W��-@n�J@���@m0x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�x+A�@�pm@��W��-@n�J@���@m4x^�@�|4b��T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^�t+A�@�xm@��W��-@n�J@���@m4x^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\t,A�@�|l@��W��-@n�J@���@m4x^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\t,A�@܄l@��W��-@n�J@���@m4y^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\p,A�@܌k@��W��-@n�J@���@m4y^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\p,A�@ܔk@��W��-@n�J@���@m4y^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\p-A�@ܘjA�W��-@n�J@���@m4y^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\p-A�@ܠjA�W��-@n�J@���@m4y^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\l-A�@	��jA�W��-@n�J@���@m4y^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\l.A�@	��jA�W��-@n�J@���@m4y^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\l.A�@	��iA�W��-@n�J@���@m4y^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\h.A�@	��iA�W��-@n�J@���@m4y^�@�|4Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\h.A�@	��iA�W��-@n�J@���@m4y^�@�|4bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\h/A�@
�iA�W��-@n�J@���@m4y^�@�|3bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\h/A�@
�iA�W��-@n�J@���@m4y^�@�|3bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\d/A�@
�iA�W��-@n�J@���@m4y^�@�|3bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\d/A�@
�iA�W��-@n�J@���@m4y^�@�|3bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\d0A�@
�iA�W��-@n�J@���@m8y^�@�|3bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�^\d0A�@��iA�W��-@n�J@���@m8y^�@�|3bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�]\d0A�@��iA�W��-@n�J@���@m8y^�@�|3bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�]\`0A�@��iK��W��-@n�J@���@m8y^�@�|3bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�]\`0A�@��iK��W��-@n�J@���@m8y^�@�|3bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�]\`1A�@��iK��W��-@n�J@���@m8y^�@�|3bs�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�\\`1A�@��iK��W��-@n�J@���@m8y^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�\\\1A�@|�iK��W��-@n�J@���@m8y^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�\\\1A�@|�iK��W��-@n�J@���@m8y^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�\\\2A�@|�iK��W��-@n�J@���@m8y^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�\\\2A�@|�iK��W��.@n�J@���@m8y^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�[\\2A�@|�iK��W��.@n�J@���@m8y^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�[\X2A�@��iK��W��.@n�J@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�[\X2A�@��iK��W��.@n�J@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�[\X3A�@��iK��W��.@n�J@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�[\X3A�@��iK��W��.@n�J@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�Z\X3A�@��iK��W��.@n�I@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=Z\T3A�@��iL�W��.@n�I@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=Z\T3A�@��iL�W��.@n�I@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=Z\T3A�@��iL�W��.@n�I@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=Y\T4A�@��iL�W��.@n�I@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=Y\T4A�@��iL�W��.@n�I@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=Y\T4A�@��hL�W��.@n�I@���@m8z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=X\P4A�@��hL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=X\P4A�@��hL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=X\P4A�@��gL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=W\P5A�@��gL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=W\P5A�@��gL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=W\P5A�@��fL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=W\P5A�@��fL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;=V\L5A�@��fL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MV\L5A�@��fL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MV\L6A�@��fL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MU\L6A�@��fL�W"�.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"   � 3�;MU\L6A�@��fL�W��.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MU\L6A�@��fL�W��.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MU\L6A�@��fL�W��.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MT\H6A�@��fL�W��.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MT\H6A�@��fL�W��.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MT\H7A�@��fL�W��.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MT\H7A�@��fL�W��.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"   � 3�;MS\H7A�@��fL�W��.@n�I@���@m<z^�@�|3Z3�T0 k� �4�82d qD�QC"3Q  ��"   � 3�;MS\H7A�@��fL�W��.@n�I@���@m<z^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MS\H7A�@<�fL�W��.@n�I@���@m<z^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MS\H7A�@<�fL�W��.@n�I@���@m<z^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MR\D7A�@<�fL�W!��.@n�I@���@m<z^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;MR\D7A�@<�fL�W!��.@n�I@���@m<z^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;M R\D7A�@<�fL�W!��.@n�I@���@m<z^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;M R\D8A�@<�fL�W!��.@n�I@���@m<z^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;M R\D8A�@<�fL�W!��.@n�I@���@m<z^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;M Q\D8A�@<�fL�W!��.@n�I@���@m<{^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;M Q\D8A�@<�fL�W!��.@n�I@���@m<{^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;M Q\D8A�@<�fL�W!��.@n�I@���@m<{^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;M Q\D8A�@L�fL�W!��.@n�I@���@m<{^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;M Q\D8A�@L�fL�W!��.@n�I@���@m@{^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;M P\@8A�@L�fL�W!��.@n�I@���@m@{^�@�|2Z3�T0 k� �4�82d qD�QC"3Q  ��"    � 3�;�tS��C��mQ+�Dw�!�/�I�k�C��Da��EQ�LZc�	T0 k� ��L��L2d qD�QC"3Q  ��:    � $ -��tS��C��mQ#�Do�!�/�I�g�C�׈Da��EQ�MZc�	T0 k� ��J��J2d qD�QC"3Q  ��:    � % *��uS��C��mQ�Dg�!�/�I�_�C�ψDa��EQ�MZc�	T0 k� ��I��I2d qD�QC"3Q  ��:    � % '��uS��C��lQ�D_�|/�I�[�C�ǈDa��EQ�MZc�	T0 k� ��G��G2d qD�QC"3Q  ��:    � % $��uS��C��lQ�DW�|/�I�W�C�Da�
�EQ�NZ3�	T0 k� �xF�|F2d qD�QC"3Q  ��:    � & !��vS�C��lQ�C�O�|/�I�O�C�Dax�EQ�NZ3�	T0 k� �tF�xF2d qD�QC"3Q  ��:    � & ��vSw�C��lQ�C�G�|/�I�K�C�Dap�EA�NZ3�	T0 k� �lC�pC2d qD�QC"3Q  ��:    � & ��w�s�C�lQ�C�?�|/�I�G�C�Dah�EA�NZ3�	T0 k� �dA�hA2d qD�QC"3Q  ��:    � & ��w�k�C�lP��C�7�|/�I�C�D��Da`S�EA�OZ3�	T0 k� �\@�`@2d qD�QC"3Q  ��:    � ' �x�[�C�lP��C�'�|/�I�;�D��DaPS�EApOZ3�	T0 k� �L@�P@2d qD�QC"3Q  ��:    � ' �x�O�C�lP��C��|/�I�7�D��D1HS�EAhOZ3�	T0 k� �D?�H?2d qD�QC"3Q  ��:    � ' �y�G�C�l���C��|/�I�3�D{�D1@S�EA`OZ3�	T0 k� �<>�@>2d qD�QC"3Q  ��:    � ' Ӡy�?�C�l���C��|/�I�/�Ds�D18S�EAXOZ3�	T0 k� �4=�8=2d qD�QC"3Q  ��:    � ' Әy�7�C�l���C��|/�I�+�Dk�D10S�EAPOZ3�	T0 k� �,=�0=2d qD�QC"3Q  ��:    � ' Ӑz�/�C�xl���C���|/�I�+�Dc�D1(S�EAHOZ3�	T0 k� �$=�(=2d qD�QC"3Q  ��:    � ' ӈz�'�C�lk���C��|/�I�'�DW�EQS�EA@OZ3�	T0 k� �=� =2d qD�QC"3Q  ��:    � ' 	Ӏz��C�dk���C��|/�I�#�DO�EQS�EA8OZ3�	T0 k� �=�=2d qD�QC"3Q  ��:    � ' �l{��C�Tk��C�י|/�I��D?�EQS�E1(OZ3�	T0 k� �<�<2d qD�QC"3Q  ��:    � ' �d{��ERLk��C�ϙ|/�I��D7�EP�S�E1 OZ3�	T0 k� �;�;2d qD�QC"3Q  ��:    � ' �\|���ERDkP��C�Ǚ|/�I��D/�EP�S�E1NZ3�	T0 k� �:�:2d qD�QC"3Q  ��:    � ' �T|���ER8kP��Eп�|/�C��D'�EP�S�E1NZ3�	T0 k� � :�:2d qD�QC"3Q  ��:    � '���L|���ER0kP��Eз�|/�C��D�EP� S�E1NZ3�	T0 k� � 9�92d qD�QC"3Q  ��:    � '���D}���ER(kP��EЯ�|/�C��D�EP�!S�@�MZ3�	T0 k� ��8��82d qD�QC"3Q  ��:    � '���4}���ERkP��EЛ�|/�C��D�EP�#S�@��LZ3�	T0 k� ��7��72d qD�QC"3Q  ��:    � '���,}���ERkP��E���|/�C��D��EP�$S�@��KZ3�	T0 k� ��6��62d qD�QC"3Q  ��:    � '��� ~���ERkP�E���|/�C���D�E@�%S�@��KZ3�	T0 k� ��5��52d qD�QC"3Q  ��:    � '���~��EQ�kP{�E���|/�C���D�E@�&S�@��JZ3�	T0 k� ��5��52d qD�QC"3Q  ��:    � '���~��EA�kPs�E�{�|/�C���D�E@�'S�E��IZ3�	T0 k� ��5��52d qD�QC"3Q  ��:    � '���~��EA�jPo�E�s�|/�C���C�ێE@�(S�E��IZ3�	T0 k� ��5��52d qD�QC"3Q  ��:    � '����~��EA�j�c�D0c�|/�C���C�ǎE@�)S�E��GZ3�	T0 k� ��4��42d qD�QC"3Q  ��:    � '��2�~��EA�j�[�D0W�|/�C���C࿎E@�*S�E��FZ3�	T0 k� ��5��52d qD�QC"3Q  ��:    � '��2�~��EA�j�S�D0O�|/�C���C෎E@x+S�E��EZ3�	T0 k� ��4��42d qD�QC"3Q  ��:    � '��2�~�EA�i�O�D0G�|/�C���C௎E@p+S�E��DZ3�	T0 k� ��3��32d qD�QC"3Q  ��:    � '��2�~w�EA�i�G�D0?�|/�C���C৏C�d,S�E��CZ3�	T0 k� ��2��22d qD�QC"3Q  ��:    � '��2�~o�EA�iP?�D07�|/�C���C���C�\,S�E��BZ3�	T0 k� ��1��12d qD�QC"3Q  ��:    � '��2�~g�EA�iP7�D0/�|/�C���C���C�T-S�E��BZ3�	T0 k� ��1��12d qD�QC"3Q  ��:    � '��2�}W�C��hP'�D0�|/�C��C���C�@-S�E��@Z3�	T0 k� �x/�|/2d qD�QC"3Q  ��:    � '��2�}O�C��gP�D0�|/�C��C�{�E�8.S�E��?Z3�T0 k� �p.�t.2d qD�QC"3Q  ��:    � '��2�}G�C��gP�D0�|/�D ��C�s�E�,.S�EЀ>Z3�T0 k� �d1�h12d qD�QC"3Q  ��:    � '��2�}?�C��gP�D0�|/�D ��C�k�E�$/S�E�x=Z3�T0 k� �\3�`32d qD�QC"3Q  ��:    � '��2�|3�C�tfP�DO��|/�D ��C�c�E�/S�E�p<Z3�T0 k� �T5�X52d qD�QC"3Q  ��:    � '��B�|+�C�lfP�DO�|/�D ��C�[�E�/S�E�h;Z3�T0 k� �L6�P62d qD�QC"3Q  ��:    � '��B�|#�C�de_��DO�|/�D ��C�S�E�0S�E�d:Z3�T0 k� �D6�H62d qD�QC"3Q  ��:    � '��Bp{�C�Td_��DOם|/�D ��C�?�E��0S�E�T9Z3�T0 k� �45�852d qD�QC"3Q  ��:    � '��Bhz�C�Ld_��DOϝ|/�D �C�7�E��1S�E�L8Z3�T0 k� �05�452d qD�QC"3Q  ��:    � '��B\z�C�Dc_��DOǞ|/�D w�C�/�C��1S�E�D7Z3�T0 k� �(6�,62d qD�QC"3Q  ��:    � '��BTz��C�<c_��DO��|/�D o�C�'�C��1S�E�@6Z3�T0 k� � 5�$52d qD�QC"3Q  ��:    � '��BLy��C�4b_��DO��|/�D g�C��C��2S�E�86Z3�T0 k� �5�52d qD�QC"3Q  ��:    � '��BDy��C�,a_��DO��|/�Dc�D �C��2S�E�05Z3�T0 k� �4�42d qD�QC"3Q  ��:    � '��B<x�߹C�$a_��DO��|/�D[�D �C�2S�E�(4Z3�T0 k� �8�82d qD�QC"3Q  ��:    � '��B4x�׹C�`_��D_��|/�DS�D �C�3S�E� 3Z3�T0 k� �<�<2d qD�QC"3Q  ��:    � '��R,w�ϹC�`_��D_��|/�DK�D��C�3S�E�3Z3�T0 k� ��>� >2d qD�QC"3Q  ��:    � '��R$w�ǸC�__��D_��|/�DC�D�C�3S�E�2Z3�T0 k� ��@��@2d qD�QC"3Q  ��:    � '��RvῸC� ^_��D_��|, E�;�D�C�4S�E�2Z3�T0 k� ��A��A2d qD�QC"3Q  ��:    � '��Ru᫷C��]_��D_w�|, E�+�E�ےC�4S�E��1Z3�T0 k� ��A��A2d qD�QC"3Q  ��:    � '��Rt᣷C��\_��D_o�|, E�#�E�ϒC�x5S�A��1Z3�T0 k� ��@��@2d qD�QC"3Q  ��:    � '��Q�tᛷC��[_��D_g�|, E��E�ǒC�p5S�A��0Z3�T0 k� ��?��?2d qD�QC"3Q  ��:    � '��Q�sᓷC��[O��D__�|, E��EￒC�d5S�A��0Z3�T0 k� ��=��=2d qD�QC"3Q  ��:    � '��Q�r�C��ZO��D_S�|, E��E﷓C�\5S�A��0Z3�T0 k� ��=��=2d qD�QC"3Q  ��:    � '��Q�r�C��YO��D_K�|,D?��EﯓC�P6S�A��/Z3�T0 k� ��<��<2d qD�QC"3Q  ��:    � '��Q�q�{�C��XO�DoC�|,D?��E陸C�H6S�A��/Z3�T0 k� ��<��<2d qD�QC"3Q  ��:    � '��Q�p�g�EаWOo�Do3�|,D?��EC�47S�A��/Z3�T0 k� ��;��;2d qD�QC"3Q  ��:    � '��Q�p�_�EШV�g�Do+�|,D?��EC�,7S�A��/Z3�T0 k� ��;��;2d qD�QC"3Q  ��:    � '��Q�o�W�EРU�_�Do#�|,D?��D?��C� 7S�A��/Z3�T0 k� ��;��;2d qD�QC"3Q  ��:    � '���o�O�EИT�[�Do�|,D?��D?{�C�7S�A��/Z3�T0 k� �x;�|;2d qD�QC"3Q  ��:    � '���n�G�EАT�S�Do�|,D?��D?s�C�8S�A��/Z3�T0 k� �p;�t;2d qD�QC"3Q  ��:    � '���n�?�EЈS�G�Do�|,D?��D?k�D8S�Aϔ/Z3�T0 k� �d;�h;2d qD�QC"3Q  ��:    � '���m�7�EЀR�;�Do�|,D?��D?c�D�8S�Aό/Z3�T0 k� �\;�`;2d qD�QC"3Q  ��:    � '���m/�E�xQ�/�Dn��|,D?��E�[�D�8S�Aτ/Z3�T0 k� �T;�X;2d qD�QC"3Q  ��:    � '���|l�E�hP� Dn�|,D?��E�K�D�9S�A�t/Z3�T0 k� �D;�H;2d qD�QC"3Q  ��:    � '���tk�C�`O�D>�|,DO��E�C�D�9S�A�l/Z3�T0 k� �<<�@<2d qD�QC"3Q  ��:    � '���lk�C�XO��D>߲|,DO��E�7�D�9S�A�d0Z3�T0 k� �4<�8<2d qD�QC"3Q  ��:    � '���dj�C�PN��D>׳|,DO��E�/�D�9S�A�\0Z3�T0 k� �,<�0<2d qD�QC"3Q  ��:    � '���\j ��C�HM��D>ϴ|,DO�E�'�D�:S�A�X0Z3�T0 k� �$<�(<2d qD�QC"3Q  ��:    � '���Tj �C�@M��D>ǵ|,DOw�E��D�:S�A�P0Z3�T0 k� �<� <2d qD�QC"3Q  ��:    � '���Li �C�8L��
D>��|,I�o�E��D�:S�A�H0Z3�T0 k� �=�=2d qD�QC"3Q  ��:    � '���Di ߲C�0L��D>��|,I�k�E��D�:S�A�@1Z3�T0 k� �>�>2d qD�QC"3Q  ��:    � '���0h ϱC� J��D>��|,I�_�E���D�;S�A�01Z3�T0 k� ��?��?2d qD�QC"3Q  ��:    � '���(hǱC�J��D>��|,I�W�E���D|;S�A�(2Z3�T0 k� ��@��@2d qD�QC"3Q  ��:    � '��� g��C�I��D>��|,I�S�E��Dt;S�A� 2Z3�T0 k� ��@��@2d qD�QC"3Q  ��:    � '���g��C�I��D>��|,I�K�E��Dl;S�A�2Z3�T0 k� ��A��A2d qD�QC"3Q  ��:    � '���f��C� H��DN��|,I�G�E��D`<S�A�3Z3�T0 k� ��A��A2d qD�QC"3Q  ��:    � '�~�f��C��G��DN��|,I�C�E�ۤDX<S�A�3Z3�T0 k� ��A��A2d qD�QC"3Q  ��:    � '�|� f��C��G�|DN{�|,I�?�E�ӥDL<S�A� 4Z3�T0 k� ��B��B2d qD�QC"3Q  ��:    � '�z��e��C��F�tDNs�|,I�;�E�ϦDD<S�A��4Z3�T0 k� ��B��B2d qD�QC"3Q  ��:    � '�x �d��C��E�`DNc�|,I�/�F��D0=S�A��5Z3�T0 k� ��C��C2d qD�QC"3Q  ��:    � '�v �d{�C��E�XDN[�|,I�+�F��C�(=S�A��5Z3�T0 k� ��D��D2d qD�QC"3Q  ��:    � '�t �ds�C��D�PDNS�|,I�'�F��C�=S�A��6Z3�T0 k� ��D��D2d qD�QC"3Q  ��:    � '�r �c�g�C��D�HDNO�|,I�#�F��C�=S�A��6Z3�T0 k� ��E��E2d qD�QC"3Q  ��:    � '�p �c�_�C��C	~@DNG�|,I�#�F��C�=S�A��7Z3�T0 k� ��E��E2d qD�QC"3Q  ��:    � '�n �c�W�C��C	~8DN?�|,I��F��C� =S�A��8Z3�T0 k� ��F��F2d qD�QC"3Q  ��:    � '�l �b�O�D�B	~0!D^7�|,I��F��I��=S�A�8Z3�T0 k� ��G��G2d qD�QC"3Q  ��:    � '�j �b�G�D�B	~(!D^/�|,I��F��I��=�A�9Z3�T0 k� �xG�|G2d qD�QC"3Q  ��:    � '�h �b�?�D�A	~ "D^'�|,E_�F��I��=�A�9Z3�T0 k� �pH�tH2d qD�QC"3Q  ��:    � '�f �a�+�D�@	~$D^�|,E_�F��I��=�A�;Z3�T0 k� �dI�hI2d qD�QC"3Q  ��:    � '�d�a�#�Dx@	�%D^�|,E_�F��I��=�A�;Z3�T0 k� �\J�`J2d qD�QC"3Q  ��:    � '�b�a��Dp?	�&D^�|,E_�E���I��=�A��<Z3�T0 k� �XI�\I2d qD�QC"3Q  ��:    � '�`x`��Dh?	� &D^�|,E_�E���I��=�A��<Z3�T0 k� �PI�TI2d qD�QC"3Q  ��:    � '�^p`��D`>	��'D]��|,E^��E���I��=�A��=Z3�T0 k� �HJ�LJ2d qD�QC"3Q  ��:    � '�\h`��DX>	��(D]��|,E^��E��I��=�A�x>Z3�T0 k� �@J�DJ2d qD�QC"3Q  ��:    � '�Z`_���DP>	}�(D]��|,E^��E�{�C�=�A�t?Z3�T0 k� �<K�@K2d qD�QC"3Q  ��:    � '�XL_��D<=	}�)Dm��|,E^��E�w�C�=�|A�d@Z3�T0 k� �0L�4L2d qD�QC"3Q  ��:    � '�VD_�߭D4<	}�*Dm��|,C���E�w�C�=�xA�\AZ3�T0 k� �(M�,M2d qD�QC"3Q  ��:    � '�T<^�׭D,<	}�*Dm��|,	C���E�s�C�=�tA�TAZ3�T0 k� � N�$N2d qD�QC"3Q  ��:    � '�R4^�ϬD$<	��+Dm��|,	C���E�s�C�=�pA�LBZ3�T0 k� �O�O2d qD�QC"3Q  ��:    � '�P�,^�ǬD;	��+Dm��|,	C���E�s�C�=�pA�HCZ3�T0 k� �O�O2d qD�QC"3Q  ��:    � '�N�$]���D;	��+Dm���,	C���E~o�C�x=�lA�@DZ3�T0 k� �P�P2d qD�QC"3Q  ��:    � '�L�]���D:	��,Dm���,	C���E~o�C�h=�dA�0EZ3�T0 k� ��R� R2d qD�QC"3Q  ��:    � '�J�]��D�:	}�,Dm���,
C���E~k�C�`=�`A�(FZ3�T0 k� ��S��S2d qD�QC"3Q  ��:    � '�H� \��D�9	}�,Dm���,
C��E~k�C�X=�\A�$GZ3�T0 k� ��S��S2d qD�QC"3Q  ��:    � '�G��\��C��9	}�,D=���,C��E~k�E�P=�XA�HZ3�T0 k� ��T��T2d qD�QC"3Q  ��:    � '�F��\��C��9	}�-D=���,C��E~k�E�H=�TA�HZ3�T0 k� ��U��U2d qD�QC"3Q  ��:    � '�E��[w�C��8M�-D=���,C��E~g�E�8=LA�JZ3�T0 k� ��W��W2d qD�QC"3Q  ��:    � '�D��[o�C��8M�.D={��,C���E~g�E�,=HA� KZ3�T0 k� ��X��X2d qD�QC"3Q  ��:    � '�C��[g�C��7M�.D=s��,C���E~c�E�$=@A��LZ3�T0 k� ��Y��Y2d qD�QC"3Q  ��:    � '�B��[_�C�7M�.I�o��,C���E~c�E�=<A��MZ3�T0 k� ��Y��Y2d qD�QC"3Q  ��:    � '�A��[W�C�7M�/I�g��,C���E~c�E�=8A��NZ3�T0 k� ��[��[2d qD�QC"3Q  ��:    � '�@��ZO�C�6=�0I�_��,C���Enc�E�=0A��OZ3�T0 k� ��]��]2d qD�QC"3Q  ��:    � '�?��Z;�C�6=�1I�S��,C�s�En_�E��=(A��PZ3�T0 k� ��_��_2d qD�QC"3Q  ��:    � (�>��Z3�C�5=�2I�O��(C�k�En_�E��= A��Qbs�T0 k� ��`��`2d qD�QC"3Q  ��:    � )�=��Z+�C��5=�2I�K��(C�c�En[�E��=A��Rbs�T0 k� ��a��a2d qD�QC"3Q  ��:    � *�<��Y#�C�|5M�3I�C��(C�_�EnW�E��>E]�Sbs�T0 k� ��\��\2d qD�QC"3Q  ��:    � +�;�xY�C�l4M�5I�;��(C�L EnW�E��>E]�Ubs�T0 k� ��Y��Y2d qD�QC"3Q  ��:    � ,�:�pY�C�`4M|6I�7��$DDEnS�E�> E]�Vbs�T0 k� ��V��V2d qD�QC"3Q  ��:    � -�9hY��I�\4Mx7I�/��$D<EnO�E�>�E]�Wbs�T0 k� �|T��T2d qD�QC"3Q  ��:    � .�8`X��I�T3�t8I�+��$D4EnK�E�>�E]�Wbs�T0 k� �xS�|S2d qD�QC"3Q  ��:    � /�8PX�I�D3�l;I�#��$D(En?�E�?�E]�Ybs�T0 k� �hS�lS2d qD�QC"3Q  ��:    � 0�8DX�ߩI�<3�h<I���$DE^;�E�?�E]�Zbs�T0 k� �dS�hS2d qD�QC"3Q  ��:    � 1�8<X�שI�43�d=E���$DE^7�E�@�E]�[Z3�T0 k� �\S�`S2d qD�QC"3Q  ��:    � 2�84W�ϩI�03�`>E���$DE^/�E�x@�E]x\Z3�T0 k� �TS�XS2d qD�QC"3Q  ��:    � 3�8$WI�$3�TAE���$D�E^'�E�dA��E]l]Z3�T0 k� �HT�LT2d qD�QC"3Q  �:    � 3�8WI�3�PBE���$D�	C��E�\A�E]d^Z3�T0 k� �LT�PT2d qD�QC"3Q  ��?    � 3�8WI�3�LDE����$D�
C��E�TB�E]\_Z3�T0 k� �PT�TT2d qD�QC"3Q  ��?    � 3�8WI�3=DEE���� D�
C��E�HC�EMT_Z3�T0 k� �TS�XS2d qD�QC"3Q  ��?    � 3�8�VI�3=<HE���� D�C��E�8D�EMDaZ3�T0 k� �XS�\S2d qD�QC"3Q  ��?    � 3�8�VI� 3=8JE���� D�C���D�0E�EM<aZ3�T0 k� �\R�`R2d qD�QC"3Q  ��?    � 3�8�V��E��3=0KE�� � D�C���D�(F�EM4bZ3�T0 k� �\R�`R2d qD�QC"3Q  ��?    � 3�8�V�w�E��2],LE��� D�C���D�G�EM0bb��T0 k� �`R�dR2d qD�QC"3Q  ��?    � 3�8�V�o�E��2](NE��� D�C���D�H�xEM(cb��T0 k� �dR�hR2d qD�QC"3Q  ��?    � 3�8�U�_�E��2] PE��� D�C���D�J�dEMcb��T0 k� �hQ�lQ2d qD�QC"3Q  ��?    � 3�8�U�W�E��1]RE��� D�C�� E��K�\EMdb��T0 k� �lQ�pQ2d qD�QC"3Q  ��?    � 3�8�U�O�E��1mSE��� EݔC��E��L�TEMdb��T0 k� �pQ�tQ2d qD�QC"3Q  ��?    � 3�8�U�C�E��1mTE��	� E݌C��E��M�Le} db��T0 k� �pP�tP2d qD�QC"3Q  ��?    � 3�8�U�;�E��1mTE��� E݄C��E��N�De|�eb��T0 k� �tP�xP2d qD�QC"3Q  ��?    � 3�8�T	�+�Eݴ0mVE��� E�tC��E��Q�4e|�fb��T0 k� �xP�|P2d qD�QC"3Q  ��?    � 3�8�T	�#�Eݬ0mWIܨ� E�lC��E��R�(e|�gb��T0 k� �|O��O2d qD�QC"3Q  ��?    � 3�8�T	��Eݨ0m XIܤ� E�dE]�E��T� e|�gZ3�T0 k� ��O��O2d qD�QC"3Q  ��?    � 3�8�xT	��Eݠ0l�XIܠ� E�\E]�E��U�e|�hZ3�T0 k� ��O��O2d qD�QC"3Q  ��?    � 3�8�pT	��E�0\�YIܜ� E�TE]�E��W�e|�iZ3�T0 k� ��O��O2d qD�QC"3Q  ��?    � 3�8�`T	���E�0\�[Iܔ� E�DE]xE��Z� e|�jZ3�T0 k� ��L��L2d qD�QC"3Q  ��"    � 3�8�XT	���E�/\�[I�� E�<E]pF�[�e|�jZ3�T0 k� �tJ�xJ2d qD�QC"3Q  ��"    � 3�8	�PS	��E�x/\�\I��$E�4E]h	F�]�e|�kZ3�T0 k� �hH�lH2d qD�QC"3Q  ��"    � 3�8	�HS	��I�p/��]I��$E�,E]`	F�_�e|�kZ3�T0 k� �\E�`E2d qD�QC"3Q  ��"    � 3�8	�8S	�ߨI�d/��^I��$E�E]PF�b�e|�mZ3�T0 k� �LC�PC2d qD�QC"3Q  ��"    � 3�8	�0S	�ۨI�\/��_E|��$E�E]HF�b�e|�mZ3�T0 k� �@A�DA2d qD�QC"3Q  ��"    � 3�8	�(S	�ӨI�X/��`E||�(E�E]@F�c�e|�nZ3�T0 k� �8@�<@2d qD�QC"3Q  ��"    � 3�8	�$S	�ϨI�P/��aE||�(E�E]8F�c�e|�nZ3�T0 k� �4?�8?2d qD�QC"3Q  ��"    � 3�8	�S	�˨I�L/��bE|x�(E�  EM0F�c�e|�oZ3�T0 k� �,>�0>2d qD�QC"3Q  ��"    � 3�8	�S	���I�@/��dE|t"�(E��"EM F�d�e|tpZ3�T0 k� �$>�(>2d qD�QC"3Q  ��"    � 3�8	�S	���I�</̼eE|p#!�(E��#EME��e�e|ppZ3�T0 k� �>� >2d qD�QC"3Q  ��"    � 3�8	�S	���I�8/��fE|l$!�(E��$EME��e�e|hqZ3�T0 k� �>�>2d qD�QC"3Q  ��"    � 3�8	��S	���I�0/��gE|l&!�(E��%EME��f�e|dqZ3�T0 k� �>�>2d qD�QC"3Q  ��"    � 3�8	��S	���I�,/��iE|h'!�(E��&EL�E��f�e|\rZ3�T0 k� �>�>2d qD�QC"3Q  ��"    � 3�8	��S	���I�$/��kEld*!�(E��)EL�E��gle|TsZ3�T0 k� �>�>2d qD�QC"3Q  ��"    � 3�8	��S	���I� /̘lEl`+!�(E��*EL�E��gde|LsZ3�T0 k� � >�>2d qD�QC"3Q  ��"    � 3�8	��S	���I�/̔nEl\-!�(F�+EL�E��h\e|HsZ3�T0 k� ��>� >2d qD�QC"3Q  ��"    � 3�8	��S	���I�/̌oEl\.!�(F�,EL�E��hTe|@tZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�8	��S	���I�/̈pElX0!�(F�.E<�E��iLe|<tZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�8	��S	���I�/̈pElP3!�(F�0E<�E��i<e|0uZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�8	��S	���I�/̄qElP4�(F�2E<�E��j�0EL,vZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�8	��S	���I�/̀sE|L5�(F�3E<�E��j�(EL$vZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�8	��S	���I�/�tvE|H8�(F�6E<�E��j�ELxZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�8	��S	���I� /�lwE|H9�(F�7CL�E��i�ELyZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�8	��S	���I� /�`xE|D9�(F�9CL�E��i�E<yZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�8	��S	���I��/�`xE|D:�(F�9CL�E��i� E<yZ3�T0 k� ��>��>2d qD�QC"3Q  �"    � 3�8	��S	���I��/�TxE|<<�(F�<CLtE��g��E<xZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�9	��S	���I��/\PxE|8=�(E��>CLpB��g��E<wZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�:	��S	���I��/\HxE|8=�(E��?CLhB� f��S��wZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�;	��S	���I��/\DyE�4>!�(E�|ACLhB�e��S��vZ3�T0 k� ��>��>2d qD�QC"3Q  �"    � 3�;	��S	��I��0\<yE�0?!�$E�xD@�`
B�dP�S��vZ3�T0 k� ��>��>2d qD�QC"3Q  �"   � 3�;	��S	��I��0\8yE�,@!� E�xF@�`	@lcP�S��uZ3�T0 k� ��>��>2d qD�QC"3Q  ��"    � 3�;�S]�E��0\0yE�(@!� E�xG@�\	@lcP�S��uZ3�T0 k� ��@��@2d qD�QC"3Q  ��"    � 3�;�S]{�E��0\(zF$B!�E�tJ@�T@laP�S��tZ3�T0 k� ��B��B2d qD�QC"3Q  ��"    � 3�;�S]w�E��0\$zF$C!�E�tL@�P@laP�S��sZ3�T0 k� ��C��C2d qD�QC"3Q  ��"    � 3�;�S]s�E��1\ yF$C!�E�tM@�P@l `P�S��sZ3�T0 k� ��D��D2d qD�QC"3Q  ��"    � 3�;�SMs�E��1\xF D!�E�tO@�L@l `P�S��sZ3�T0 k� ��E��E2d qD�QC"3Q  ��"    � 3�;�SMo�E��1\xF E!�E�tP@�H@l$_P�S��rZ3�T0 k� ��E��E2d qD�QC"3Q  ��"    � 3�;�SMk�E��2\wE� F�E�tR@�D@l(^P|S��rZ3�T0 k� ��F��F2d qD�QC"3Q  ��"    � 3�;�SMg�E��3\vE� G�E�tT@�@@l,]PlS��pZ3�T0 k� ��G��G2d qD�QC"3Q  ��"    � 3�;��S�c�M\�4\vE� H�E�tV@�<@l0]PhS��oZ3�T0 k� ��E��E2d qD�QC"3Q  ��"    � 3�;�|S�c�M\�4\uE� I�E�xW@�<@l4\P`S��nZ3�T0 k� ��D��D2d qD�QC"3Q  ��"    � 3�;�tS�_�M\�5\tB� J�E�xX@�8 @l8[PXS��nZ3�T0 k� ��D��D2d qD�QC"3Q  ��"    � 3�;�pS�_�M\�5\tB� J�E�xZ@�4 @l8[PPS��mZ3�T0 k� ��C��C2d qD�QC"3Q  ��"    � 3�;�lS�[�M\�6\sB� K�E�|[@�7�@l<ZPLS��lZ3�T0 k� ��C��C2d qD�QC"3Q  ��"    � 3�;�dS�W�M\�6\ sB� K� E�|\@�3�@l<ZPDS��kZ3�T0 k� ��C��C2d qD�QC"3Q  ��"    � 3�;�`S�W�M\�7[�rB� K� E��^@�/�@l@ZP<S��jZ3�T0 k� ��D��D2d qD�QC"3Q  ��"    � 3�;�XS�S�M\�8[�rB� K� E��_@�/�@l@ZP8S��jZ3�T0 k� ��D��D2d qD�QC"3Q  ��"    � 3�;�TS�S�M\�8[�qB� K��E��`@�+�@lDZP0S��iZ3�T0 k� ��E��E2d qD�QC"3Q  ��"    � 3�;�HS�O�M\�9[�pB�$L��E��b@�'�@lHZP$S��hZ3�T0 k� ��F��F2d qD�QC"3Q  ��"    � 3�;	�@SK�Ml�:[�pB�$L��E��c@�#�@lLZPS��gZ3�T0 k� ��G��G2d qD�QC"3Q  ��"    � 3�;	�<SG�Ml�:[�pB�(L��E��d@�#�@lPZPS��fZ3�T0 k� ��I��I2d qD�QC"3Q  ��"    � 3�;	�4SG�Ml�;[�oB�(L��B��e@��@lTZPS��eZ3�T0 k� ��J��J2d qD�QC"3Q  ��"    � 3�;	�0SC�Ml�;[�oB�,L��B��f@��@lTZPS��eZ3�T0 k� ��K��K2d qD�QC"3Q  ��"    � 3�;	�,SC�Ml�<[�oB�,L��B��g@��@lX[PS��dZ3�T0 k� ��K��K2d qD�QC"3Q  ��"    � 3�;	�$S?�Ml�<[�oB�,L��B��h@��@l\[P S��cZ3�T0 k� ��L��L2d qD�QC"3Q  ��"    � 3�;	� S?�Ml�=[�nB�0L��B��h@��@l\[_�S��cZ3�T0 k� ��L��L2d qD�QC"3Q  ��"    � 3�;	�S;�Ml�=[�nB�4L��B��i@��@l`[_�S��bZ3�T0 k� ��M��M2d qD�QC"3Q  ��"    � 3�;	�S;�Ml�=[�nB�8L��B��j@��@ld[_�S��bZ3�T0 k� ��M��M2d qD�QC"3Q  ��"    � 3�;	�S7�M\�>[�nB�8L��B�i@��@ld[_�S��aZ3�T0 k� ��M��M2d qD�QC"3Q  ��"    � 3�;                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��^� ]�(V(U 8 �� P��   � �	    ��H��     Q��H��    �i   	        _		 Z�;           ���    ���   0		 
 
          8�;     
	  ���O     8�V��    ���            � �1          �     ���    	!
           8�         ��     8���           	      �) �
         �      ���   H
           fG�   � �	    �?K�     fG��?K�           
           N		 Z�;          �0�  %  ���  0	 

          W��  � �     .�2�     W���2�                     v
	 Z�;          ��    ���   @	
           .�        B���
     .ׯ���
     3                      ���.              �  ���    8

 '             I��       V����     I�����4    �� �                � ��        �@     ��H   H
D
 
          �Ҹ�        j����    �Һ�����    ��             
   �         �     ��@   (
 
           {E        ~�P�     {�P �     O i               e �         �      ��@   0	
           ��          ���Y�     ����^l      ��               
  ��         	 !�     ��@   H	$
          2��       ����o     2�2���o    ��               
     �         
 h�     ��B   03 
           ����
	      � �ث     �� �ث                              ���              �  ��@   P		 5                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          o�  ��        ��҇     o��҇         "                  x                j  �       �                              ��        ��         �                                                            �                         �H���?�2�������P���� ����� 
   	             
  C   � �� ���K       �D �c@ �D d@ �d  d` ɤ  d� �� d� Ǆ  \� �� ]  �� ]  �  ]@ 
�\ W  �D f� �d g  Є g  Ф g@���� � �� �[� �� \� H� _� 
�� V� 
�\ W  
�� W� 
�� W� 
�\ W� � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }`���� ����� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����;�� 3�� �  ������  
�fD
��L���"����D" � j  "  B   J jF�"      �j * , .��
��
��"   "D�j�
�� " �
� �  �  
�      ��     ��           ��     ��       I    ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �"D      ��m �  ���        � �  ��        �        ��        �        ��        �    ��    (�� =��        ��                         襩 4  ����                                     �                 ����             ����%��   3�;                 10 Dale Hawerchuk                                                                                   3  3      � �
�	4k� �L k� �"kj �: kr �� �� �*CB �	CF �
CJ � � � �K � K �B� �% B� �K. �K6& � K9  � K: �C- � C"3 �C#& �C%. � C'6 �B� � B� �B� �B� � B�! �k~? � k�/ l!c� � � "c� � d#kV r$k^ �&%"� �& &"� �'� �(
� �&)"� �& *"� �+"� �,*� � �-"�
 � ."� w/� w0
� �1)�} � 2*Om � 3*Km � 4*J} �5)�m6)�}; 7*IUK 8*PES 9*O][  *HES  *R][ <*Ge[  *KE[  *KE;  *LU                                                                                                                                                                                                                         �� R         �     @         �     ^ P E `  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    ��4�� ��������������������������������������������������������   �4, B� 0 � �� ��@2�@Y�J���x����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   l  	  +        0$�J      h                             ������������������������������������������������������                                                                                                                                         �    ���                      ��                  
   �� ��������������������� � ������������ �� �������������� ����������� ������ ���������������� � ����� �����  ��� �������� �������� ��������������� ������� �������� � ������� ������ ��������� ����������������������������� ����                                   �    +    ��  D��J      	e  	                           ������������������������������������������������������                                                                                                                                           �    ���i                      �  �            
 	    �� �������������������� � ���� �������������� ����������� ������������������������������������������ ������� ��������������� � ��������������������������������� ������ ������������ ������ �������� ���������������� ��������������������� �  �������                                                                                                                                                                                                                                                                                                                           �             


            �   }�         ���z        8�      0�                                   R
                         ���F��������  >      6�������������������������������������������������  �����  6���������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 8 F <                                  � !�� �\                                                                                                                                                                                                                                                                                       
)n1n  1�1n                a      `      a      a                  m                                                                                                                                                                                                                                                                                                                                                                                                                
@ h  	>�  J�  M#�  J#�  EZm�  �N )�UJ��������˖���˖�������˖�v����n�                       � i          �   &  AG� �   �                    �                                                                                                                                                                                                                                                                                                                                        7 H   �          #             !��                                                                                                                                                                                                                            Y   �� �� Ѱ��      �� I      �� ��������������������� � ������������ �� �������������� ����������� ������ ���������������� � ����� �����  ��� �������� �������� ��������������� ������� �������� � ������� ������ ��������� ����������������������������� ������ �������������������� � ���� �������������� ����������� ������������������������������������������ ������� ��������������� � ��������������������������������� ������ ������������ ������ �������� ���������������� ��������������������� �  �������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ?      3                             I     �  �����J����      ��     p�      �         �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �� ��  � ��     � ��   	 ��  p �� �� ��     -�  �@  'l >�������J J  'l -�  �@  'l   )  �1   �    ��    ��  � �� ��   �z � �N ��  � �� ��   	 �� �� ��  �� �� �  �� �� �z � ��� �$  �  �� �       �   d   ���� e�����  g��� 	       f ^�         �� B 3            ��_R���2�������J����  ��      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                                                         �� �����虙������(��������������񙙘�!                �  �������                           �       �  "(� """ �"" ""  "   �      �   �"��"""�"""�"""�"""�����������������������������������""�".�"/��"���!���.���/���-���""����������.���-������/�������   ��  �  .� /�� "�� "� "-�                                ""�  �(��""! ("" �"  �"   ����������������陙����.��� 陙/���.���"���"!��"��".���!♒""����������������̎���""�""",""/ �-� /� "�� "�� . /� �                    �                                           ""陂".��""� � �          �"(��(""������� ��        ""!�"!������������           ��     �                       wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  ""   "! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  ""   "! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �            " ""   ""     " ""   "" "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                          �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                            �  �˰ ��� �wp ���                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                    ""  ."  �"    �   ��  �   �                  �  �  �  �                                       �  �   ��                     �    � �  ��                  ���                                                                                                                                                                          �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                                � ���             �  �� �  �� �  ��                        �              ����������             �� �  �  �      �   �                             ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                      �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                                  � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         "  " �" ��" ��- �ۼ w۽��ݹ����� ��� ��  ˼  ��  ˼  ��  H�  �D  J�  J�  �  �  �  �  
�  �  �  �  ,�  " "" �" �"�   ˰  ��  wp ��ډ�v���r�̸��˰��� ��  ��  ��  ��  ̸  ��  ��  DC  C4@ T4@ T40 T30 T30 S;� H�  ��  ��  ��  ""  "  �""� "�/��        �   �   �      �  �   �   �   �   �              �   �   �   �             ���� �                        " "" """ �"  �   �   �                              � ��                  �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                   UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �           J� �D�M�D���4���ˠ ��� ̽� ��� ��ٰ�۰"˰""+�""!��"�  �                        �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H��        �� ��� ۻ� }݉ ��� ��� ��� �˼ ��� �ٚ��ک��М��J� "                           � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �                        �� ̻ ��   �������  �                     �  �   �  �  ��  �  ��  �                                                                                                                                                                                                                          	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                   �   ������  ��                      �   �                      �������  ���    �                    �   ���                       ���                � �������������               �  �     �   �  �  �                                                                                                                  �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                             �� ��������p��}`     �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��  ��  ���  �   ��  ��  ��  �  �   ��  ��                                                                                                                                                                                       	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                       ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ���          �  ��� ݼ� w{� �װ vw�                    �   ���                            �   �                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                            �� ̽      D   J   J   J  �  ��  ��  ʘ ̠ "  " �"" �""  �"                      �    ���� �              �  �� ��  �    � ���                                  � �������������  �                                                                                                                                                      �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                             �  ��� ܽ� ��p �}`�   �   �      �                                � �� ���H���     ̰ �˻���ݹ��w���&ɧvvɪ�p              �  �� �� �� ��                         ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                           �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��                  �          �         �   �  �  �   �               �   �                               � ����ݼ� ����                                                                                                                                                                             �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""��������D�M����""""�������D�M�M""""�����AMAD������""""��������D��""""������MM�����""""���������D�""""������������������""""������������������������"""$���4���4���4���4���4���4ffffffffffffffffff333DDDffffffffffffffffffffffff3333DDDDafaafffaffDDffff3333DDDDfFfFDfFFfFffdFffff3333DDDDfaffaffaffafffDfffff3333DDDDADAFaFadFfDffff3333DDDDafffDfdFdffff3333DDDDDDFFDfFFfdFffff3333DDDDAffAffaffafffDffffff3333DDDDffffffffffffffffffffffff3333DDDDfff4fff4fff4fff4fff4fff43334DDDD"""������������������""""������������������������""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""���������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��������������D�����3333DDDDI����D��DI����3333DDDDADAIA����D������3333DDDD��������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(����������������� � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(����������������� 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5���������������� x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x���������������� w w x y�������H���������������������������������H������yxww����������������  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(���������������� , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,���������������� +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+���������������� 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5���������������� =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=����������������     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( ���������������� � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � ����������������� � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � ����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
�	4k� �L k� �"kj �: kr �� �� �*CB �	CF �
CJ � � � �K � K �B� �% B� �K. �K6& � K9  � K: �C- � C"3 �C#& �C%. � C'6 �B� � B� �B� �B� � B�! �k~? � k�/ l!c� � � "c� � d#kV r$k^ �&%"� �& &"� �'� �(
� �&)"� �& *"� �+"� �,*� � �-"�
 � ."� w/� w0
� �1)�} � 2*Om � 3*Km � 4*J} �5)�m6)�}; 7*IUK 8*PES 9*O][  *HES  *R][ <*Ge[  *KE[  *KE;  *LU3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������=�K�K�S�[��<�K�R�G�T�T�K� � � � � � � �=��;�������������������������������������������+�R��7�G�I�3�T�T�O�Y� � � � � � � � � ��=�@�������������������������������������������.�G�R�K��2�G�]�K�X�I�N�[�Q� � � � � � ��=�@�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������=��;� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ������������������=�@� �� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 