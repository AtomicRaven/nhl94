GST@�                                                            \     �                                                     @                    ���2�����	 ʴ������̸������z���        �h      #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"     �j@ �    ��
  �                                                                               ����������������������������������      ��    bb= QQ0 4 111 44              		 

                     ��� �   � �                 nnE ))         88�����������������������������������������������������������������������������������������������������������������������������o  b  o   4  +c  c  'c            �        	  
      	G  7�  V(  	(                  n  1          :8 �����������������������������������������������������������������������������                                (  0   |  S�   @  #   �   �                          �                                                     '        )n)nE  1n    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE 0 �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ߾@ k� x l��Y| K���K�A[��-��^;�3��T0 k� ����c�t B%�0d    ��?    ����@߾@ g� | l��Y| K���K�A[��-��^3�3��T0 k� ����c�t B%�0d    ��?    ����@߾@ g� | l��Y| K���K�A[��-�^/�3��T0 k� ����c�t B%�0d    ��?    ����@߾@ g� | l��Y| K���K�A[��-{�^'�3��T0 k� ����c�t B%�0d    ��?    ����@߿@ g� | l��Y| K���K�A[��-s�^#�3��T0 k� ����c�t B%�0d    ��?    ����@߿@ c� | l��Y| K���K�A\�-o�^�3��T0 k� ����c�t B%�0d    ��?    ����@߿@ c� | l��Y{�K���K�A\�-k�^�3��T0 k� ����c�t B%�0d    ��?    ����@߿@ c� | l��Y{�K����K�A\�-c�^�3��T0 k� ����c�t B%�0d    ��?    ����@߿@ c� | l��Y{�K����K�A\�-_�^�3��T0 k� ����c�t B%�0d    ��?    ����@��@ _� | l��Y{�K����K�A\�-[�^�3��T0 k� ����c�t B%�0d    ��?    ����@��@ _� | l��Y{�K����K�A\�-W�]��3��T0 k� ����c�t B%�0d    ��?    ����@��@ _� � l��Y{�K����K�A\�-S�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ _� � l��Y{�K����K�A\�-O�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ _� � l��Y{�K����K�A\�-G�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ [� � l��Y{�K����K�A\�-C�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ [� � l��Y{�K���K�A\�-?�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ [� � l��Y{�K���K�A\�-;�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ [� � l��Y{�K���K�A\�-7�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ [� � l��Y{�E��K�A\�-3�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ [� � l��Y{�E��K�A\�-/�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ W� � l��Y{�E��K�A\�-+�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ W� � l��Y{�E��K�A\�-'�m��3��T0 k� ����c�t B%�0d    ��?    ����@��@ W� � l��Y{�E��K�A\�-#�=��3��T0 k� ����c�t B%�0d    ��?    ����@��@ W� � l��Y{�E���K�A\�-�=��3��T0 k� ����c�t B%�0d    ��?    ����@��@ W� � l��Y{�E���K�L�-�=��3��T0 k� ����c�t B%�0d    ��?    ����@��@ S� � l��Y{�E���K�L�-�=��3��T0 k� ����c�t B%�0d    ��?    ����@��@ S� � l��Y{�E���K�L�-�=��3��T0 k� ����c�t B%�0d    ��?    ����@��@ S� � l��Y{�E���K�L�-�=��3��T0 k� ��� c�t B%�0d    ��?    ����@��@ S� � l��Y{�E���K�L�-�=��3��T0 k� � �c�t B%�0d    ��?    ����@��@ S� �
 l��Y{�E}#��K�L�-�=��3��T0 k� ��c�t B%�0d    ��?    ����@��@ S� �
 l��Y{�E}'��K�L�-��s�3��T0 k� ��c�t B%�0d    ��?    ����@��@ O� �
 l��Y{�E}+��K�L���o�3��T0 k� ��c�t B%�0d    ��?    ����@��@ O� �
 l��Y{�E}/��K�L���g�3��T0 k� ��c�t B%�0d    ��?    ����@��@ O� �
 l��Y{�E}/�|K�L���_�3��T0 k� ��c�t B%�0d    ��?    ����@��@ O� �
 l��Y{�E}3�|K�L���[�3��T0 k� ��c�t B%�0d    ��?    ����@��@ O� �	 l��Y{�E}7�|K�L���S�3��T0 k� ��c�t B%�0d    ��?    ����@��@ O� �	 l��Y{�Em7�|K�L���K�3��T0 k� �� c�t B%�0d    ��?    ����@��@ O� �	 l��Y{�Em;�|K�L,����G�3��T0 k� � �$c�t B%�0d    ��?    ����@��@ K� �	 l��Y{�Em?�|K�L,����?�3��T0 k� �$�(c�t B%�0d    ��?   ����@��@ K� �	 l��Y{�Em?��K�L,����?�3��T0 k� �$�(c�t B%�0d    ��?    ����@��@ K� �	 l��Y{�EmC��K�L,�����;�3��T0 k� �(�,c�t B%�0d    ��?    ����@��@ K� �	 l��Y{�D=C��K�L,�����7�3��T0 k� �,�0c�t B%�0d    ��?    ����@��@ K� �	 l��Y{�D=C��O�L,�����3�3��T0 k� �0�4c�t B%�0d    ��?    ����@��@ K� � l��Y{�D=G��O�L,�����3�3��T0 k� �4�8c�t B%�0d    ��?    ����@��@ K� � l��Y{�D=G��O�L,����/�3��T0 k� �4�8c�t B%�0d    ��?    ����@��@ K� � l��Y{�D=G��O�L,����+�3��T0 k� �8�<c�t B%�0d    ��?    ����@��@ K� � l��Y{�D=G��O�L,����'�3��T0 k� �<�@c�t B%�0d    ��?    ����@��@ K� � l��Y{�D=G��S�L,����#�3��T0 k� �@�Dc�t B%�0d    ��?    ����@��@ K� � l��Y{�D=G��S�L,��߸��3��T0 k� �D�Hc�t B%�0d    ��?    ����@��@ K� � l��Y{�DMK��S�L,��۸]�3��T0 k� �D�Hc�t B%�0d    ��?    ����@��@ K� � l��Y{�DMK��W�L,��ӷ]�3��T0 k� �H�Lc�t B%�0d    ��?    ����@��@ K� � l��Y{�DMK��W�L,��϶]�3��T0 k� �L�Pc�t B%�0d    ��?    ����@��@ K� � l��Y{�DMG��[�L,��ǵ]�3��T0 k� �P�Tc�t B%�0d    ��?    ����@��@ K� � l��Y{�DMG��[�L,��ô]�3��T0 k� �P�Tc�t B%�0d    ��?    ����@��@ K� � l��Y{�EmG��_�L,����]�3��T0 k� �T�Xc�t B%�0d    ��?    ����@��@ K� � l��Y{�EmG��_�L,����]�3��T0 k� �X�\c�t B%�0d    ��?    ����@��@ K� � l��Y{�EmG��c�L,����]�3��T0 k� �\�`c�t B%�0d    ��?    ����@��@ K� � l��Y{�EmG��c�L,����]�3��T0 k� �`�dc�t B%�0d    ��?    ����@��@ K� � l��Y{�EmC��g�L,����\��3��T0 k� �`�dc�t B%�0d    ��?    ����@��@ K� � l��Y{�E]C��k�L,����\��3��T0 k� �d�hc�t B%�0d    ��?    ����@��@ K� � l��Y{�E]C��k�L,����\��3��T0 k� �h�lc�t B%�0d    ��?    ����@��@ K� � l��Y{�E]?��k�L,����\��3��T0 k� �l�pc�t B%�0d    ��?    ����@��@ K� � l��Y{�E]?��k�L,����\�3��T0 k� �l�pc�t B%�0d    ��?    ����@��@ K� � l��Y{�E];��o�L,���l�3��T0 k� �p�tc�t B%�0d    ��?    ����@��@ O� � l��Y{�C�7��o�L,���l�3��T0 k� �t�xc�t B%�0d    ��?    ����@��@ O� � l��Y{�C�7��o�L,���l�3��T0 k� �x�|c�t B%�0d    ��?    ����@��@ O� � l��Y{�C�3��o�L,���l�3��T0 k� �x�|c�t B%�0d    ��?    ����@��@ O� � l��Y{�C�/��o�L,���l�3��T0 k� �|��c�t B%�0d    ��?    ����@��@ O� � l��Y{�C�/��o�L,���l�3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E]+��s�L,��l�3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E]'��s�L,�{�lߥ3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E]#��s�L,�{�lߤ3��T0 k� ����c�t B%�0d    ��?   ����@��@ O� � l��Y{�E]��w�L,�w�lۣ3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E]�w�L,��s�lۢ3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EM�{�L,��s�lס3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EM�{�L,��s�lנ3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EM�{�L,��o�lӟ3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EM�{�L,��o�lϟ3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EM��L��o�lϞ3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EM��L��o�l˝3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EL����L��o�l˜3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E<����L��o�lǛ3��T0 k� ����c�t B%�0d    ��?   ����@��@ O� � l��Y{�E<����L��o�lǛ3��T0 k� ����c�t B%�0d    ��?   ����@��@ O� � l��Y{�E<���L��o�lÚ3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E<�܏�A\��o�lÙ3��T0 k� ����c�t B%�0d    ��?   ����@��@ O� � l��Y{�E<�܏�A\��o�l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E<�ܓ�A\��o�l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E<�ܓ�A\��s�l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E<߱ܗ�A\��s�l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E,۱ܗ�A\��s�l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E,ױܛ�A\��w�l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E,ӱܟ�A\��w�l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E,ϱܣ�A\��w�l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E,ϰܧ�A\��{�l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E,ϰܧ�A\��{�l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�E,ϯܫ�A\���l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EϮ쫼A\����l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eϭ쯻A\����l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EϬ쯻A\����l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eϫ쳺A\����l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EϪ췹A\����l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eϩ췹A\����l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EϨ컸A\����l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eϧ컷A\���l��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eϧ쿷A\���\��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EϦ쿶A\���\��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eϥ�öA\���\��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eϥ�õA\���\��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EϤ�ǵA\���\��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�EϤ�ǵA\���\��3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eϣ�ǴA\������3��T0 k� ����c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eϣ�ǴA\������3��T0 k� ��� c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eϣ�˴A\������3��T0 k� � �c�t B%�0d    ��?    ����@��@ O� � l��Y{�EϢ�˴A\������3��T0 k� � �c�t B%�0d    ��?    ����@��@ O� � l��Y{�EϢ�˴A\������3��T0 k� ��c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eӡ�˳A\������3��T0 k� ��c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eӡ�˳A\������3��T0 k� ��c�t B%�0d    ��?    ����@��@ O� � l��Y{�Eӡ�˳A\������3��T0 k� ��c�t B%�0d    ��?    ����@�@ O� � l��Y{�E�ӡ˳A\������3��T0 k� ��c�t B%�0d    ��?    ����@�@ O� � l��Y{�E�נ˳A\������3��T0 k� ��c�t B%�0d    ��?    ����@�@ O� � l��Y{�E�נ˳A\���L��3��T0 k� ��c�t B%�0d    ��?    ����@�@ O� � l��Y{�E�۠˳A\���L��3��T0 k� ��c�t B%�0d    ��?    ����@�@ O� � l��Y{�E�۠˳A\���L��3��T0 k� �� c�t B%�0d    ��?    ����@�@ O� � l��a��D�۠L˳A\���L��3��T0 k� �� c�t B%�0d    ��?    ����@��@ b��s�=��Y|/�C�'�r�kE����.S?����T0 k� �����c�t B%�0d   ��;   ��� ��@ b��s�>	��Y|/�C�#�b�jEq���.S;����T0 k� �����c�t B%�0d    ��;   ��� ��@ b��s�>	��Y|/�C��b�iEq��3�/S7����T0 k� �����c�t B%�0d    ��;   ��� ��@ b��s�>	��Y|/�C��b�iEq��3�/S3����T0 k� �����c�t B%�0d    ��;   ��� ��@ b��s�?	��Y|/�C��b�gEq��3�0S+����T0 k� �����c�t B%�0d    ��;   ��� �#�@ R��c�?	.��a�/�C��b�fEq��3�1C+����T0 k� �����c�t B%�0d    ��+   ��� ��'�@ R��c�?	.��a�/�C��b�fEq���1C+����T0 k� �����c�t B%�0d    ��+   ��� ��+�@ R��c�?	.��a�/�C��b�eEq���2C'�s��T0 k� �����c�t B%�0d    ��+   ��� ��3�@ R��c�?	.��a�/�C���b�cEq���2C#�s��T0 k� �����c�t B%�0d    ��+   ��� ��7�@ ���c�?	��a�/�C���R�bEq���2C#�s��T0 k� �����c�t B%�0d    ��+   ��� ��;�@ ���c�?	��a�/�C���R�aEq���2��s��T0 k� �����c�t B%�0d    ��+   ��� ��;�@ ���c�>	��a�/�C���R�`Eq���2��s��T0 k� �����c�t B%�0d    ��+   ��� ��?�@ ���S�>	��a�/�C���R�_Ea���2��s��T0 k� �����c�t B%�0d    ��+   ��� ��C�@ ���S�>	��a�/�C���R�_Ea���2��s��T0 k� �����c�t B%�0d    ��+   ��� ��C�@ ���S�>	.��a�/�C���R�^Ea���2��s��T0 k� �����c�t B%�0d    ��+   ��� ��G�@ ��S�=	.��Y|/�C���R�\Ea����1��s��T0 k� �����c�t B%�0d    ��+   ��� ��G�@ ����=	.��Y|/�C���R�[Eb���1���s��T0 k� �����c�t B%�0d    ��+   ��� ��K�@ ����=	.��Y|/�C���R�[Eb���1������T0 k� �����c�t B%�0d    ��+   ��� ��K�@ ����=	��Y|/�C����ZD2���0������T0 k� �����c�t B%�0d    ��+   ��� ��K�@ ����=	��Y|/�C����YD2���0������T0 k� �����c�t B%�0d    ��+   ��� ��K�@ ����=	��Y|/�C����XD2 ��/������T0 k� �����c�t B%�0d    �+   ��� ��K�@ �{���<	þY|/�C����WD2��.���s��T0 k� �l �p c�t B%�0d    ��/   ��� ��K�@ �s���<	.þY|/�C����VEb��-���s��T0 k� �`�dc�t B%�0d    ��/   ��� ��K�@ �g���<	.þY|/�C����UEb��-���s��T0 k� �T�Xc�t B%�0d    ��/   ��� ��K�@ R_���<	.þY|/�C����TEb��,���s��T0 k� �H�Lc�t B%�0d   ��/   ��� ��K�@ RW���<	.þY|/�C����TEb��+���s��T0 k� �<�@c�t B%�0d   ��/   ��� ��G�@ RK���;	.þY|/�C����SEb
��*���s��T0 k� �,	�0	c�t B%�0d   ��/   ��� ��G�@ RC���;	þY|/�C����REb��)���s��T0 k� � �$c�t B%�0d   ��/   ��� ��G�@ R;���;	þY|/�C�{��QEb��(������T0 k� ��c�t B%�0d   ��/   ��� ��C�@ R/���;	þY|/�C�w��PEb��'¿����T0 k� ��c�t B%�0d   ��/   ��� ��?�@ B���;	þY|/�E�g��NEb��%·����T0 k� ����c�t B%�0d   ��/   ��� ��?�@ B���;�þY|/�E�_��MER��$³����T0 k� ����c�t B%�0d   ��/   ��� ��;�@ B���;�ǾY|/�E�[��LER��#¯����T0 k� ����c�t B%�0d    ��/   ��� ��;�@ B���:�ǾY|/�E�S��JER��!«����T0 k� ����c�t B%�0d    ��/   ��� ��7�@ A���:�ǾY|/�E�K��IER�� «����T0 k� ���c�t B%�0d    ��/   ��� ��7�@ A���:�ǾY|/�E�C��HER��B�����T0 k� ���c�t B%�0d    ��/   ��� |�3�@ A���:�˾Y|/�E�;�b�GER��B��s��T0 k� ���c�t B%�0d    ��/   ��� w�+�@ A���:�˾Y|/�E�/�b|EER��B��s��T0 k� �!��!c�t B%�0d    /�/   ��� r�+�@ A���:�ϾY|/�C�'�bxCER��B��s��T0 k� �x#�|#c�t B%�0d    ��/   ��� m�'�@ A���:�ϾY|/�C��btBER ��2��s��T0 k� �l%�p%c�t B%�0d    ��/   ��� h�#�@ A���9�ӾY|/�C��bpAC�!��2��s��T0 k� �`'�d'c�t B%�0d    ��/   ��� g4�@ 1���9�ӾY|/�C��bl@C�"��2��s��T0 k� �L*�P*c�t B%�0d    ��'   ��� f4�@ 1���9�׾Y|/�C��bh>C�#��2��s��T0 k� �D)�H)c�t B%�0d    ��'   ��� e4�@ 1���9�ۿY|/�C���R`<C�&��2��s��T0 k� �<.�@.c�t B%�0d    ��'   ��� c4�@ 1���9�߿Y|/�C��R\:C�'��2�s��T0 k� �82�<2c�t B%�0d    ��'   ��� a4�@ 1��9�߿Y|/�C��RX9C�(��2{�s��T0 k� �44�84c�t B%�0d    ��'   ��� _4�@ 1s��9���Y|/�C��RT8C�*	Ӏ2{�s��T0 k� �06�46c�t B%�0d    ��'   ��� ]4�@ 1k�x9���Y|/�C�۲RL7C�+	Ӏ2w�s��T0 k� �,7�07c�t B%�0d    ��'   ��� [3��@ 1c�t8���Y|/�C�ӱRH5C� ,	�|
2s�s��T0 k� �$7�(7c�t B%�0d    ��'   ��� Y3��@ A[�l8���Y|/�C�˱RD4C��-	�|
2s�s��T0 k� � 7�$7c�t B%�0d    ��'   �   W3��@ AS�d8���Y|/�C�ðR<3C��.	�|	2o�s��T0 k� �7� 7c�t B%�0d    ��'   �  U3��@ AK�\8���Y|/�C�R82C��/	�|	2o�3��T0 k� �7�7c�t B%�0d    ��'   �  SC��@ A;�P8���Y|/�C�R82C��1	�|2k�3��T0 k� �6�6c�t B%�0d    ��'   �  RC��@ A3�H8���Y|/�C�R41C��2	�|2k�3��T0 k� �6�6c�t B%�0d    ��'   �  QC��@ A+��@8���Y|/�C�R01C��3	�|2g�3��T0 k� �6�6c�t B%�0d    ��'   �  OC��@ A#��88���Y|/�C�R(0EQ�4	�|2g�3��T0 k� �6�6c�t B%�0d    ��'   �  MC��@ A��08��Y|/�C���R$/EQ�5	�|2g�3��T0 k� � 5�5c�t B%�0d    ��'   �  Kc��@ A��(8��Y|/�C���B /EQ�6	�|2g�3��T0 k� ��8� 8c�t B%�0d    ��'   �  Ic��@ A�� 7��Y|/�C��B.EQ�7	�|2c�3��T0 k� ��9��9c�t B%�0d    ��'   �  Gc��@ A��7��Y|/�D w�B.EQ�8	�|2c�3��T0 k� ��:��:c�t B%�0d    ��'   �  Ec��@ P���7��Y|/�D o�B-EQ�9	�|"c�3��T0 k� ��:��:c�t B%�0d    ��'   �  Cc��@ P���7��Y|/�D g�B-EQ�:	�|"c�3��T0 k� ��;��;c�t B%�0d    ��'   �  AS��@ P����7��Y|/�D _��-EQ�;	�|"_�3��T0 k� ��6��6c�t B%�0d    ��'   �  ?S��@ P����7��Y|/�D W�� ,EA�<	�|"_�3��T0 k� ��3��3c�t B%�0d    ��'   �  =S��@ P����7��Y|/�D K���+EA�>�|"_�3��T0 k� ��/��/c�t B%�0d    ��'   �  ;S��@ P����7��Y|/�D C���+EA�>�|�_�3��T0 k� ��-��-c�t B%�0d    ��'   �  9㗺@ 0����7��Y|/�D ;���*EA�?�|�_�3��T0 k� ��+��+c�t B%�0d    ��'   �  7㏸@ 0����7��Y|/�D 3�a�*Eь@�|�_�3��T0 k� �+��+c�t B%�0d    ��'   �  5ㇷ@ 0����7��Y|/�D +�a�)EфA�|�_�3��T0 k� �*��*c�t B%�0d    ��'   �  3��@ 0���6��Y|/�D#�a�)EрA�|�c�3��T0 k� �*��*c�t B%�0d    ��'   �  1�{�@ 0���6��Y|/�D�a�)E�xB�|�c�3��T0 k� �)��)c�t B%�0d    ��'   �  /�s�@ 0���6��Y|/�D�a�(E�pC�|�c�3��T0 k� �|)��)c�t B%�0d    ��'   �  -�k�@ 0���6��Y|/�D�Ѽ(E�hD�|�c�3��T0 k� �|(��(c�t B%�0d    ��'   �  +�c�@ 0���6��Y|/�D�Ѵ'E�`D�|�g�3��T0 k� �|&��&c�t B%�0d    ��'   �  )�[�@ 0���6��Y|/�D��Ѭ'E�XE�|�g�3��T0 k� �x%�|%c�t B%�0d    ��'   �  &�S�@  ���6��Y|/�D�Ѥ'E�TF�|�g�3��T0 k� �t$�x$c�t B%�0d    ��'   �  #�K�@  ��|6��Y|/�D�ќ&EQLF�|�h 3��T0 k� �p$�t$c�t B%�0d    ��'   �   �G�@  ��t6��Y|/�D�є&EQDG�|h3��T0 k� �l$�p$c�t B%�0d    ��'   �  �?�@  ��l6��Y|/�D۞�%EQ<HS|l3��T0 k� �h�lc�t B%�0d    ��'   �  �7�@  ��d6��Y|/�DӞ�%EQ4HS|l3��T0 k� �`�dc�t B%�0d    ��'   �  �'�@  �P6��Y|/�C�Ý�t$EQ$JS|p3��T0 k� �P�Tc�t B%�0d    ��'   �  ��@  {�H6O�Y|/�Cﻜ�l$EQJS|t3��T0 k� �H�Lc�t B%�0d    ��'   �  ��@  w�@6O�Y|/�Cﳜ�d#EQKS|x3��T0 k� �@�Dc�t B%�0d    ��'   �  ��@  p 86O�Y|/�C﫜�\"EQKS|x	3��T0 k� �8�<c�t B%�0d    ��'   �  ��@  l06O�Y|/�C�T"EQLS||3��T0 k� �0�4c�t B%�0d    ��'   �  ���@ l(5O�Y|/�I����L!EP�MS|�3� T0 k� �(�,c�t B%�0d    ��'   �  	���@ h5O�Y|/�I����D E@�MS|�3� T0 k� � 
�$
c�t B%�0d    ��'   �  �@ h5O�Y|/�I����< E@�NS|�3� T0 k� ��c�t B%�0d    ��'   �  �@ d
5O�Y|/�I����4E@�NS|�3� T0 k� ��c�t B%�0d    ��'   �  ߠ@ d5O�Y|/�I����,E@�OS|�3� T0 k� � �c�t B%�0d    ��'   �  נ@ d�5O�Y|/�I���$E@�OS|�3�T0 k� ����c�t B%�0d    ��'   � ��ϟ@ `�5���Y|/�I�w��E@�OS|�3�T0 k� ����c�t B%�0d    ��'   � ��Ǟ@ `�5���Y|/�I�s��E@�OS|�3�T0 k� ����c�t B%�0d    ��'   � ����@ `�5���Y|/�I�o��E@�PS|�3�T0 k� ����c�t B%�0d    ��'   � ����@ `�5���Y|/�I�g��E@�PS|�3�T0 k� ����c�t B%�0d    ��'   � ����@ `�5���Y|/�I�c���E@�PS|�3�T0 k� ��
��
c�t B%�0d    ��'   � ����@ �`�5���Y|/�I�_���E@�PS|�3�T0 k� ����c�t B%�0d    �'   � ����@ �`��5���Y|/�I�[� �E0�PS|�3�T0 k� ���c�t B%�0d    ��/   � ����@ �`�5���Y|/�I�W� �E0�PS|"�3�T0 k� ���c�t B%�0d   ��/   � ����@ �d�5���Y|/�I�S� �E0�PS|"� 3�T0 k� ���c�t B%�0d   ��/   � ����@ �d�5���Y|/�I�O� �E0�PS|"�"3�T0 k� � �� c�t B%�0d   ��/   � ���@ �d �5���Y|/�I�K� �E0|PS|"�#3�T0 k� ������c�t B%�0d   ��/   � ��w�@ �h!�5���Y|/�I�G� �E0tPS|"�%3�T0 k� �����c�t B%�0d   ��/   � ��o�@ �h"�5���Y|/�I�C�0�E0lPS|2�&3�T0 k� �o��s�c�t B%�0d   ��/   � ��c�@ �h#�5���Y|/�I�?�0�E0dOS|2�'3�T0 k� �c��g�c�t B%�0d   ��/   � ��[�@ �l$�|5���Y|/�I�;�0�C@`OS|2�)3�T0 k� �W��[�c�t B%�0d   ��O   � ��S�@ �l%�p5���Y|/�I�7�0�C@XOS|2�*3�T0 k� �K��O�c�t B%�0d   ��O   � ��K�@ �p&�h5���Y|/�I�3�0�C@PNS|2�+3�T0 k� �?��C�c�t B%�0d   ��O   � ��C�@ �t'�`4���Y|/�I�/�@�C@LNS|2�,3�T0 k� �3��7�c�t B%�0d   ��O   � ���;�@ �t(�X4���Y|/�I�+�@�C@DMS|2�-3�T0 k� �'��+�c�t B%�0d   ��O   � ���3�@ �x(�P4޿�Y|/�I�'�@�C@<MS|2�-3� T0 k� ����c�t B%�0d   ��O   � ���+�@ px)�H4޻�Y|/�I�#�@�C@8LS|2�.3� T0 k� ����c�t B%�0d   ��O   � ���#�@ p|*�@4޷�Y|/�I��@�C@0LS|B�/3� T0 k� ����c�t B%�0d   ��O   � ����@ p�*�44���Y|/�I��@�C@,KS|B�03� T0 k� ������c�t B%�0d   ��O   � ��R�@ p�+�,4���Y|/�I��@xC@$JS|B�03��T0 k� ������c�t B%�0d   ��O   � ��R�@ p�+�$4�� Y|/�I��@tC@IS|B�13��T0 k� ������c�t B%�0d   ��O   � ��Q��@ p�+�4��Y|/�I��@pC@IS|B�23��T0 k� ������c�t B%�0d   ��O   � ��Q��@ `�+�4��Y|/�I��@hCPH�|��33��T0 k� ������c�t B%�0d   ��O   � ��Q�@ `�,�4��Y|/�I��@dCPG�|��43��T0 k� ������c�t B%�0d   ��O   � ��Q�@ `�,�4��Y|/�I��@\
CPF�|��53��T0 k� ������c�t B%�0d   ��O   � ��Qߋ@ `�, �4��Y|/�I���@X
CP E�|� 63��T0 k� ������c�t B%�0d   ��O   � ��Q׋@ `�, �4��Y|/�I���@T	C_�D�|� 63��T0 k� ������c�t B%�0d   ��O   � ��Aϊ@ `�, �4��Y|/�I���@L	C_�C3x�73��T0 k� ������c�t B%�0d   ��O   �  ��AÊ@ `�, �4��Y|/�I��@HC_�B3x�83��T0 k� �{���c�t B%�0d   ��O   �����A��@ `�, �4��	Y|/�I��@DC_�A3x�93��T0 k� �o��s�c�t B%�0d   ��O   �����A��@ 0�, �4��
Y|/�C��@@C_�@3x�:3��T0 k� �c��g�c�t B%�0d   ��O   �����A��@ 0�+ �4�|
Y|/�C��@8C_�?3t�;3��T0 k� �W��[�c�t B%�0d   ��O   ����}���@ 0�+ �4�xY|/�C�ߚ@4C_�>3t�<3��T0 k� �K��O�c�t B%�0d   ��O   ����z���@ 0�* �5�xY|/�C�ۚ@0Co�=3p�<3��T0 k� �?��C�c�t B%�0d    ��O   ����w���@ 0�) �5�tY|/�C�ך0,Co�<3p�=3��T0 k� �/��3�c�t B%�0d    ��O   ����s���@ 0�( �6�pY|/�C�Ӛ0(Co�:Cp�>3��T0 k� �#��'�c�t B%�0d    .�O   ����p��@ 0�(�6�lY|/�C�˚0 Co�9Cl�>3��T0 k� ����c�t B%�0d    ��O   ����m�w�@ 0�'�7�hY|/�C�ǚ0Co�8Ch�?3��T0 k� ����c�t B%�0d    ��O   ����j�o�@ 0|&�7�hY|/�C0Co�7Ch�?3��T0 k� �����c�t B%�0d    ��O   ����g�c�@ 0|%�7�dY|/�C0Co�5Cd �@3��T0 k� �����c�t B%�0d    ��O   ����d�[�@ 0x$�8�`Y|/�CPCo�4Cg��@3��T0 k� ����c�t B%�0d    ��O 	  ����a�S�@ 0t#�8�\Y|/�CPCo�2Cc��A3��T0 k� �۳�߳c�t B%�0d    ��O 	  ����^�K�@ @p"�9�XY|/�C���PCo�1C_��A3��T0 k� �ϱ�ӱc�t B%�0d    ��O 	  ����[�C�@ @l!�9�TY|/�C���_� Co�/C[��A3��T0 k� �ï�ǯc�t B%�0d    ��O 	  ����X�;�@ @h x9�PY|/�C���_� C�.C[�c A3��T0 k� ������c�t B%�0d    ��O 	  ����V�/�@ @dt:�LY|/�C���_��C�,CW�c B3��T0 k� ������c�t B%�0d    ��O 	  ����T�'�@ @`l:�HY|/�C���_��C�+SS�c B3��T0 k� ������c�t B%�0d    ��O 	  ����R��@ `\�d;�@Y|/�Eއ�_��C�)SO�b�B3��T0 k� ������c�t B%�0d    ��O 	  ����P��@ `T�\;�<Y|/�E��_��C�(SK�b�B3��T0 k� ������c�t B%�0d    ��O 	  ����N��@ `P�T;�8Y|/�E�w�_��C�&SG�b�B3��T0 k� �s��w�c�t B%�0d    ��F 	  ����L��@ `L�L<�4Y�/�E�o�_��C�$SC�b�B3��T0 k� �c��g�c�t B%�0d    ��F 	  ����J���@ `H�D<�0Y�/�E�g�O��C�#S?�b�B3��T0 k� �W��[�c�t B%�0d    ��F 
  ����H��@ `D�<<�(Y�/�E�c�O��C�!S;�b�B3��T0 k� �K��O�c�t B%�0d    ��F 
  ����G��@ `<�4=�$Y�/�E�[�O��C�S7�b�A3��T0 k� �?��C�c�t B%�0d    ��F 
  ����F��@ `8�(=� Y�/�E�S�O��C�S3�b�A3��T0 k� �;��?�c�t B%�0d    ��F 
  ����E�ۉ@ `4� =�Y�/�E�K�O��CO|S/�b�A3��T0 k� �3��7�c�t B%�0d    ��F 
  ����D�ϊ@ `,�>�Y�/�E�C�߫�COxS+�R�A3��T0 k� �+��/�c�t B%�0d    ��F 
  ����C�Ǌ@ P(�>�Y�/�E�;�ߣ�COxS'�R�A3��T0 k� �#��'�c�t B%�0d    ��F 
  ����B࿊@ P �>�Y�/�E�3�ߛ�COtS#�R�@3��T0 k� ����c�t B%�0d    ��F 
  ����A්@ P� ?�Y�/�E�+�ߓ�COpS�R�@3��T0 k� ����c�t B%�0d    ��F 
  ����@ொ@ P��?> Y�/�E�#�ߋ�E�lS�R�@3��T0 k� ����c�t B%�0d    ��F 
  ����?࣊@ P
��?=�Y�/�E��߃�E�h��R�@3��T0 k� ����c�t B%�0d    ��F 
  ����>���@ P	��?=� Y�/�E���{�E�d����@3��T0 k� ������c�t B%�0d    ��F 
  ����=���@ P��@=� Y�/�E���s�E�`����?3��T0 k� �����c�t B%�0d    ��F 
  ����<���@ _���@=� Y�/�A���k�E�\�����?3��T0 k� ����c�t B%�0d    ��F   ����;���@ _���@=� Y�/�A����c�E�X	�����?3��T0 k� �ӭ�׭c�t B%�0d    ��F   ����:�{�@ _���A=�!Y�/�A���W�E�T�����?3��T0 k� �Ǭ�ˬc�t B%�0d    ��F   ����9�o�@ ����A��!Y�/�A���O�E�P�����?3��T0 k� ����ëc�t B%�0d    ��F   ����8�g�@ ����A��!Y�/�A���G�E�P�����?3��T0 k� ������c�t B%�0d    ��F   ����8�_�@ ����A��!Y�/�A�۟�?�E�L����>3��T0 k� ������c�t B%�0d    ��F   ����8�W�@ �� �B��!Y�/�A�ӟ�7�E�H����>3��T0 k� ������c�t B%�0d    ��F   ����8�O�@ ����B��!Y�/�A�ˠ�/�E�@����>3��T0 k� ������c�t B%�0d    ��F   ����8�C�@ ����B�!Y�/�A�à�#�E�< ����>3��T0 k� ������c�t B%�0d    ��F   ����8�;�@ ���B�!Y�/�E]����E�;�����>3��T0 k� ������c�t B%�0d    ��F   ����8�3�@ ���C�!Y�/�E]����E�7����>3��T0 k� ������c�t B%�0d    ��F   ����8 +�@ ��xC�!Y�/�E]����E�3����=3��T0 k� ������c�t B%�0d    ��F   ����8 #�@ ��pC� Y�/�E]����E�/����=3��T0 k� �����c�t B%�0d    ��F   ����8 �@ ��dC�� Y�/�E]�����E�'����=3��T0 k� �w��{�c�t B%�0d    ��F   ����8 �@ ��\D�� Y�/�E퓤���E�#����=3��T0 k� �o��s�c�t B%�0d    ��F   ����8 �@ ���TD�� Y�/�E틤N��C�����=3��T0 k� �g��k�c�t B%�0d    ��F   ����8��@ ��LD��Y�/�E탥N��C�����|=3��T0 k� �_��c�c�t B%�0d    ��F   ����8��@ �w�DD��Y�/�E�{�N��C�����t=3��T0 k� �[��_�c�t B%�0d    ��F   ����8�@ �k�<D�|Y�/�E�s�N��C�����p<3��T0 k� �S��W�c�t B%�0d    ��F   ����8�@ �c�4E�xY�/�E�o�N��C���w��h<3��T0 k� �K��O�c�t B%�0d    ��F   ����8ۋ@ �[�,E�pY�+�E�g�N��C��o��`<3��T0 k� �C��G�c�t B%�0d    ��F   ����8ˌ@ �G�E�hY�+�A�W�N��C���_�T<3��T0 k� �/��3�c�t B%�0d    ��F   ����8Ì@ �?�E�`Y�+�A�O����C���W�L<3��T0 k� �#��'�c�t B%�0d    ��F   ����8��@ �7�F�\Y�+�A�G����C���O�D<3��T0 k� ����c�t B%�0d    ��F   ����8��@ �/� F�XY�+�A�?����C���G�<<3��T0 k� ����c�t B%�0d    ��F   ����8��@ #��F�PY�+�A�7����C���?�4;3��T0 k� ����c�t B%�0d    ��F   ����8��@ ��F�LY�+�A�/����C���7�,;3��T0 k� ����c�t B%�0d    ��F   ����8��@ ���FHY�+�A�'���C���/�$;3��T0 k� ������c�t B%�0d    ��F   ����8��@ ���GDY�+�A���w�C���'�;3��T0 k� �����c�t B%�0d    ��F   ����8��@ ���G@Y�+�A���k�C����;3��T0 k� ����c�t B%�0d    ��F   ����8{�@ ���G<Y�'�A���c�C����;3��T0 k� ����c�t B%�0d    ��F   ����8s�@ ����G8Y�'�A���[�C����;3��T0 k� �߾��c�t B%�0d    ��F   ����8k�@ ���G�4Y�'�A���S�C�����;3��T0 k� �׿�ۿc�t B%�0d    ��F   ����8�c�@ ���G�0Y�'�A����K�C������:3��T0 k� ������c�t B%�0d    ��F   ����8�[�@ ���G�,Y�'�A���C�C������:3��T0 k� ������c�t B%�0d    ��F   ����8�G�@ ���F�$Y�#�A���/�C������:3��T0 k� ������c�t B%�0d    ��F   ����8�?�@ ��>�F} Y�#�A�߶�'�D����:3��T0 k� ������c�t B%�0d    ��F   ����8O7�@ ��>�F} Y�#�E�׷��Dw����:3��T0 k� ������c�t B%�0d    ��F   ����8O/�@ ��>�F}Y�#�E�ϸ��Do����:3��T0 k� ������c�t B%�0d    ��F   ����8O'�@ ��>xF}Y�#�E�ǹ��Dg����:3��T0 k� ������c�t B%�0d    ��F   ����8O�@ ��>pE}Y�#�E쿺��D_����:3��T0 k� ������c�t B%�0d    ��F   ����8O�@ ^��>dE}Y�#�E컻���DW����:3��T0 k� ������c�t B%�0d    ��F   ����8O�@ ^��>\E}
Y�#�E쳼���DO����:3��T0 k� ������c�t B%�0d    ��F   ����8O�@ ^��>TD�	Y��E������DG����93��T0 k� ������c�t B%�0d    ��F   ����8N��@ ^��>LD�Y��E������D?����93��T0 k� ������c�t B%�0d    ��F   ����8N�@ ^��>DD�Y��E������D7����93��T0 k� ������c�t B%�0d    ��F   ����8��@ ^{�><C�Y��E������D/����x93��T0 k� ������c�t B%�0d    ��F   ����8�ߏ@ ^s�>4C� Y��E������D'����p93��T0 k� ������c�t B%�0d    ��F   ����8�א@ ^g�N,B��Y��E������D����h93��T0 k� ������c�t B%�0d    ��F   ����8�Ǒ@ ^g�NA��Y��E�{����D��o��T93��T0 k� ������c�t B%�0d    ��F   ����8���@ N_�NA��Y��E�w����D��g��L93��T0 k� ������c�t B%�0d    ��F   ����8���@ NS�N@��Y��E�o����D���_��D93��T0 k� �����c�t B%�0d    ��F   ����8���@ NK�N @��Y��E�k����D���W��<93��T0 k� ������c�t B%�0d    �F   ����?���@ NC�M�?��Y��H�c����D���O��093��T0 k� ������c�t B%�0d    ��O   ����F���@ N;�M�?�� Y��H�_�M��D���G��(83��T0 k� ������c�t B%�0d    �O   ����E���@ N3�M�>���Y��H�W�M�D���?�� 83��T0 k� ������c�t B%�0d    ��O   ����D���@ N'�M�>���Y|�H�S�Mw�D���7��83��T0 k� ������c�t B%�0d   ��O   ����C���@ N�M�=���Y|�H�K�Mo�C����/��83��T0 k� ������c�t B%�0d   ��O   ����B�{�@ N�]�<���Y|�H�G�Mg�C����'��83��T0 k� �����c�t B%�0d   ��O   ����A�s�@ N�]�<���Y|#�H�C�M_�C������83��T0 k� �����c�t B%�0d   ��O   ����@�k�@ N�]�;���Y|#�H�;�mW�C������83��T0 k� ܷ����c�t B%�0d   �O    ����@N[�@ N�]�:���Y|#�H�3�mG�EM������83��T0 k� ܯ����c�t B%�0d   �O    ����@NS�@ M����9���Y|#�H�+�m?�EM�� ����83��T0 k� ܫ����c�t B%�0d   ��O    ����@NK�@ M����8���Y|#�H�'�m7�EM�� ����83��T0 k� ܫ����c�t B%�0d   ��O    ����@NC�@ M����8���Y|#�H�#�m3�EM�� ����73��T0 k� ̧����c�t B%�0d   ��O    ����@N;�@ M����7���Y|#�H��]+�EM�� ����73��T0 k� ̣����c�t B%�0d   ��O    ����@N3�@ M����6���Y|#�H��]#�I}{� ���73��T0 k� ̟����c�t B%�0d   ��O    ����@N+�@ M����6���Y|'�H��]�I}o� ���7"s��T0 k� ̛����c�t B%�0d   ��O    ����@#�@ M���x5���Y|'�H��]�I}c� ���6"s��T0 k� ̗����c�t B%�0d   ��O    ����@�@ ���t5���Y|'�H��]�I}[� ����6"s��T0 k� �����c�t B%�0d  	 ��O    ����@�@ ���l4���Y|'�H��M�I}O� ����6"s��T0 k� �����c�t B%�0d  	 ��O    ����@�@ ���d4���Y|'�H��M�C�C� ��0�5"s��T0 k� �����c�t B%�0d  	 ��O    ����@�@ ���\3���Y|'�H��M�C�7� ��0�5"s��T0 k� �����c�t B%�0d  
 ��O    ����@��@ ���X2���Y|'�H��L��C�/���0x5"s��T0 k� �����c�t B%�0d  
 ��O    ����@��@ ���P2���Y|'�H��L��C�#���0p4"s��T0 k� �����c�t B%�0d  
 ��O    ����@�@ ���H1���Y|'�H��<��C����0h4"s��T0 k� ����c�t B%�0d  
 ��O    ����@�@ ���D1���Y|'�H���<��C����0`3"s��T0 k� {���c�t B%�0d   ��O    ����@�@ ���<0���Y|'�H���<��C����0T3"s��T0 k� w��{�c�t B%�0d   ��O    ����@ߢ@ ���80���Y|+�H���<��C����0L23��T0 k� s��w�c�t B%�0d   ��O    ����@ۢ@ ��0/���Y|+�H���<� C���w�0D23��T0 k� �s��w�c�t B%�0d   ��O    ����@ӣ@ w��,/���Y|+�H���L� C���o�0<13��T0 k� �l �p c�t B%�0d   ��O    ����@ϣ@ o��$.���Y|( H���L�C���g�0403��T0 k� �h�lc�t B%�0d   ��O    ����@ǣ@ k�� .���Y|( H���L�C���[�0,03��T0 k� �d�hc�t B%�0d   ��O    ����@ä@ c��-���Y|(H���L�C���S�@$/3��T0 k� �`�dc�t B%�0d   ��O    ����@��@ _��-���Y|(E���L�C����K�@/3��T0 k� �\�`c�t B%�0d   $�O    ����@��@ W��,���a�(E���\�C����C�@.3��T0 k� �`�dc�t B%�0d   ��O    ����@��@ S��,���a�(E���\�C����;�@-3��T0 k� �d�hc�t B%�0d   ��O    ����@��@ O��,���a�(E���\�C����3�@ -3��T0 k� �h�lc�t B%�0d   ��O   ����@��@ G�� +���a�(E���\�C����+�O�,3��T0 k� �l�pc�t B%�0d   ��O    ����@��@ C���+���a�(F��\�C����#�O�+"���T0 k� �p�tc�t B%�0d   ��O    ����@��@ ;���*���a�(F��l�C�����O�*"���T0 k� �t�xc�t B%�0d   ��O    ����@��@ 7���*���a�,F��l�C�����?�*"���T0 k� �t�xc�t B%�0d  
 ��O    ����@��@ 3���)���a�,F��l�C����?�)"���T0 k� �x�|c�t B%�0d  
 ��O    ����@��@ /���)���a�,F��l�I|w���?�("���T0 k� �|��c�t B%�0d  
 ��O    ����@��@ '���)���a�,@��l�I|s����?�'"���T0 k� ����c�t B%�0d  
 ��O    ����@��@ #���(��a�,@��|�I|k����?�'"���T0 k� ����c�t B%�0d  	 ��O    ����@�@ ���(��Y|,@��|�I|c����?�&"���T0 k� ����c�t B%�0d  	 ��O    ����@{�@ ���'��Y|,@��|�I|[����?�%"���T0 k� ����c�t B%�0d  	 ��O    ����@w�@ ���'��Y|,@��|�E�W����?�%"���T0 k� ����c�t B%�0d   ��O    ����@o�@ ���'��Y|,@k��|�E�O����?�$"���T0 k� ܔ��c�t B%�0d   ��O    ����@k�@ ���&���Y|,@k����	E�C����?�#3��T0 k� ܘ��c�t B%�0d   ��O    ����@g�@ ���&���Y|,@k����	E�3����?�#3��T0 k� ܜ��c�t B%�0d   ��O    ����@c�@ ���&���Y|,@k����	E�'����?�"3��T0 k� ܠ��c�t B%�0d   ��O    ����@_�@ ����%���Y|,	@k����
C�����?�"3��T0 k� ܠ��c�t B%�0d   ��O    ����@[�@ ����%���Y|,	B�����
C�����?�!3��T0 k� ����c�t B%�0d   ��O    ����@W�@ ����%���Y|,	B�����
C�����Ox 3��T0 k� ����c�t B%�0d   ��O    ����@S�@ ����$���Y|,
B����|C�����Op 3��T0 k� ����c�t B%�0d   ��O    ����@O�@ ����$���a�0
B���|C����Ol3��T0 k� ����c�t B%�0d   ��O    ����@K�@ ����$���a�0
B���xC�߬��Od3��T0 k� ����c�t B%�0d   ��?    ����@G�@ ����#���a�0B���tC�ӫ��O`3��T0 k� ���c�t B%�0d   ��?   ����@C�@ ����#���a�0B���tC�ǫ{�OX3��T0 k� ���c�t B%�0d   ��?    ����@?�@ ����#���a�0B���pCۻ�o�OT3��T0 k� ����c�t B%�0d   ��?    ����@;�@ ����#���a�0C��pCۯ�g�OL3��T0 k� ����c�t B%�0d    ��?    ����@7�@ ����#���a�0C��lCۣ�_�OH3��T0 k� ����c�t B%�0d    ��?    ����@7�@ ����#���a�,C��lCۛ�W�O@3��T0 k� ����c�t B%�0d    ,�?    ����@3�@ ����# l��a�,C��lCۛ�O�O<3��T0 k� ����c�t B%�0d    ��?    ����@/�@ ���# l��a�,C��lC۟�G�O43��T0 k� ����c�t B%�0d    ��?   ����@+�@ ���" l��a�(C��hCۣ�?�O03��T0 k� ����c�t B%�0d   ��?    ����@'�@ ���" l��Y|(C#��hCۣ�7�O,3��T0 k� ����c�t B%�0d   ��?    ����@#�@ ���" l��Y|(C'��hCۧ�/�O$3��T0 k� ���c�t B%�0d   ��?    ����@#�@ ���" l��Y|(E,+��dCۧ�'�O 3��T0 k� ���c�t B%�0d   ��?    ����@�@ ���" l��Y|$E,/��dC۫��O3��T0 k� ���c�t B%�0d   ��?    ����@�@ ���|! l��Y|$E,3��dC۫��O3��T0 k� �	��	c�t B%�0d   ��?    ����@�@ ���x! l��Y|$E,7��dCۯ��O3��T0 k� �	��	c�t B%�0d   ��?    ����@�@ ���t  l��Y|$E,;��dCۯ��O3��T0 k� ��	��	c�t B%�0d   ��?    ����@�@ ���t  l��Y| EC��dC۳���O3��T0 k� ��	��	c�t B%�0d   ��?    ����@�@ ���t  l��Y| EG��dA[����O3��T0 k� ��	��	c�t B%�0d   ��?    ����@�@ ���p  l��Y| EK�\dA[����N�3��T0 k� ��	��	c�t B%�0d   ��?    ����@�@ ��p  l��Y| EO�\`A[����N�3��T0 k� ��	� 	c�t B%�0d   ��?    ����@�@ ��l  l��Y|ES�\`A[�����N�3��T0 k� � 
�
c�t B%�0d   ��?    ����@�@ ��l l��Y|B�[�\`A[�����N�3��T0 k� �
�
c�t B%�0d   ��?    ����@��@ ��h l��Y|B�_�\`A[�����N�3��T0 k� �
�
c�t B%�0d   ��?    ����@��@ ��h l��Y|B�c��\A[�����N�3��T0 k� �
�
c�t B%�0d   ��?    ����@��@ ��h l��Y|B�k��\A[î��N�3��T0 k� �
�
c�t B%�0d   ��?    ����@��@ ��h l��Y|B�o��\A[î��N�3��T0 k� �
�
c�t B%�0d   ��?    ����@��@ ���d l��Y|K�s��XA[Ǯ��N�3��T0 k� �
�
c�t B%�0d   ��?    ����@�@ ���d l��Y|K�{��XA[Ǯ��N�3��T0 k� ��c�t B%�0d   ��?    ����@�@ ���d l��Y|K���TA[˯��N�3��T0 k� �� c�t B%�0d   ��?    ����@�@ ���d l��Y|K����TA[˯��N�3��T0 k� � �$c�t B%�0d   ��?    ����@�@ ���d l��Y|K����P
A[ϯ��N�3��T0 k� �$�(c�t B%�0d   ��?    ����@�@ ���d l��Y|K����P	A[ϯ��N�3��T0 k� �(�,c�t B%�0d   ��?    ����@�@ ���h l��Y|K����P	A[ϰ�{�N�3��T0 k� �,�0c�t B%�0d    ��?    ����@�@ ���h l��Y|K����LA[Ӱ�s�N�3��T0 k� �0�4c�t B%�0d    ��?    ����@�@ ���h l��Y|K����LA[Ӱ�k�N�3��T0 k� �4�8c�t B%�0d    ��?    ����@�@ ���h l��Y|K���HA[װ�c�N�3��T0 k� 8�<c�t B%�0d    /�?    ����@߶@ �� h l��Y|K���HA[װ�[�N�3��T0 k� 8�<c�t B%�0d    ��?    ����@߶@ �� h l��Y|K���HA[ױ�S�>�3��T0 k� <�@c�t B%�0d    ��?    ����@߶@ �� l l��Y|K���DA[۱�K�>�3��T0 k� @�Dc�t B%�0d    ��?    ����@߷@ �� l l��Y|K���DA[۱�C�>�3��T0 k� D�Hc�t B%�0d    ��?    ����@߷@ �� l l��Y|K����DA[߱�;�>�3��T0 k� H�Lc�t B%�0d    ��?   ����@߷@ �� l l��Y|K����D A[߱�3�>�3��T0 k� L�Pc�t B%�0d    ��?    ����@߸@ �� l l��Y|K����G�A[߲�+�>�3��T0 k� P�Tc�t B%�0d    ��?    ����@߸@ �� l l��Y|K����G�A[�#�>�3��T0 k� T�Xc�t B%�0d    ��?    ����@߸@ �� p l��Y|K����G�A[��>�3��T0 k� X�\c�t B%�0d    ��?    ����@߹@ �� p l��Y|K���|G�A[��>�3��T0 k� �X�\c�t B%�0d    ��?    ����@߹@ � p l��Y|K���|G�A[��>�3��T0 k� �\�`c�t B%�0d    ��?    ����@߹@ � p l��Y|K�æ|G�A[��>�3��T0 k� �`�dc�t B%�0d    ��?    ����@߹@ � p l��Y|K�å|G�A[���>�3��T0 k� �d�hc�t B%�0d    ��?    ����@ߺ@ {� p l��Y|K�ǥ|G�A[���>�
3��T0 k� �h�lc�t B%�0d    ��?    ����@ߺ@ {� p l��Y|K�Ǥ|G�A[���>�
3��T0 k� �l�pc�t B%�0d    ��?    ����@ߺ@ {� t l��Y|K�ˣ|G�A[���>�	3��T0 k� �p�tc�t B%�0d    ��?    ����@ߺ@ w� t l��Y|K�ϣ|G�A[���>|	3��T0 k� �t�xc�t B%�0d    ��?    ����@߻@ w� t l��Y|K�Ϣ|G�A[���>x3��T0 k� �x�|c�t B%�0d    ��?    ����@߻@ w� t l��Y|K�ӡ|G�A[���>t3��T0 k� �x�|c�t B%�0d    ��?    ����@߻@ s� t l��Y|K�ӡ|G�A[���Np3��T0 k� �|��c�t B%�0d    ��?    ����@߻@ s� t l��Y|K�נ|G�A[���Nh3��T0 k� ����c�t B%�0d    ��?    ����@߼@ s� t l��Y|K�ן|G�A[�-��Nd3��T0 k� ����c�t B%�0d    ��?    ����@߼@ s� t l��Y|K�۟|G�A[�-��N`3��T0 k� ����c�t B%�0d    ��?    ����@߼@ o� x l��Y|K�۞�G�A[��-��N\3��T0 k� ����c�t B%�0d    ��?    ����@߼@ o� x l��Y|K�ߞ�G�A[��-��NX3��T0 k� ����c�t B%�0d    ��?    ����@߽@ o� x l��Y|K�ߝ�G�A[��-��NP3��T0 k� ����c�t B%�0d    ��?    ����@߽@ o� x l��Y| K���G�A[��-��NL3��T0 k� ����c�t B%�0d    ��?    ����@߽@ k� x l��Y| K���K�A[��-��NH 3��T0 k� ����c�t B%�0d    ��?    ����@߽@ k� x l��Y| K���K�A[��-��NC�3��T0 k� ����c�t B%�0d    ��?    ����@߾@ k� x l��Y| K���K�A[��-��N?�3��T0 k� ����c�t B%�0d    ��?    ����@                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��/ ]�(((' � ���g          ��A��    �� {�AH=    �,             
   ��         ��     ���   
0	          �n       �  (�    �n  (�               ��      	 ����        �0       ���   (
          ���L          �hc    �����hR    �C                 �         $`     ���   8�

          ��           �%��     ��%�z    �� ]              
   �$           �     ���   (	          ��;
          .�%�    ��;
�%�                   
    �$          #�     ���   P
B           5� 
     B��;�     /���>?     `��                      ��              	  ���  8		 1             ��4� M X
     V�6��    ��H;�6u�    �s�             ���@         "p�   
  ��@ @0	%          ��ݔ  $ P     j�2i�    ��ݔ�2i�                     # 	���@          #p     ��@ 0
 
         ���K   
	   ~��    ���x�"2    ����          	���@         ��  �  ��H   8
          ���s  1 1     ��+W�    ��� �*�i     ��                ���@         	 ��     ��@   8         ���  $ $    ��.$�    �����-�     �&              X���@         
   �     ��@ P	         ��Q� ��     � �b�    ��Q� �b�                             ���|            (  ��@    P                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          ��  ��        ����     ���)Q    p
G "                x                j  �   �   �                              ��       ���         ��           "                                                �                         �A  ��%�%���6�2��+�. ������� 
      	          
     �e �R�G       �d �h@ ��  i@ �d i� AD �j� BD  k� B� l ���J ����X ����J ����X ����X ����  ����. ����< ����J ����X � �  s@ 
� V� 
�< V� 
�\ W  
�< W� 
�� W� 
�\ W� � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� �R� 
�< U� 
�� V  
�| V ���� ����� ����� � 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����@������ �  ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"     �j @�    �
� �  �  
� ��    ��     ��  �    ��  ��     ��%      ��    ��     ��          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �?%      �� � �  ���        �
 �  ���        �        ��        �        ��        �    ��     I� !��        ��                         ��  0 � ���                                     �                ���              �
���%��  ���@�� F�2            �HFD y Yake gilny    0:00                                                                        7  7     �"�""�9KBPKJH KL`k~ �8 k� �C �	C � �
C6 �C.C6* �c� � c� � c� � �c� � � c� � �cj � � cp � � cq � �kV � �k^ � � k` � �B� � �B� b �T a �S"�- "�?"�-*�<8 "� �8 !"� �("� �(#
� � x$"* z �%"2 z � &"@ z �'": � � ("P � �)!� � *"* z+"< � ,"2 z8-"6 z8."
 �@ /"L �X 0"R �`  "K �`  "K �`  "K �`  "K �@ 5"D �` 6"K �`  "K �`  "K �` 9"G �`  "K � �;*4F �  *Nf �=!� �>!� � ".                                                                                                                                                                                                                         �� P `       �     @         �     W P E f  ��                    	�������������������������������������� ���������	�
��������                                                                                          ��    ��`�� ��������������������������������������������������������   �4, J  < Q�� b
 ��� ł��@����@��A������H���_�                                                                                                                                                                                                                                                                                                              4"@r ��"                                                                                                                                                                                                                                            �       
     �  L�J      ��                             ������������������������������������������������������                                                                                                                                     g   ��           �  ;          ��                 	 	 ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ���                                    0         D�J    	  �U                             ������������������������������������������������������                                                                                                                                      {     �      �        �        �  �          	  
 	 
 	 	 ���������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������           �                                                                                                                                                                                                                                       
                                                                       �             


             �  }�         ������������      $��������������������  *�����    ��������������������     'p������������������������                                           R�                    y�               ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" A C 6                	                 � E&
U �\        �t�S$
�C$+TA                                                                                                                                                                                                                                                              )n)nE  1n                                a      m                                                                                                                                                                                                                                                                                                                                                                                                                     > �  >�  
�  (�  J�  D7a�  �����q����~�̎���˖�!��� ���p��H�g�����                 | � :�� r	       	  	�   & AG� �   �                 �                                                                                                                                                                                                                                                                                                                                      p I B   �                        !��                                                                                                                                                                                                                            Y��   �� �� �      �� Z  �� ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ������������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������             $ffllf���flll����llll����ll�l����l��������l�l���fl�Ƹ��ˈ�l���ƪ�˻��˪��˫�̼�ff�f�f��ff�lff���flll���˼ff�̼ffffff�ffffffffffff���̶�ff�fff����flflfl��ffll�fl�lʻ�̻��l̻��˻�l�ll����l�l�����ll����̼��������l�l�����lll�����l�l���ʬƬ�fl��flffff��ffl�f�f�f�f��fˉ�f���f��ffl�ffffffff�fffƬ��Ɖ����ffffffffffff�fffff�ffffffflf�fllfff�ffffffffffffffl�fffl��l�����l������ll��f���fll�����fll�f���ffllff�ffflff��klflj����ffff�ffffffl�fk��f���f�Ƽf�̖f��ff�fl�f��fʨ�����ʩ����̚��l����ll�Ɖ�������˙�����̺���ʙ�f����l��f�k���lj���̛lll�˪̪fˬ��̛�kllll���lll�f���f�l�f���lf��f���ll����l��l�����l��������l������l�f���f���j��ɫ��ɘ��i���i���ʈ�����������������������������������������������������ʋ̼Ɖ��l�����������j���j�������̩���ɩ�̺����f�ƺl�l�f��yl�̙f�ƨ��l�f�ƨ���flf�����ff�l����ffllf���flll����f�{�f�z��ʊ��jy��f����x��ƚ��̙�����������������ʪ��˚��̺���˺����˼fff˺�̚�����˪����������������˪��̪�f���l���˻�ƫ̻l�˻jƨf�ƙl�̊f��{l�̛ll̦���flll����flll����llll����lllf���i�fk��l��lɉ��̩��fj�fff���ƪ��ˊ��i������f�˺���ʬl̪��̉��l�����������������˫�l�������˼�ll�fɼlʩ�������f�ˬ�l��l˛�Ʃ�l̚�ff�˻f�ʙ�lll�����ll�l����l�l�����ffflffff$�I    /      D   #�                         4     �  �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �f ��     �f �$ ^$ �@       �       �     �   r 
� �     �f ��        p���� ��   p���� �$ ^h  ��   p   	  ��     �           �� �   6   
���(�� x    �     ����� ��   ����� �$ ^$      
[�   �z �   $   & � ��� �� � ���5O �  �� �       �  ��   ��������2����  g��� 	 �     f ^�         �� C��      �      ��/x���2�������J����  ��      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "" "  """""" "!   " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                              "! "   "      ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  ""   "! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                      �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �                   �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������            �۰ ̽  �̰ ̻� ˸� ��U@��T@UUUJ  ���� �                           �   ��  ���  � �    �                                                                                                                                       ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r` "�"�����   �� �          ����   �       �                                   �    ���  ��                    ��  ��  ���     ��   �  ��  �  �  �         � �������������  �                                                                                                                                                      �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �        �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                   �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �              "      �           �  �   �   ��  �            ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                            � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                                         	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                       ���  +"  "" ���������                   �                        ���� ��� ����            �� ���  ��                                                                                                                                                                                                                         �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �    ���                              �������  �                     �  �   �  �  ��  �  ��  �                                                                                                                    �  �  ��  �                                                                        �� ̽ ̽ ۽�}ک z�� ���
���
��̙�������̽��̘�̙��
� �	�"� �"  .  �
 �  �               �    ���                                    �   ̰  ��  ݚ� ��� ̽� �ͻ ��� �˘ ̸��ˉUP��UZ�UUJETDUDDUU33ET335[3�� ؚ  ��  +   "  �  ��   � �        �   �   @   �   �   �   �   �   �"  ""  !� �� ��  �               �   ������  ��                   �                        ���� ��� ����                            �    � �  ��                  ���                              �   ���                            �   �    ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         �� 
�� ��� ��� ��� ��� ��� ����˭ۻ�؉+��  8�  �E �U �U �T �@  ��  
� ,� "� ""  "   ��  ��� ��� ̸��̺��̸����� ̽� ȉ  ��  4S  UT  DC  C0  33  3  �   ��  �" �"  ""  "�/�����            �  ��� ̻� {�� w}ڠ    �   �� "�" ��" �                                       �   �   ��  � " ��"  "                     �                             ���                         �  ��                    �����                      �  �  �   �   ��  �                            �   ���                            �   �                    �   �� �       �  �  ��  �   �   �   �                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                  � �� ��  ��             �  �˰ ��� �wp ���                                                                                                                                                                             �  �   ��  �   �  �  �  ��  ��  ��  I�  T:  UJ  T   T  T  J  T�  �� 
�� � �  �˰ ��� ��p���p��� ��� ˹� ̻� �̙ ̼� ˼� �ܘ �٪�؋�Ѓ=�Ш3� �C  �0  ��  ;"� "/ �� ��  ��� ,� ""/ """  ���     �      �                           �  ��  �  ��  �              �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ���   �       �                        �   ��  ���  � �    �                                                                                                                                            �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �                   �   �   �   "   "   "  !�    ��                ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                                                                                                                                                                                            �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                     �                        �         �  �� �  �� ��                                                                                                                                                   �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=LL����������D����3333DDDD    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����������A������ x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx""""�������I�I������ w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww""""�������I��D���I�������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(�D�M�D���M������3333DDDD �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""�����AMAD������ M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M""""������������������ � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�fFfFDfFFfFffdFffff3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DDFFDfFFfdFffff3333DDDD 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5""""wwwwwwwGGD x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x""""wwwwwwqwAqwAwA w w x y�������H���������������������������������H������yxww""""wwwwqwqAwAqAqAq  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(A�A�A�A��LD�����3333DDDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,�A�LDL�L�D�L�����3333DDDD +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+""""wwwwwwDGAD 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5""""wwwwqqDAAq =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=""""wwwwwwwGGwGGwGwGw     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( UQUUQUUQUUQUUUDUUUUU3333DDDD � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � �DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq"�""�9KBP" KJ`KKHk~ �8 k� �C �	C � �
C6 �C.C6* �c� � c� � c� � �c� � � c� � �cj � � cp � � cq � �kV � �k^ � � k` � �B� � �B� b �T a �S"�- "�?"�-*�<8 "� �8 !"� �("� �(#
� � x$"* z �%"2 z � &"@ z �'": � � ("P � �)!� � *"* z+"< � ,"2 z8-"6 z8."
 �@ /"L �X 0"R �`  "K �`  "K �`  "K �`  "K �@ 5"D �` 6"K �`  "K �`  "K �` 9"G �`  "K � �;*4F �  *Nf �=!� �>!� � ".3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0����������������������������������������� ��=�K�X�X�_��B�G�Q�K� � � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������2�0�.� ��"�������������������������������������2�0�.�	�
�������������������� � � � � � �����������������������������������������%��������������������,�>�0� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            