GST@�                                                            \     �                                               �   �   �                  � 2�����	 J���������������~���        h     	#    ~���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    
 �j� � 
 ���
��
�"     "�j��   * ��
  ��                                                                              ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             �F  )1          == �����������������������������������������������������������������������������                                �   9       �   @  &   �   �                                                                                 '       )n)n1n  )�1F    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    C��4 oO�q$K������|+�_;�\rAP< @��JA;�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
C��3 oS�a(K������|+�_;�XrAP< @��JA;�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
C��1 oS�a(K������|+�_;�XrAP< @��JA;�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
C��0 oS�a,K����Â|+�_;�TqAP< @��JA?�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
C��. oS�a0K����˂|+�_;�TqAP< @��JA?�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
C��- oS�a4K����ς|+�_;�TqAP< @��JA?�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C��+ oS�14K����ׂ|+�_;�PqAP< @��JA?�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C��* oS�18K����ہ|+�_;�PqAP< @��JAC�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C��( oS�18K�����|+�_;�PqAP< @��JAC�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C��' oS�1<
K�����|+�_;�LqAP< @��JAC�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C��% oS�1<	K�����|+�_;�LpAP< @��JAC�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C��# oS�1@K�����|+�_;�LpAP< @��JAC�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C��" oS�1@K������|+�_;�HpAP< @��JAG�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C��  oS�1@K������|+�_;�HpAP< @��JAG�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C�� oS�A@K�����|+�_;�HpAP< @��JAG�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C�� oS�AD K�����|+�_;�DpAP< @��JAG�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C�� oS�AG�K�����|+�_;�DpAP< @��JAG�3� T0 k� �k��o�e2$  (u1'T   ��   ��� 
C�� oS�AG�K�����|+�_;�DpAP< @��JAK�3� T0 k� �k��o�e2$  (u1'T   ��   ��� 
C�� oW�AG�K�����|+�_;�@oAP< @��JAK�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C�� oW�AG�K�����|+�_7�@oAP< @��JAK�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C�� oW�AG�K����'�|+�_7�@oAP< @��JAK�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C�� oW�AG�K����+�|+�_7�<oAP< @��JAK�3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
C�� oW�1G�K����/�|+�_7�<oAP< @��JAO�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�� oW�1G�K����3�|+�_7�<oAP< @��JAO�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�� oW�1G�K����7�|+�_7�<oAP< @��JAO�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C��
 oW�1G�K����?�|+�_7�8oAP< @��JAO�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�� oW�1G�K����C�|+�_7�8oAP< @��JAO�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�� oW�1G�K����G�|+�_7�8nAP< @��JAO�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�� oW�1C�K����K�|+�_7�8nAP< @��JAS�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�� oW�1C�K����O�|+�_7�4nAP< @��JAS�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�� oW�1C�K����S�|+�_7�4nAP< @��JAS�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C��� oW�1C�K����W�|+�_7�4nAP< @��JAS�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C��� oW�1C�B����[�|+�_7�4nAP< @��JAS�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C��� oW�1C�B����_�|+�_7�0nAP< @��JAS�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C��� oW�1C�B����c�|+�_7�0nAP< @��JAS�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C��� oW�1C�B����g�|+�_7�0nAP< @��JAW�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C��� oW�AC�B����k�|+�_7�0nAP< @��JAW�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C��� oW�AC�B����k�|+�_7�0nAP< @��JAW�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�� oW�AC�B����o�|+�_7�,mAP< @��JAW�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�{� o[�AC�B����o�|+�_7�,mAP< @��JAW�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�{� o[�AC�B����s�|+�_7�,mAP< @��JAW�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�w� o[�AC�E���w�|+�_7�,mAP< @��JAW�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�s� o[�AC�E���w�|+�_7�(mAP< @��JA[�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�o� o[�AC�E���{�|+�_;�(mAP< @��JA[�3� T0 k� �o��s�e2$  (u1'T   ��   ��� 
C�k� o[�AC�E���{�|+�_;�(mAP< @��JA[�3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
C�g� o[�AC�E����|+�_;�(mAP< @��JA[�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
C�g� o[�A?�E����|+�_;�(mAP< @��JA[�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
C�c� o[�A?�E�����|+�_;�(mAP< @��JA[�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
C�c� o[�A?�E�����|+�_?�$mAP< @��JA[�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
C�_� o[�A?�E�����|+�_?�$mAP< @��JA_�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
C�_� o[�A;�E�����|+�_?�$mAP< @��JA_�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
C�_� o[�A7�B������|+�_C�$mAP< @��JA_�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
K�[� o[�A7�B�����|+�_C�$lAP< @��JAc�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
K�W� o[�A3�B�����|+�_C� lAP< @��JAc�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
K�W� o[�A3�B�����|+�_G� lAP< @��JAc�3� T0 k� �s��w�e2$  (u1'T   ��   ��� 
K�S� o[�A/�B�����|+�_G� lAP< @��JAg�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
K�S� o[�A/�B�����|+�_G� lAP< @��JAg�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
K�O� o[�A+�B�����|+�_K� lAP< @��JAg�3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
K�O��[�A+�K�����|+�_K� lAP< @��JAg�3� T0 k� �k��o�e2$  (u1'T   ��   ��� 
K�K��[�A'�K�����|+�_O� lAP< @��JAk�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
K�K��[�A'�K�����|+�_O�lAP< @��JAk�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
K�G��[�A#�K�����|+�_S�lAP< @��JAk�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K�G��[�A#�K���|+�_S�lAP< @��JAo�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
K�C��[�A�K���|+�_S�lAP< @��JAo�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
K�C��[�A�K���|+�_W�lAP< @��JAo�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
K�?��[�A�K���|+�_W�lAP< @��JAo�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
L?��[�A�K���|+�_[�lAP< @��JAs�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
L;��[�A�K�����|+�_[�lAP< @��JAs�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
L;��_�A�K�����|+�_[�lAP< @��JAs�3� T0 k� �[��_�e2$  (u1'T   ��   ��� 
L7��_�A�K�����|+�__�lAP< @��JAs�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
L7��_�A�K�����|+�__�kAP< @��JAw�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
L3��_�A�K�����|+�_c�kAP< @��JAw�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
L3��_�A�K�����|+�_c�kAP< @��JAw�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
L3��_�A�K�����|+�_c�kAP< @��JAw�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
L/��_�A�K�#����|+�_g�kAP< @��JA{�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
L/��_�A�K�#����!�+�_g�kAP< @��JA{�"�� T0 k� �[��_�e2$  (u1'T   ��    ��� 
L+��_�A�K�#��É!�+�_g�kAP< @��JA{�"�� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L+��_�1�K�'��Ê!�+�_k�kAP< @��JA{�"�� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L'��_�1�K�'��Ǌ!�+�_k�kAP< @��JA{�"�� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L'��_�1�K�'��ǋ!�+�_k�kAP< @��JA�"�� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L'��_�1�K�+��ǋ!�+�_o�kAP< @��JA�"�� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L#��_�1�K�+��ǋ!�+�_o�kAP< @��JA�"�� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L#��_�1�K�+��ǌ!�+�_o�kAP< @��JA�"�� T0 k� �_��c�e2$  (u1'T   ��   ��� 
L#��_�0��K�/��ǌ!�+�_s�kAP< @��JA�"�� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�0��K�/��ǌ!�+�_s�kAP< @��JA��"�� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�0��K�/��ǌ!�+�_s�kAP< @ÝJA��"�� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�0��K�3��Ǎ|+�_w�kAP< @ÞJA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�0��K�3��Ǎ|+�_w�kAP< @ÞJA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�0��K�3��ǎ|+�_w�kAP< @ßJA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�`��K�7��ǎ|+�_{�kAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�`��K�7��Ǐ|+�_{�kAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�`��K�7��Ǐ|+�_{�kAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�`��K�;��Ï|+�_�kAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�`��K�;��Ï|+�_�kAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�`��K�;��Ï|+�_�kAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�P��K�;�࿐|+�_�kAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�P��K�?��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�P��K�?��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�P�K�?��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_�P�K�?��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_���K�C��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_���K�C�@��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_���K�C�@��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_���K�C�@��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_���K�G�@��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
L��_���K�G�@��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K���_��K�G�@��!�+�_��jAP< @��JA��"s� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K���_��K�G�@��|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K���c�ߠK�K�@��|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K���c�ߠK�K�@��|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K���c�۟K�K����|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K���c�۟K�K����|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K���c�מK�K����|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K���c�מK�O����|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K����c�מK�O����|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K����c�ӝK�O����|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K����c�ӝK�O����|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K����c�ϜK�O����|+�_��jAP< @��JA��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
K��� oc�ϜB�O���|+�_��jAP< @��JA��3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
K��� oc�˜B�O��{�|+�_��jAP< @��JA��3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
K��� oc� ˛B�O��w�|+�_��jAP< @��JA��3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
K��� oc� ˛B�S��s�|+�_��jAP< @��JA��3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
K��� oc� ǛB�S��k�|+�_��jAP< @��JA��3� T0 k� �w��{�e2$  (u1'T   ��    ��� 
K����c� ǚB�S��g�|+�_��jAP< @��JA��3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
K����c� ÚB�W��c�|+�_��jAP< @��JA��3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
K����c� ÚB�W��_�|+�_��jAP< @��JA��3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
L ���c� ÙB�[��[�|+�_��jAP< @�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ���c� ��B�[�	pW�|+�_��jAP< @�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ���c� ��B�_�	pS�|+�_��jAP< @{�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ���c� ��B�_�	pO�|+�_��jAP< @{�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ��c� ��B�c�	pK�|+�_��jAP< @{�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ��c� ��B�c�	pG�|+�_��jAP< @w�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ��c� ��B�c�	�C�|+�_��jAP< @w�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ��c� ��B�g�	�?�|+�_��jAP< @w�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ��c� ��B�g�	�?�|+�_��jAP< @s�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ��c� ��B�k�	�;�|+�_��jAP< @s�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ��c� ��B�o�	�;�|+�_��jAP< @s�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
L ��c� ��B�o�	p7�|+�_��jAP< @o�JA��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
\$'_;� ǰA[�  �k�|é��)A\��-�Ls�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\$'_;� ǰA[�  �k�|ǩ��)A\��-�Lk�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\$(_;� ǰA[�  �k��Ǩ��)A\��-�Lg�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\$(_7� ǰA[�  �k��Ǩ��)A\��-ߜLc�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\$(_7� ǰA[�  �k��˧��*A\��-ۜL_�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\$(_7� ǰA[�  �k��˧��*A\��ۜL[�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\$(_7� ǰA[�  �k��Ϧ��*A\��לLW�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\$(_7� ǯA[�  �k��Ϧ��*A\��לLS�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\$(_7� ǯA[�  �k��ӥ��*A\��ӜLO�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\$(_3� ǯA[�  �k��ץ��*A\��ӜLK�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\$(_3� ǯA[�  �k�|פ��*A\��ϜLG�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\((_3� ǯA[�  �k�|ۤ��*A\���ϜLC�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\((_3� ǯA[�  �k�|ۣ��*A\���˜L?�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\()_3� ǯA[�  �k�|ߣ��*A\���ǜL;�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\()_/� ǯA[�  �k�|ߢ��*A\���ǜL7�"���T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\()_/� ǯA[�  �k�|���*A\���ÜL3�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\()_/� ǯA[�  �k�|���*M���K�/�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\()_/� ǯA[�  �k�|���*M���K�+�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\()_/� ǯA[�  �k�|���*M���K�'�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\,)_/� ǯA[�  �k�|���*M���K�'�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\,)_+� ǯA[�  �k�|���*M���K�#�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\,)_+� ˯A[�  �k�|���*M���K��3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\,)_+� ˯A[�  �k�|���*M���C��3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\0)_+� ˯A[�  �k�|���*M�����C��3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\0)_+� ˯A[�  �k�����*M�����C��3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\0)_+� ˯A[�  �k������*M�����C��3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\4)_+� ˮA[�  �k������*M,�����C��"s��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\4)_'� ˮA[�  �k������)M,�����EM�"s��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\4*_'� ˮA[�  �k������)M,�����EM�"s��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\8*_'� ˮA[�  �k������(M,�����EL��"s��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\8*_'� ˮA[�  �k������(M,�����EL��"s��T0 k� ���#KP 4a2$  (u1'T  ��_  ����8\8*_'� ˮA[�  �k�����'M,����EL��"s��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\<*_'� ˮA[�  �k�����&M,���{�E<��"s��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\<*_'� ˮA[�  �k�����&M,���w�E<��"s��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\<*_'� ˮA[�  �k�����&M,��o�E<��"s��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\@*_#� ˮA[�  �k���� %M��k�E<��"s��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\@*_#� ˮA[�  �k���� %M��g�E<��"s��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\@*_#� ˮA[�  �k����$M��c�E<��3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\D*_#� ˮA[�  �k����#M��[�E<��3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\D*_#� ˮA[�  �k����"M��W�E<��3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\D*_#� ˮA[�  �k����!M��S�E<��3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\H*_#� ˮA[�  �k����!M��O�E<ӿ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\H*_#� ˮA[�  �k���� M��O�E<Ͼ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\H*_#� ˮA[�  �k����M��K�E<˽3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\L*_� ˮA[�  �k����A\��K�E,Ǽ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\L+_� ˮA[�  �k���� A\��G�E,ǻ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\L+_� ˮA[�  �k���$A\��G�E,ú3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\P+_� ˮA[�  �k���(A\��C�E,��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\P+_� ˮA[�  �k���,A\��-C�E,��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\P+_� ˮA[�  �k���0A\��-?�E,��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\P+_� ˮA[�  �k���4A\��-?�E,��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\T+_� ˮA[�  �k���8A\��-;�E,��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\T+_� ˮA[�  �k���<A\��-;�E,��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\T+_� ˮA[�  �k���@A\��-7�E,��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\X+_� ˮA[�  �k���DA\��-7�E,��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\X+_� ˮA[�  �k���HA\��-3�E,��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\X+_� ˭A[��  �k���LA\��-3�E,��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\X+_� ˭A[��  �k����TA\��-3�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\\+_� ˭A[��  �k����XA\��-/�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\\+_� ˭A[��  �k����\A\��-/�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\\+_� ϭA[��  �k����`A\��-+�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\\+_� ϭA[��  �k����`A\��-+�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\`+_� ϭA[��  �k����dA\��-+�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\`+_� ϭA[��  �k����dA\��-'�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\`,_� ϭA[��  �k����hA\��-'�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\`,_� ϭA[��  �k�}��lA\��-'�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\d,_� ϭA[��  �k�}��p
A\��-#�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\d,_� ϭA[��  �k�}��t
A\��-#�E��3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\d,_� ϭA[��  �k�|���t
A\��-�E���3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\d,_� ϭA[��  �k�|���|
A\��-�E���3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\d,_� ϭA[��  �k�|���	A\��-�E���3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\h,_� ϭA[��  �k�����	A\��-�E�Û3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\h,_� ϭA[��  �k�����A\��-�E�Ú3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\h,_� ϭA[��  �k�����M��-�E�Ǚ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\h,_� ϭA[��  �k������M��-�E�˙3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\h,_� ϭA[��  �k������M��-�E�˘3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\l,_� ϭA[��  �k�����M��-�E�ϗ3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\l,_� ϭA[��  �k�����M��-�E�ӗ3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\l,_� ϭA[��  �k�����M��-�E|ז3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\l,_� ϭA[��  �k���|�M��-�E|ז3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\l,_� ϭA[��  "�k���|�M��-�E|ە3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\l,_� ϭA[��  "�k���|�M��-�E|ߕ3��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\p,_� ϭA[��  "�k���|�M��-�E|�3��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\p,_� ϭA[��  "�k���|� M,��-�E|�3��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\p,_� ϭA[��  "�k������M,��-�E|�3��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\p,_� ϭA[��  "�k������M,��-�E|�3��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\p,_� ϭA[��  "�k������M,��-�E|�3��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\t,_� ϭA[��  "�k������M,��-�D��3��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\t,_� ϭA[��  "�k������M,��-�D��3��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\t-_� ϭA[��  "�k������M,���D��3��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\t-_� ϭA[��  "�k���\��M,���D��3��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\t-_� ϭA[��  �k���\��M,���D��3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\t-_� ϭA[��  �k�M�\��M���D��3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\t-_� ϭA[��  �k�M�\��M���D��3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\x-_� ϭA[��  �k�M�\��M���D��3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\x-_� ϭA[��  �k�M�\��M����E|�3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\x-_� ϭA[��  �k�M�\��M����E|�3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\x-_� ϭA[��  �k���]�M����E|�3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\x-_� ϭA[��  �k��#�]�M����E|�3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\x-_� ϭA[��  �k��#�]�M����E|�3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\x-_� ϭA[��  �k��'�]�M����El�3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\|-_� ϭA[��  �k��'�]�A\����El�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\|-_� ϭA[��  "�k��'�]�A\����El�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\|-_� ϭA[��  "�k��'�]�A\����El�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\|-_� ϭA[��  "�k��+�m�A\����El�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\|-_� ϭA[��  "�k��+�m�A\����D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\|-_� ϭA[��  "�k��+�m#�A\����D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\|-_� ϭA[��  "�k��+�m'�A\����D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\|-_� ϭA[��  "�k��+�m+�A\����D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  "�k��+�m/�M����D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  "�k��+�m/�M����D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  "�k��+�m3�M����D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  "�k��+�m7�M����D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k��+�m;�M��]�D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k��+�m?�M��]�D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k��+�m?�M��]�D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k��+�mC�M��]�D<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k�+�mG�M��]�L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k�+�mK�M��]�L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k�+�mK�M,��]�L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k�+�mO�M,��]�L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k�+�mS�M,���L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k�+�mS�M,���L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k�+�mW�M,���L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�-_� ϭA[��  �k�+�m[�M,���L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�+�m[�M,���L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�+�m_�M,���L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�+�mc�M,���L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�/�mc�M���L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�/�mg�M���L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-/�mg�M���L<�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-/�mk�M���LL�3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-/�mo�M���LL�3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-/�mo�M���LL�3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-3�ms�M���LL�3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-3�ms�M���LL�3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-3�mw�M���LL�3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-3�mw�A\���LL�3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-3�m{�A\���LL�3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-3�m{�A\���LL�3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-7�m�A\���LL�3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-7�m�A\���LL�3��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-7�m��A\���LL�3��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-7�m��A\���LL�3��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-7�m��A\���LL�3��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-7�]��A\���LL�3��T0 k� ���#[P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-7�]��A\���LL�3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-;�]��A\���LL�3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-;�]��A\���LL�3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-;�]��A\���LL�3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-;�]��A\���LL�3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-;����A\���LL�3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-;����A\���LL�3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-;����A\���LL�3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-?����A\���LL�3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-?����A\���LL�3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-?�}��A\���LL�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-?�}��A\���LL�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-?�}��A\���LL�3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-?�}��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-?�}��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-?�}��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-C�m��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-C�m��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-C�m��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-C�m��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-C�m��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-C�m��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-C�m��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-C�m��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ϭA[��  �k�-C�m��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ӬA[��  �k�G�]��A\���LLߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ӬA[��  �k�G�]��A\���L<ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ӬA[��  �k�G�]��A\���L<ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ӫA[��  �k�G�]��A\���L<ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ׫A[��  �k�G�]��A\���L<ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ׫A[��  �k�G�훷A\���L<ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ׫A[��  �k��G�훶A\���L<ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� תA[��  �k��G�헵A\���L<ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ۪A[��  �k��G�퓵A\���A�ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ۪A[��  �k��G�폴A\���A�ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ۩A[��  �k��G�폳A\���A�ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ۩A[��  �k��G�틲A\���A�ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ۩A[��  �k��G�퇲A\���A�ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ߩA[��  �k��G�탱A\���D�ߘ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ߨA[��  �k��G���A\���D�ߙ3��T0 k� ���#�P 4a2$  (u1'T  ��_   ����8\�._� ߨA[��  �k��G��{�A\���D�ߙ3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\�._� ߨA[��  �k��C��w�A\���D�ߚ3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\�._� ߨA[��  �k��C��o�A\���D�ߚ3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\�._� �A[��  �k��C��k�A\���D�ߚ3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k��C��k�A\���D�ߛ3��T0 k� ���$P 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k��C��k�A\���D�ߛ3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k��C��g�A\���D�ߛ3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k��C��c�A\���D�ߛ3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k�M?��_�A\����D�ߛ3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k�M;��[�A\����D�ۜ3��T0 k� ���#;P 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k�M;��[�A\����D�ۜ3��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k�M7��W�A\����D�ۜ3��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k�M7��S�A\����D�ۜ3��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k�M7�O�A\����D�ۜ3��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k�M3�O�A\����D�ۜ3��T0 k� ���#KP 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k�M3�K�A\����A�ۜ3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k�M/�G�A\����A�ۜ3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k��+�C�A\����A�ۜ3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k��+�	�C�A\����A�ۜ3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k��+�	�C�A\�����A�ۜ3��T0 k� ���#kP 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k��'�	�?�A\�����A�ۜ3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8\�/_� �A[��  �k��'�	�?�A\�����A�ۜ3��T0 k� ���#{P 4a2$  (u1'T  ��_   ����8@��2 ��� � @o8# o;�|  �+��(2AP<  ��A �#3� T0 k� �  � e2$  (u1'T   ��/    �   2@��2 ��� � @o8# o;�|  �+��(2AP<  ��A �#3� T0 k� �  � e2$  (u1'T   /�/    �   2@��2 ��� � @o8# o;�|  �+��(2AP<  ��A �#3� T0 k� ������e2$  (u1'T   ��/    �   2@��2 ��� � @o8# o;�|  �+��(2AP<  ��A �#3� T0 k� ������e2$  (u1'T   ��/    �   2@��2 ��� � @o8# o;�| @+�@(2AP< P��A �#3� T0 k� ������e2$  (u1'T   ��/    �   2@��2 ��� � @o8# o;�| @+�@(2AP< P��A �#3� T0 k� ������e2$  (u1'T   ��/    �   2@��2 ��� � @o8# o;�|  @+�@(2AP< P��A �#3� T0 k� ������e2$  (u1'T   ��/    �   1@��2 ��� � @o8" o;�|  @+�@(2AP< P��A �#3� T0 k� ������e2$  (u1'T   ��/    �   1A_�2 ��� � CO8" o;�|$ @+�@(2AP< P��C@�"3� T0 k� ������e2$  (u1'T   ��/    �   0A_�2 o�� � CO8" ;�|$  +� (2AP< ���C@�"3� T0 k� ������e2$  (u1'T   ��/    �   0A_�2 o�� � CO8" ;�|$  +� (2AP< ���C@�"3� T0 k� ������e2$  (u1'T   ��/    ��� 0A_�2 o�� � CO8! ;�|$  +� (2AP< ���C@�!3� T0 k� ������e2$  (u1'T   ��    ��� 0A_�2 o�� � CO8! ;�|(  '� (2AP< ���C@�!3� T0 k� ������e2$  (u1'T   ��    ��� 0A��2 o�� o� CO8  ;�|(  '� (2AP< ���C@�!3� T0 k� ������e2$  (u1'T   ��    ��� 0A��2 o�� o� CO8 O;�|+��'� `(2AP< ���C@� 3� T0 k� ������e2$  (u1'T   ��    ��� 0A��2 o�� o� CO8O;�|+��� `(2AP< ���C@�3� T0 k� ������e2$  (u1'T   ��    ��� 0A��2 o�� o� E�8O;�|+��� `(2AP< ���C@�3� T0 k� ������e2$  (u1'T   �    ��� .A��2 o�� o� E�8O;�|+��� `(2AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� -A��2 o�� �� E�8O;�|+��� `(2AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� ,A��2 o�� �� E�8�;�|+�P�@(2AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� +A��2 o�� �� E�8�;�|+�P�@(3AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� *A��2 o�� �� E�8�;�|+�P�@(3AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� )A��2 o�� �� E�8�;�|+�P�@(3AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� (BO�2 o��O� E�8�;�|+�P�@(4AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� 'BO�2 o��O�E�8�;�|+�P�@(4AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� &BO�2 o��O�E�8�;�|+�P�@(5AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� %BO�2 o��O�E�8�;�|+�P�@(5AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� $BO�2 o��O�E�4�;�|+�P�@(6AP< ���CP�3� T0 k� ������e2$  (u1'T   ��    ��� #@�2 o��O�E�4�;�|+�P��(6AP< ���IP�3� T0 k� ������e2$  (u1'T   ��    ��� "@�2 o��O�E�4;�|+�P��(7AP< ���IP�3� T0 k� ������e2$  (u1'T   ��    ��� !@�2 o��O�E�0;�|+�_���(8AP< ���IP�3� T0 k� ������e2$  (u1'T   ��    ���  @�2 o��_�E�0;�|+�_���(9AP< ���IP�3� T0 k� ������e2$  (u1'T   ��    ��� @�2 o��_�E�,;�|+�_���(:AP< `��IP�3� T0 k� ������e2$  (u1'T   ��    ��� B��2 o��_�E�(o;�|+�_���(;AP< `��IP�3� T0 k� ������e2$  (u1'T   ��    ��� B��2 o��_�E�(o;�|+�_���(<AP< `��I`�3� T0 k� ������e2$  (u1'T   ��    ��� B��2 o��_�	E�$o;�|+�_���(=AP< `��I`�3� T0 k� ������e2$  (u1'T   ��    ��� B��2 o��/�
E� o;�|+�_���(>AP< `��I`�3� T0 k� ������e2$  (u1'T   ��    ��� B��2 o��/�E� o7�|+�_���$?AP< 0��I`�3� T0 k� ������e2$  (u1'T   ��    ��� E��2 o��/�E�	o7�|+�_���$AAP< 0��I`�
3� T0 k� ������e2$  (u1'T   ��    ��� E��2 o��/�E�o3�|+�_���$BAP< 0��E0�	3� T0 k� ������e2$  (u1'T   ��    ��� E��2 o��/�E�o3�|+�_��� DAP< 0��E0�	3� T0 k� ������e2$  (u1'T   ��    ��� E��2 o��/�Eoo/�|+�_��� EAP< ��E0�3� T0 k� ������e2$  (u1'T   ��    ��� E��3 o��/�Eoo/�|+�����FAP< ��E0�3� T0 k� ������e2$  (u1'T   ��    ��� E��3 o��/�Eoo+�|+�����GAP< ��E0�3� T0 k� ������e2$  (u1'T   ��    ��� E� 4 o���Eoo'�|+�����JAP< ��E �3� T0 k� ������e2$  (u1'T   ��    ��� D�4 o���Eo?'�|+�����KAP< ��E �3� T0 k� ������e2$  (u1'T   ��    ��� D�5 o���E?#�|+�_���LAP< ��E �3� T0 k� ������e2$  (u1'T   ��    ��� D�5 o���E ?�|+�_���NAP< ��E �3� T0 k� ������e2$  (u1'T   ��    ��� D�6 o���E�?�|+�_���OAP< ��E � 3� T0 k� ������e2$  (u1'T   ��    ��� D�7 o����E�o�|+�_���RAP<  ��E ��3� T0 k� ������e2$  (u1'T   ��    ��� D� 8 o����E�o�|+�_���SAP<  ��E ��3� T0 k� ������e2$  (u1'T   ��    ��� D�$9 o���E�o�|+�_��� UAP<  ��E ��3� T0 k� ������e2$  (u1'T   ��    ��� D�(: o{���E�o�|+�_����VAP<  ��E��3� T0 k� ������e2$  (u1'T   ��    ��� D�,: o{���E~��o�|+�_����XAP<  ��E��3� T0 k� ������e2$  (u1'T   ��    ��� D�0; ow��� E~��o�|+�_����YAP<  ��E��3� T0 k� ������e2$  (u1'T   ��    ��� D�8< os���!E~���|+�_����[AP<  ��E��3� T0 k� ������e2$  (u1'T   ��    ��� 
D�@> oo���#E����|+�_����^AP<  ��J@��3� T0 k� ������e2$  (u1'T   �    ��� 
D�H? ok�� $E����|+�_����_AP< @��J@��3� T0 k� �����e2$  (u1'T   �    ��� 
D�L@ og��%E����|+�_���aAP< @��J@��3� T0 k� �{���e2$  (u1'T   ��    ��� 
D�TA oc��%E�����|+�_���bAP< @��J@��3� T0 k� �w��{�e2$  (u1'T   ��    ��� 
D�XB oc��&E�����|+�_���dAP< @��J@��3� T0 k� �w��{�e2$  (u1'T   ��   ��� 
E�`C o_�'F����|+�_���eAP< @��J@��3� T0 k� �s��w�e2$  (u1'T   ��    ��� 
E�dD o[�(F����|+�_���gAP< @��J@��3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
E�lE o[� )F�����|+�_���hAP< @��J@��3� T0 k� �o��s�e2$  (u1'T   ��    ��� 
E�tE oW�$*F����|+�_��iAP< @��J@��3� T0 k� �k��o�e2$  (u1'T   ��    ��� 
E�xF oS�,+F����|+�_{��kAP< @��J@��3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
E��G oS��0+E�����|+�_w��lAP< @��J@��3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
E��H oO��8,E�����|+�_w��mAP< @��J@��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E��I oO��<-E�����|+�_s��oAP< @��J@��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E��J oK��D-E�����|+�_o��pAP< @��J@��3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E��J oG��H.E�����|+�_k��qAP< @��J@��3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
E��K oG��P.E�����|+�_k��rAP< @��JA�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
E��K oC��T/E�����|+�_g��sAP< @��JA�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
E��L oC��\/E�����|+�_c��uAP< @��JA�3� T0 k� �W��[�e2$  (u1'T   ��    ��� 
E��L oC��d0E�����|+�__��vAP< @��JA�3� T0 k� �W��[�e2$  (u1'T   ��    ��� 
E��M oC��h0E����|+�__��wAP< @��JA�3� T0 k� �W��[�e2$  (u1'T   ��    ��� 
E��M oC��p0E����|+�_[��xAP< @��JA�3� T0 k� �W��[�e2$  (u1'T   ��    ��� 
E��M oC�pt1B����|+�_W��yAP< @��JA�3� T0 k� �W��[�e2$  (u1'T   ��    ��� 
E��N oC�p|1B����|+�_W��yAP< @��JA�3� T0 k� �W��[�e2$  (u1'T   ��    ��� 
E��N oG�p�1B����|+�_S��yAP< @��JA�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
E��N oG�p�1B����|+�_O��xAP< @��JA�3� T0 k� �[��_�e2$  (u1'T   ��    ��� 
E��N oG�p�1B����|+�_O��xAP< @��JA�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
E��N oG�p�1B����|+�_K��xAP< @��JA�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
E� N oG�p�1K����|+�_G��xAP< @��JA�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
E�N oG�p�0K����|+�_G��wAP< @��JA�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
E�M oG�p�0K����|+�_C��wAP< @��JA�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
E�M oG�p�0K����|+�_C��wAP< @��JA�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
CAM oG���/K����|+�_C��wAP< @��JA�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
CA$L oK���/K���#�|+�_C��vAP< @��JA�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
CA,L oK���/K���'�|+�_C��vAP< @��JA�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
CA0K oK���.K���/�|+�_C��vAP< @��JA�3� T0 k� �_��c�e2$  (u1'T   ��    ��� 
CA8K oK���.K���3�|+�_C��vAP< @��JA#�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�@J oK���-K���7�|+�_C��vAP< @��JA#�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�DJ oK���,K���;�|+�_C�|uAP< @��JA#�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�LI oK���,K���?�|+�_?�|uAP< @��JA'�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�PH oK���+K���G�|+�_?�xuAP< @��JA'�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�XG oK���*K���K�|+�_?�xuAP< @��JA'�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�\F oK���)K���O�|+�_?�tuAP< @��JA+�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�dE oK���(K���W�|+�_?�ttAP< @��JA+�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�hD oK���'K���[�|+�_?�ptAP< @��JA+�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�pC oO���'K���c�|+�_?�ptAP< @��JA/�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�tB oO���&K���g�|+�_?�ltAP< @��JA/�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E�xA oO���$K���o�|+�_?�ltAP< @��JA/�3� T0 k� �c��g�e2$  (u1'T   ��    ��� 
E��@ oO�� #K���s�|+�_?�hsAP< @��JA/�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
E��? oO�q"K���{�|+�_?�hsAP< @��JA3�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
E��= oO�q!K����|+�_?�dsAP< @��JA3�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
E��< oO�q K�����|+�_?�dsAP< @��JA3�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
E��; oO�qK�����|+�_?�dsAP< @��JA7�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
E��: oO�qK�����|+�_?�`sAP< @��JA7�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
E��8 oO�qK�����|+�_?�`rAP< @��JA7�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
E��7 oO�qK������|+�_;�\rAP< @��JA7�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
E��6 oO�q K������|+�_;�\rAP< @��JA;�3� T0 k� �g��k�e2$  (u1'T   ��    ��� 
                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��4r ]�)�)� � ����T  � �     � ;��    ��� ;��    �x��             �� 
          ���    ���   	          ��p�   � �
	   ���t    ��p���q       -           v �� 
�        ���  #  ���  0
&         ����   � �
	    ,h/    ��� ,�    ���N   	        u�� 
         ��    ���   8
         ����  + +      ����    �����+/    ��/             M
 �� 
           )��    ���   @

          ����   � �	    . �C    ��պ �    !��   	           
		�� 
          �0�     ���  8	          ��4�  ��      B�
�Z    ��4��
�Z                             ���@               �  ���     

 0            ��U�         V���    ��b��랍    �?"              	   �8         �     ��@   8(          j9�        j��h�     j<���r�    ���j             	 ���8         ��     ��@   8
           �   	    ~ H�      � H�                  	    �8         �@     ��J    

'		          ����  $ $       � �    ��� Bt    
�N               �� �         	 ��     ��@   X
	         ��;� � �
    � gd�    ��b6 gM�    ��Y                   �         
 �
`     ��P   8
            � ��     � ��       � ��                            �����              �  ��@    0 0                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��R  ��        ���6�    ��R��3�       - "                x                j  �       �                         ��    ��        ���      ��  ��           "                                                �                          ;�� ,�� �
����   g �������         	 
       
  x   |W� ���F       �� e� �� _@ � _` �$  _� �d _� �� _� �� _� �� b  �  b@ D� `e� E�  f� E�  f� � n@ � �t� �  u� � �r@ �  s@ 
�< V� 
� V� 
�\ W  �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� � }`���� � 
�| V  
�| V� 
�� V� 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� 
 ������  ������  
�fD
��L���"����D" � j  "  B   J jF�"     
�j � � 
��
��
��"     "�j��   * �
� �  �  
� ��    ��     ���      ��    ��     ���            ��     �           � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �&&'      �� T ���        � �T ���        �        ��        �        ��        �    ��    ��l B��        ��                         T�) ,   ���                                     �                ����             �������%��  �� 
 2               27 Jeremy Roenick      1:39                                                                        3  2      �!cjj9crzB� � � B� � B� � �B� � � B� � � B� � 	� � 
� �K � K" � �cV � c^ � � . � �C/ � �C7 � � C9 � �k~  � k�  �c� � � c� � �C � � C � � C � � C � � C � � C � �J� � �J� � � J� � �  J� � w!k� � "k� �  #k� �-$"� �- %"� �&� �'
� �-("� �- )"� �*"� �+*� � �,"� � � -"� �.� � � 
� � 
�1"2 t02"6 t03"
 �8 4"L �P 5"R �X  "K �07"6 t08"
 �8 9"L �P :"R �X  "K �X  "K �` =*G\`  *K<_  *G\                                                                                                                                                                                                                         �� R @       �     @ 
         �     W P E e  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    ��   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, <  6 )  � @��@Q��@���A#� �4�h �)��                                                                                                                                                                                                                                                                                                                   �                                                                                                                                                                                                                                                   �    ,     �   :�J      �                             ������������������������������������������������������                                                                    
                                                                  �    �    �        p      p�                   
     ���������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ����                         
       �   ! !    ��  4�J      	u  	                           ������������������������������������������������������                                                                                                                        
                   ]  �   )            �      �  ��               	 
     � ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� ������������������                                                                                                                                                                                                                                                             
                                        	                    �             


             �  }�                    +#        V                                                           ��������    ��������������������������������  R}��������������������     N�����������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" A C 6                                 � 5Hq� �\                                                                                                                                                                                                                                                                                            )n)n1n  )�1F                m      m      m                        k                                                                                                                                                                                                                                                                                                                                                                                                                > �  	>�  J�  @#�  H#�  Cm�  �̞����� ������p������̎���̎�� �N �����|                ���   S p        �   & AG� �  �                 �                                                                                                                                                                                                                                                                                                                                        K N   �                      !��                                                                                                                                                                                                                            Y��   �� �� ��      �� 6      ���������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ����� ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� ������������������             $����������������˪�������������������������������������f��ff��ff�������̺�ff�fffffffffffffffffff����ƹ��ffʻfff�fffjffffffffffff��������������������ʺ��l���f˪������������������������������������������������������������������fff�fff�fff�ffk�ffi�ff��ff��ff�ffffffff�fff�x�����w��xx�������wfffffff�ffff�fffww��ww�x����wx��fk��ff��ff��ffʹffj��fʪ�f�ˊ�k������������ʚ��������������������������������������������˫��ʫ��ff��fl��fl��ff̫fff�ffʬ�f���f�����������wu���w��l������f����W��������xww��Wy�l����x������k���W�fi���j���j���f����˘�����y�y�y����������������������������������������������������ʻ����ʫɚ�����l���ƨ�lƘ�j���k���̜i���j���kxx���wx������wx������������ƈx����������������wW����w�������������������������z����������˫��̺������������������������������������������������������������ʺ������k������������������������������������������x�j���˙�x�˘��̩�x������x���xx�x������x������wx���˫��ʫ����������˪�����ʻ��������������������������������������ʻ�ʻ�����ʪ̫����˺��������������������˪�����f���k��f��fǶW�g���k���̻���f������������������x�������˩f̺�����uw�����w��x�wXx��˪�����������l����l���i��ƹx�f�������������������ʫUW��UUU�UUUX      ?      2     ��                       7     �   �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p��  5� � ��    �@���6 ��  �@���6 �$ ^$ �r@  �@  �r@   5 
�V ��   5 
   ���  ��   ���  �$ ^$   �        8 
e �� 8 � �$���  � ��� �� � ��� � �� � � ��� �  �      �      �������2����   g���        f ^�         �� ���            ��4����2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                               	                 �  ��� �UU���U              �	���UUU�UUUUUU      	� ��U�UUUUUUUUUUUUUUUUUUU    ��� U^��UUU�UUU^UUUUUUUUUUUU            �   �   ^�  U�  UY�    � 	UU 	��  	�  	�  �^ 	��    �	UY�������UUUUUUU��UU��UU�U�UUUUUUUUUUUUUUUUUUUUUUUUUUUU^UUUYUU^�U^� U� ^�  �  ��  �   �   ��UU ��U �U  �U  ��            U^� UU� UU� UU� ���                    	   �       	   	   	    �UUU�UU���U  	�� �����U�UUU�UUUUUUYUUUYUUUYUUU^UUU^UUUUUUUUUUUU�   �   �   �   �   � �^���U^��            	����UUU�UUU�UUUUUU^            ��  U�  Y�  �  �      �   �   �   	                ���Y���U��Y�^�U��U ��^ 	� 	� UUUU�UUUUUUUU^�U^����� �        UUUUUUUUUUUUUUUUUUUU�������    UUU�UU^�UU�U� Y�  ��          �                               wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "" "  """ ""   "! " ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ ""   "! " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """"! "   "      ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        "  " �" ��" ��- �ۼ w۽��ݹ����� ��� ��  ˼  ��  ˼  ��  H�  �D  J�  J�  �  �  �  �  
�  �  �  �  ,�  " "" �" �"�   ˰  ��  wp ��ډ�v���r�̸��˰��� ��  ��  ��  ��  ̸  ��  ��  DC  C4@ T4@ T40 T30 T30 S;� H�  ��  ��  ��  ""  "  �""� "�/��        �   �   �      �  �   �   �   �   �              �   �   �   �             ���� �                        " "" """ �"  �   �   �                              � ��                  �  �˰ ��� �wp ���    �   ��  ���  � �    �                                                                                                                                      "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��                   � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                              �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��  ��  �   ��  �                  ��                                 � ���� ��   � � �                           �   �                                                                                                        �   �   �   �  
� 	�� �� ���	���
���	������+�ݼ� �  
C  �U  �T 
UC 
UT ED  �D  ��  �  �   " �"  �     �        �   ��  ��  ��  w�  ��  ��� ��� ̻� ̻���˩�̽��̽� ˉ� ��  340 UT0 DD0 330 33  C  C  
�  �  ,�  ""  "  �� ��     �      �   ��  �  ��  �             �  �   �   ��  �             ��  ��  �                            �   �    �   �       �   �   �                .                      ��� ���� �����                                                                                                                                                                                                 0 0#0  03  10         �  �  � 
�� ��} ˚w
���	����+� �+� ��� ",  "�  ". 34 DC3 DD3 �DC ��  ��  
"   "  "  ""  "!    �                    �   �   �   w   m�  g�� z�� ����̹���˙�̼̰������������蜚��L��>\���" ""  ""  �+ "	��"� �����.�"��"! "  ��           /   ��  �   �    �  ���  ��� ��  �                        �   �   �                            �   �   �   �   �      �                    ��� ���� ��                                                                                                                                                                                                                   �� �����ݼڜ��ک��ک��z�	��� 
�� 
�� 	�� ̘ ɪ  ��  �  �� �� ������������ ���  � � � �� �� ������ ��                      �   ��  ��  �̰ ��� ��˰�̻��̻���������ˉ�U��EP�ET �I� ٕ  �D� �L� ��� ��" ����/�"�"�""�����                         /�� �                                         �  ��  �� ��  ��                  �   ��� �̰       �  �� Ș ��  ��  �                                                                                                                                                                                                                                     	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                      �   �   �   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw     �����                     �"�!/"�  �                     �   ��  ���  � �    �                                                                                                                                                     �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �        �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                              "  .���"    �     �                                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  �   �   �   �   �       �     �"  "  �   "                                    �   �   �            �� �� �� g} �� vw                       �   �      ��   �  ��  �  �  �         � �������������  �                                �   �                                                                                                        �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �      �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                       � ��                  �  �˰ ��� �wp ���      � �������������  �                                                                                                                                             �   �   �   � 
�w ��� ș����	���
���	������ ݼ� ݼ� �� �� 	�� �� 3E 34 D@ ��  ��  ʢ  ""� "/  ��� �      �    �   ��  ��  �p  �p  w   ��  ��� ��� ��� ˻� ̼˰��ː�۹�̽��̽����˸� "��@ DJ� EZ� DU� EZ  DL̘ 	�������" �""�"/��"� ��                    � ��� "  �         �    �  �       �   �   ��  �   �   �   �       ����   �       �                                   �    ���  ��                    ��  ��  ���              �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                                           �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                     �                             �   �   �   �   �   �                                                                                                                                                �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""��������������������""""������DDM�D��""""�������MM�M�M""""��������DD�A��""""�������MAA�MA""""��������AA�A""""����������M�MA""""������������M���M���M���"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUQUUQUUUUUUQUUUUUUUU3333DDDDUUUUDEEDDTEUUUU3333DDDDAEAEQQUDTDUUUU3333DDDDQUQUQDUDDUUUU3333DDDDAADAUAUEDUTUUUU3333DDDDADAEAQAUEDUTUUUU3333DDDDUDUQEUQUUQUEUDUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=""""��������AA�A    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ADA�LL��L�D����3333DDDD x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(XxLL����������D����3333DDDD w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""����������A������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(""""�������I�I������ �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�""""�������I��D���I������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`�D�M�D���M������3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(MD�M�A�����MD�����3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(�""""�����AMAD������ � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(�""""������������������ � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(��H��J�AD�DH�D����3333DDDD � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(�""""�������DD����� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq!cjj9crzB� � � B� � B� � �B� � � B� � � B� � 	� � 
� �K � K" � �cV � c^ � � . � �C/ � �C7 � � C9 � �k~  � k�  �c� � � c� � �C � � C � � C � � C � � C � � C � �J� � �J� � � J� � �  J� � w!k� � "k� �  #k� �-$"� �- %"� �&� �'
� �-("� �- )"� �*"� �+*� � �,"� � � -"� �.� � � 
� � 
�1"2 t02"6 t03"
 �8 4"L �P 5"R �X  "K �07"6 t08"
 �8 9"L �P :"R �X  "K �X  "K �` =*G\`  *K<_  *G\3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������=�N�K�U�X�K�T��0�R�K�[�X�_� � � � � � �-�1�B�������������������������������������������1�G�X�_��<�[�Z�K�X� � � � � � � � � � �-�1�B�����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������-�2�3� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�1�B� ��!������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            