GST@�                                                           �`�                                                      ���                       ���2���2
 ʲ����������8���~���        �h     #    ~���                                d8<n    �  ?     r����  �
fD�
�L���"����D"� j   " B   J  jF�"     "�j  " ���
��
�"    B�jl �   B ��
  �                                                                               ����������������������������������       ��    =bo 0Q 4g 11  4              	� 
                     �� � �  �                 �n� 	)         88�����������������������������������������������������������������������������������������������������������������������������o  b  o   1  +    '           �                  	  7  V  	                  E  "          := �����������������������������������������������������������������������������                                ��  �   o   f�   @  #   �   �                                                                                '     	�)n�  "E    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E f �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    M�}ۼD��E��; m��� �k��MD�����=\2Z3�T0 k� ��C��C(%2't �8t B  ��G    � �8M�}�D��E��:-��� �k��ND�#����-T3Z3�T0 k� ��@��@(%2't �8t B  ��G    � �8M�}�D��E��9-��� �k��ND�'����-P4Z3�T0 k� ��>��>(%2't �8t B  ��G    � �8M�}��D��E��8-��� �g��OD�+����-D7Z3�T0 k� ��?��?(%2't �8t B  ��G    � �8]�}��D��E��7-��� �c��OD�/����-@9Z3�T0 k� ��@��@(%2't �8t B  ��G    � �8]�~�E�E��6-��� �c��OD�/�޷�-<:Z3�T0 k� ��@��@(%2't �8t B  ��G    � �8]�~�E#�E��5-��� �_��PD�3�ޯ�-8<Z3�T0 k� ��@��@(%2't �8t B  ��G    � �8]�~�E'�E��3��� �[��PD�7�ޣ�-0?Z3�T0 k� ��A��A(%2't �8t B  ��G    � �8]�~'�E+�E��2��� �W�� PD�8 ޛ�-,@Z3�T0 k� ��A��A(%2't �8t B  ��G    � �8]�~+�E/�E��1��� �S�� PD�<ޓ�-(BZ3�T0 k� ��A��A(%2't �8t B  ��G    � �8]�~3�E3�E��0��� �O���PI�<ޏ�-$CZ3�T0 k� ��A��A(%2't �8t B  ��G    � �8]�n?�E;�E��.��� �G���PI�@ޏ�$CZ3�T0 k� ��A��A(%2't �8t B  �G    � �8]�nG�Eo;�E��.�� ^C���PI�D
^��$DZ3�T0 k� ��A��A(%2't �8t B  �G    � �8m�nK�Eo?�E��-�� ^C���PI�D^�� EZ3�T0 k� ��A��A(%2't �8t B  ��G    � �8m�nW�EoC�E��+�� ^G�\�QI�H^��FZ3�T0 k� ��G��G(%2't �8t B  ��G    � �8m�n_�EoG�E��*�� ^G�\�QI�L^� GZ3�T0 k� ��K��K(%2't �8t B  ��G    � �8m�nc�EoG�E��)�� ^G�\�QI�L^{� HZ3�T0 k� ��O��O(%2't �8t B  ��G    � �8m�ng�EoG�E��(�� ^G�\�QI�P^{� HZ3�T0 k� ��Q��Q(%2't �8t B  ��G    � �8m�nk�EoK�E��'��� ^G�\�QI�P^w� IZ3�T0 k� ��S��S(%2't �8t B  ��G    � �8m�no�EoK�E��'��� ^G���QA�T^s� JZ3�T0 k� ��M��M(%2't �8t B  ��G    � �8m�ns�EoK�E��&��� ^G���QA�T^o� JZ3�T0 k� ��H��H(%2't �8t B  ��G    � �8m�^w�D?K�E��%��� ^K��QA�X^k� KZ3�T0 k� ��D��D(%2't �8t B  ��G    � �8m�^{�D?O�E��%��� ^K��QA�X^g� LZ3�T0 k� ��A��A(%2't �8t B  ��7    � �8}�^��D?O�El�$��� ^K��QA�\^c� MZ3�T0 k� ��>��>(%2't �8t B  ��7    � �8}�^��D?O�El�#��� ^K��QA�\ ^_� MZ3�T0 k� ��=��=(%2't �8t B  ��7    � �8}�^��D?O�El�#��� ^O��PA�`"^[� NZ3�T0 k� �|<��<(%2't �8t B  ��7    � �8}�^��D?O�El�"��� ^O��PA�`#^[� NZ3�T0 k� �x;�|;(%2't �8t B  ��7    � �8}�^��D?O�El�"��� ^O��PA�d%^W� OZ3�T0 k� �p:�t:(%2't �8t B  ��7    � �8}�^��D?K�El�!��� ^O��OA�d&^S�  PZ3�T0 k� �h9�l9(%2't �8t B  ��7    � �8}�^��D?K�El�!��� ^S���OA�d'^O�  PZ3�T0 k� �p8�t8(%2't �8t B  ��7    � �8}�^��D?K�El� ��� ^S���NA�h)^O�  QZ3�T0 k� �t8�x8(%2't �8t B  ��7    � �8}�N��D?K�El� ��� ^S��xNA�h*^K� �QZ3�T0 k� �t7�x7(%2't �8t B  ��7    � �8}�N��DOG�El���� ^S��pMA�l+^G� �RZ3�T0 k� �t7�x7(%2't �8t B  ��7    � �8M�N��DOG�A����� ^S��lMA�l-^G� �RZ3�T0 k� �p6�t6(%2't �8t B  ��7    � �8M�N��DOG�A����� ^W��dLA�l.^C� �SZ3�T0 k� �p5�t5(%2't �8t B  ��7   � �8M�N��DOC�A����� ^W��`KA�p/^?� �SZ3�T0 k� �l5�p5(%2't �8t B  ��7    � �8M�N��DOC�A����� ^W��XJA�p0^?� �TZ3�T0 k� �h4�l4(%2't �8t B  ��7    � �8M�N��DO?�A����� ^W��TIA�p2^;� �TZ3�T0 k� �`3�d3(%2't �8t B  ��7    � �8M�N��DO;�E���� ^W��PHA�t3^7� �UZ3�T0 k� �\2�`2(%2't �8t B  ��7    � �8M�N��DO;�E���� ^[��HHA�t4^7� �UZ3�T0 k� �T1�X1(%2't �8t B  ��7    � �8M����DO7�E���� ^[�DGA�t5^3� �VZ3�T0 k� �X2�\2(%2't �8t B  ��7    � �8M����DO7�E���� ^[�@EA�x6^3� �VZ3�T0 k� �\2�`2(%2't �8t B  ��7    � �8M����DO3�E���� ^[�8DA�x7^/� �WZ3�T0 k� �\2�`2(%2't �8t B  ��7    � �8M����D_/�E����� ^[�4CA�x8^+� �WZ3�T0 k� �X2�\2(%2't �8t B  ��7    � �8M����D_+�E���#�� ^_�0BA�|:^(  �WZ3�T0 k� �X1�\1(%2't �8t B  ��7    � �8]�N��D_'�E���#�� ^_�,AA�|;^$ �XZ3�T0 k� �X0�\0(%2't �8t B  ��7    � �8]�N��D_'�E���#�� ^_�(@A�|<^$ �XZ3�T0 k� �h3�l3(%2't �8t B  �7    � �8]�N��D_#�E���#�� ^_��$?A��=^  �YZ3�T0 k� �t5�x5(%2't �8t B  ��?    � �8]�N��D_�E|��#�� ^_�� >A��>^  �YZ3�T0 k� ��7��7(%2't �8t B  ��?    � �8]�N��D_�E|��'�� ^_��=A��?^ �ZZ3�T0 k� ��9��9(%2't �8t B  ��?    � �8]�>��D_�E|��'�� ^c��<A��@^ �ZZ3�T0 k� ��;��;(%2't �8t B  ��?    � �8]�>��D_�E|��'�� ^c��;A��A^ �ZZ3�T0 k� ��;��;(%2't �8t B  ��3    � �8]>��D_�E|��'�� ^c��:A��B^ �[Z3�T0 k� ��:��:(%2't �8t B  ��3    � �8]>��D_�El��+�� ^c��9A��C^ �[Z3�T0 k� ��6��6(%2't �8t B  ��3    � �8]>��DoEl��+�� ^c��8A��C^ �[Z3�T0 k� ��3��3(%2't �8t B  ��3    � �8]N�Do El��+�� ^c��7A��D^	 �\Z3�T0 k� �|1��1(%2't �8t B  ��3    � �8m
N�Dn�El��+�� ^g��6A��E^
 �\Z3�T0 k� �t1�x1(%2't �8t B  ��3    � �8mN�Dn�El��+�� ^g�� 5A��F^
 �]Z3�T0 k� �h0�l0(%2't �8t B  ��3    � �8mN{�Dn�	A���/�� ^g�	�4A��G^ �]Z3�T0 k� �`/�d/(%2't �8t B  ��3    � �8mN{�En�A���/�� ^g�	�3A��H^ �]Z3�T0 k� �X/�\/(%2't �8t B  ��3    � �8mNw�En�A���/�� ^g�	�2A��I^ �^Z3�T0 k� �T.�X.(%2't �8t B  ��3    � �8mNw�En�A�| �/�� ^g�	�1A��J^ �^Z3�T0 k� �P.�T.(%2't �8t B  ��3    � �8mNw�En�A�| �/�� ^g�	�0A��J^ �^Z3�T0 k� �L-�P-(%2't �8t B  ��3    � �8�Ns�En�L<x!�3�� ^k�	�/A��K^ �_Z3�T0 k� �T*�X*(%2't �8t B  ��3    � �8�Ns�En�L<t!�3�� ^k�	�.A��L^  �_Z3�T0 k� �\'�`'(%2't �8t B  ��3    � �8�Ns�En�L<t!�3�� ^k�	�.A��M^  �_Z3�T0 k� �\%�`%(%2't �8t B  ��3    � �8�No�En�L<p"�3�� ^k�	�-A��M]� �`Z3�T0 k� �\%�`%(%2't �8t B  ��3    � �8�!^o�E^�L<l"�3�� ^k�	�,A��N]� �`Z3�T0 k� �`$�d$(%2't �8t B  ��3    � �8�#^o�E^�L<l#�3�� ^k�	�+A��O]� �`Z3�T0 k� �`#�d#(%2't �8t B  ��3    � �8�%^k�E^� L<h#�7�� ^k�	�*A��P]� �`Z3�T0 k� �\#�`#(%2't �8t B  ��3    � �8�'^k�E^�"L<d#�7�� ^o�	�+A��P]� �aZ3�T0 k� �\#�`#(%2't �8t B  ��3    � �8�)^k�E^�#L<d$�7�� ^o�	�+A��Q]� �aZ3�T0 k� �X$�\$(%2't �8t B  ��3    � �8�*�g�L�%L<`$�7�� ^o�	�+A��R]� �aZ3�T0 k� �T$�X$(%2't �8t B  ��3    � �8�,�g�L�'LL\$�7�� ^o�	�,A��S]� �bZ3�T0 k� �T$�X$(%2't �8t B  ��3    � �8�.�c�L�)LL\%�7�� ^o�	�,A��S]� �bZ3�T0 k� �P%�T%(%2't �8t B  ��3    � �8�0�c�L�+LLX%�;�� ^o�	�,A��T]� �bZ3�T0 k� �L%�P%(%2't �8t B  ��3    � �8�1�_�L�,LLX%�;�� ^o�	�-A��U]� �bZ3�T0 k� �L%�P%(%2't �8t B  ��3    � �8�3�_�L�.LLT&�;�� ^o�	�-A��U]� �cZ3�T0 k� �H&�L&(%2't �8t B  ��3    � �8�5�[�L�0LLT&�;�� ^o�	�-A��V]� �cZ3�T0 k� �H&�L&(%2't �8t B  ��3    � �8�6�W�L�2LLP&�;�� ^s��.A��V]� �cZ3�T0 k� �D&�H&(%2't �8t B  ��3    � �8�8�W�L�3LLL'�;�� ^s��.A��W]� �cZ3�T0 k� �D'�H'(%2't �8t B  ��3    � �8�9�S�L�5LLL'�;�� ^s��.A��X]� �dZ3�T0 k� �@'�D'(%2't �8t B  ��3    � �8�;�O�L.�6LLH'�?�� ^s��.A��X]� �dZ3�T0 k� �@'�D'(%2't �8t B  ��3    � �8�=�O�L.�8LLH'�?�� ^s��.A��Y]� �dZ3�T0 k� �<'�@'(%2't �8t B  ��3    � �8�>>K�L.�:LLD(�?�� ^s� �.A��Y]� �dZ3�T0 k� �8(�<((%2't �8t B  ��3    � �8�@>G�L.�;LLD(�?�� ^s� �.A��Z]� �eZ3�T0 k� �8(�<((%2't �8t B  ��3    � �8�A>G�L.�=LL@( n?�� ^s� �.A��[]� �eZ3�T0 k� �4(�8((%2't �8t B  ��3    � �8�B>C�L.�>LL@) n?�� ^s� �/A��[]� �eZ3�T0 k� �4)�8)(%2't �8t B  ��3    � �8�D>?�L.|@LL<) nC�� ^s� �/A��\]� �eZ3�T0 k� �0)�4)(%2't �8t B  ��3    � �8�E>?�L.xALL<) nC�� ^w� �/A��\]� �fZ3�T0 k� �0)�4)(%2't �8t B  ��3   � �8�G>;�L.tBLL8) nC�� ^w� �/A��]]� �fZ3�T0 k� �0)�4)(%2't �8t B  ��3    � �8�HN;�L.pDLL8*�C�� ^w���/A��]]� �fZ3�T0 k� �,*�0*(%2't �8t B  ��3    � �8�IN7�L.pELL8*�C�� ^w���/A��^]� �fZ3�T0 k� �,*�0*(%2't �8t B  ��3    � �8�KN3�L.lFLL4*�C�� ^w���/A��^]� �fZ3�T0 k� �(*�,*(%2't �8t B  ��3    � �8�LN3�L.hHLL4*�G�� ^w���/A��_]� �gZ3�T0 k� �(*�,*(%2't �8t B  ��3    � �8�MN/�L.dILL0+�G�� ^w���/A��_]� �gZ3�T0 k� �$+�(+(%2't �8t B  ��3    � �8�N�+�L.dJLL0+�G�� ^w���/A��`]� �gZ3�T0 k� �$+�(+(%2't �8t B  ��3    � �8�P�+�L.`LLL,+�G�� ^w���/A��`]� �gZ3�T0 k� � +�$+(%2't �8t B  ��3    � �8�Q�'�L.\MLL,+�G�� ^w���/A��a]�  �gZ3�T0 k� � +�$+(%2't �8t B  ��3    � �8�R�#�L.XNLL,,�G�� ^w���0A��a]�  �hZ3�T0 k� � ,�$,(%2't �8t B  �3    � �8�S�#�L.XOLL,,�K�� ^w���0A��b]�! �hZ3�T0 k� ,,� ,(%2't �8t B  ��?    � �8�T��L.TQLL,,�K�� ^{���0A��b]�! �hZ3�T0 k� ,,� ,(%2't �8t B ��?    � �8�V��L.PRLL0,�K�� ^{���0A��b]�! �hZ3�T0 k� ,,�,(%2't �8t B �?    � �8�W��L.PSR\4,�K�� ^{���1A��c]�" �hZ3�T0 k� ,,�,(%2't �8t B ��?    � �8�X��L.LTR\8,�K�� ^{���1A��c]�" �hZ3�T0 k� ,,�,(%2't �8t B ��?    � �8�Y��L.HUR\<,�K�� ^{���1A��d]�" �iZ3�T0 k� ,,�,(%2't �8t B ��?    � �8�Z��L.HVR\@+�O�� ^{�� 2A��d]�# �iZ3�T0 k� �,�,(%2't �8t B ��?    � �8�[��L.DWR\@+�O�� ^{�2A��e]�# �iZ3�T0 k� �,�,(%2't �8t B ��?    � �8�\�L.DXR\D+�O�� ^{�3A��e]�# �iZ3�T0 k� �-�-(%2't �8t B ��?    � �8�]�L.@YR\H+�O�� ^{�3A��e]�$ �iZ3�T0 k� �-�-(%2't �8t B ��?    � �8�^�L.<ZR\L+�O�� ^{�3A��f]�$ �iZ3�T0 k� �-�-(%2't �8t B ��?    � �8�_�L.<[RlP+�O�� ^{�4A��f]�$ �jZ3�T0 k� <-�-(%2't �8t B ��?    � �8�`�L.8\RlT+�O�� ^{�4A��g]�% �jZ3�T0 k� <-�-(%2't �8t B ��?    � �8�a�L.8]RlX+�S�� ^{�4A��g]�% �jZ3�T0 k� <-�-(%2't �8t B ��?    � �8�b��L.4^RlX*�S�� ^{� 5A��g]�% �jZ3�T0 k� <-�-(%2't �8t B ��?    � �8�c��L.4_Rl\*�S�� ^�$5A��h]�& �jZ3�T0 k� <-�-(%2't �8t B ��?    � �8�d��L.0`Rl`*�S�� ^�(5A��h]�& �jZ3�T0 k� �-�-(%2't �8t B ��?    � �8�e���L.0aRld*�S�� ^�(6A��h]�& �kZ3�T0 k� �-�-(%2't �8t B ��?    � �8�e���L.,bR|h*�S�� ^�,6A��i]�& �kZ3�T0 k� � .�.(%2't �8t B ��?    � �8�f���L.,cR|h*�S�� ^�06A��i]�' �kZ3�T0 k� � .�.(%2't �8t B ��?    � �8�g���L.(dR|l*�S�� ^�47A��i]�' �kZ3�T0 k� � .�.(%2't �8t B ��?    � �8�h���L.(eR|p*�W�� ^�87A��j]�' �kZ3�T0 k� +�.� .(%2't �8t B ��?    � �8�i���L.$fR|t*�W�� ^�<7A��j]�' �kZ3�T0 k� +�.� .(%2't �8t B ��?    � �8�j���L$fR|t*�W�� ^�@8A��j]�( �kZ3�T0 k� +�.��.(%2't �8t B ��?    � �8Mk���L gR|x)�W�� ^�@8A��k]�( �kZ3�T0 k� +�.��.(%2't �8t B ��?    � �8Mk���L hR||)�W�� ^�D8A��k]�( �lZ3�T0 k� +�.��.(%2't �8t B ��?    � �8Ml���LiR||)�W�� ^�H8A��k]�( �lZ3�T0 k� ��.��.(%2't �8t B ��?    � �8Mm���LjR|�)�W�� ^�L9A��l]�) �lZ3�T0 k� ��.��.(%2't �8t B ��?    � �8Mn���LjR|�)�W�� ^�P9A��l]�) �lZ3�T0 k� ��/��/(%2't �8t B ��?    � �8Mp���C�kR|�)�[�� ^� P9A��l]�) �lZ3�T0 k� ��/��/(%2't �8t B ��?    � �8	]q���C�lR|�)�[�� ^� T9A��l]�) �lZ3�T0 k� ��/��/(%2't �8t B ��?    � �8	]r���C�mR|�)�[�� ^� X:A��m]�* �lZ3�T0 k� K�/��/(%2't �8t B ��?   � �8	]r���C�mR|�)�[�� ^�� X:A��m]�* �lZ3�T0 k� K�/��/(%2't �8t B ��?    � �8	]s=��C�nR|�)�[�� ^�� \:A��m]�* �mZ3�T0 k� K�/��/(%2't �8t B ��?    � �8	]t=��C�oR|�)�[�� ^�� `;A��m]�* �mZ3�T0 k� K�/��/(%2't �8t B ��?    � �8	]u=��C�pR|�(�[�� ^�� d;A��n]�+ �mZ3�T0 k� K�/��/(%2't �8t B ��?    � �8	mv=��C�pR|�(�[�� ^�� d;A��n]�+ �mZ3�T0 k� ��/��/(%2't �8t B ��?    � �8	mu=��C� qR|�(�[�� ^�� h;A��n]�+ �mZ3�T0 k� ��/��/(%2't �8t B ��?    � �8	mu=��C��rR|�(�[�� ^�� l;A��o]�+ �mZ3�T0 k� ��0��0(%2't �8t B  ��?    � �8	mu=��C��rR|�(�[�� ^�� l<A��o]�+ �mZ3�T0 k� ��0��0(%2't �8t B  ��?    � �8	mu=��C��rR|�(�_�� ^�� p<A��o]�, �mZ3�T0 k� ��0��0(%2't �8t B  -�?    � �8u=��C��rR|�(�_�� ^�� p<A��o]�, �mZ3�T0 k� +�0��0(%2't �8t B  ��?    � �8t=��C��rR|�(�_�� ^�� t<A��o]�, �nZ3�T0 k� +�0��0(%2't �8t B  ��?    � �8tM��C��sR|�(�_�� ^�� x=A��o]�, �nZ3�T0 k� +�0��0(%2't �8t B  ��?    � �8tM��C��sR|�(�_�� ^�� x=A��o]�, �nZ3�T0 k� +�0��0(%2't �8t B  ��?    � �8tM��C��sR|�(�_�� ^�� |=A��o]�- �nZ3�T0 k� +�0��0(%2't �8t B  ��?    � �8� tM��E]�tR|�(�_�� ^�� |=A��o]�- �nZ3�T0 k� ��0��0(%2't �8t B ��?    � �8� tM��E]�uR|�(�_�� ^�� �=A��p]�- �nZ3�T0 k� ��0��0(%2't �8t B ��?    � �8��tͳ�E]�uR|�(�_�� ^�� �>A��p]�- �nZ3�T0 k� ��1��1(%2't �8t B ��?    � �8��tͯ�E]�vR|�( n_�� ^�� �>A��p]�- �nZ3�T0 k� ��1��1(%2't �8t B ��?    � �8��tͫ�E]�vR|�' nc�� ^�� �>A��p]�- �nZ3�T0 k� ��1��1(%2't �8t B ��?    � �8��tͧ�EM�vR|�' nc�� ^�� �>A��p]�. �nZ3�T0 k� ;�1��1(%2't �8t B ��?    � �8��tͤEM�vR|�' nc�� ^�� �>A��p]�. �nZ3�T0 k� ;�1��1(%2't �8t B ��?    � �8��t͠EM�vR|�' nc�� ^�� �?A��p]�. �oZ3�T0 k� ;�1��1(%2't �8t B ��?    � �8��s͜EM�vR|�'�c�� ^�� �?A��p]�. �oZ3�T0 k� ;�1��1(%2't �8t B ��?    � �8��s��C��vR|�'�g�� ^�� �?A��p]�. �oZ3�T0 k� ;�1��1(%2't �8t B  ��?    � �8��s��	C��vR|�'�g�� ^�� �?A��p]�/ �oZ3�T0 k� ��1��1(%2't �8t B  ��?    � �8��s��C��vR|�'�g�� ^�� �@A��p]�/ �oZ3�T0 k� ��2��2(%2't �8t B  ��?    � �8��r��C��vR|�'�g�� ^�� �@A��p]�/ �oZ3�T0 k� ��2��2(%2't �8t B  ��?    � �8��r��C��vR|�'�g�� ^�� �@A��o]�/ �oZ3�T0 k� ��2��2(%2't �8t B  ��?    � �8��q��C��vR|�'�g�� ^�� �@A��o]�/ �oZ3�T0 k� ��2��2(%2't �8t B  ��?    � �8��q�|C��vR|�'�g�� ^�� �@A��o]�/ �oZ3�T0 k� +�2��2(%2't �8t B  ��?    � �8��p�xC��vR|�'�g�� ^�� �@A��o]�/ �oZ3�T0 k� +�2��2(%2't �8t B  ��?    � �8��p�tC��vR|�'�g�� ^�� �AA��o]�0 �oZ3�T0 k� +�2��2(%2't �8t B  ��?    � �8��o�pC��vR|�'�g�� ^�� �AA��o]�0 �oZ3�T0 k� +�2��2(%2't �8t B  ��?    � �8��n�lC��vR|�'�g�� ^�� �AA��o]�0 �oZ3�T0 k� +�2��2(%2't �8t B  ��?    � �8��n�hC��vR|�'�c�� ^�� �AA�|o]�0 �oZ3�T0 k� ��2��2(%2't �8t B  ��?    � �8��m�dC��vR|�'�c�� ^�� �AA�|o]�0 �oZ3�T0 k� ��2��2(%2't �8t B  ��?    � �8��m�`C��vR|�&�c�� ^�� �AA�xn]�0 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��l�\!C��uR|�&�c�� ^�� �BA�tn]�0 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��l�X#C��uR|�&�_�� ^�� �BA�pn]�1 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��k�T$C��uR|�&�_�� ^�� �BA�ln]�1 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��k=P&C��uR|�&�\ � ^�� �BA�ln]�1 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��k=L(C��tR|�&�X� ^�� �BA�hn]�1 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��j=H*C��tR|�&�X� ^�� �BA�dm]�1 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��j=D,C��tR|�&�T� ^�� �BA�`m]�1 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��j=@.C��sR|�&�T� ^�� �BA�`m]�1 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��j=<0C��sR|�&�P� ^�� �CA�\m]�1 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��jM81C��sR|�&�P� ^�� �CA�Xm]�1 �oZ3�T0 k� ��3��3(%2't �8t B  ��?    � �8��iM43C��sR|�&�L� ^�� �CA�Tl]�2 �oZ3�T0 k� ��4��4(%2't �8t B  ��?    � �8��iM45C��rR|�&�L� ^�� �CA�Pl]�2 �oZ3�T0 k� ��4��4(%2't �8t B  ��?    � �8��hM07C��rR|�&�H	� ^�� �CA�Ll]�2 �oZ3�T0 k� ��4��4(%2't �8t B  ��?    � �8��hM,9C��qR|�&�D
� ^�� �CA�Hl]�2 �oZ3�T0 k� ��4��4(%2't �8t B  ��?    � �8��g	](:C��qR|�&�D� ^�� �CA�Hk]�2 �oZ3�T0 k� ��4��4(%2't �8t B  ��?    � �8��g	](<C��qR|�&�@� ^�� �CA�Dk]�2 �oZ3�T0 k� ��4��4(%2't �8t B  ��?    � �8��f	]$=C͈pR|�&�<� ^�� �DA�@k]�2 �oZ3�T0 k� ��4��4(%2't �8t B  ��?    � �8��f	]$?C̈́pR|�&�8� ^�� �DA�<k]�2 �oZ3�T0 k� ��4��4(%2't �8t B  ��?    � �8��e	] @C̀oR|�&�8� ^�� �DA�8j]�2 �oZ3�T0 k� ��4��4(%2't �8t B  ��?    � �8��d	m BC�|nR|�&�4� ^�� �DA�4j]�3 �oZ3�T0 k� ��4��4(%2't �8t B  ��?    � �8\�c	mCC�xnR|�&�0� ^�� �DA�0j]�3 �oZ3�T0 k� ��4��4(%2't �8t B  ��?   � �8\�c	mDE�tmR|�&�,� ^�� �DA�,i]�3 �oZ3�T0 k� ��5��5(%2't �8t B  ��?    � �8\�b	mEE�plR|�&�(� ^�� �DA�(i]�3 �oZ3�T0 k� ��5��5(%2't �8t B  ��?    � �8\�a	mFE�hlR|�&�$� ^�� �DA�$i]�3 �pZ3�T0 k� ��5��5(%2't �8t B  ��?    � �8\�`	]GE�dkR|�&� � ^�� �DA� i]�3 �pZ3�T0 k� ��5��5(%2't �8t B  ��?   � �8\�`	]HE�`jR|�&� � ^�� �EA� h]�3 �pZ3�T0 k� ��5��5(%2't �8t B  ��?    � �8\�_	]IE�`jR|�&�� ^�� �EA� h]�3 �pZ3�T0 k� ��5��5(%2't �8t B  ��?    � �8\�^	]JE�`jR|�&�� ^�� �EA� h]�3 �pb��T0 k� ��5��5(%2't �8t B  ��?    � �8\�]	]KE�`jR|�&�� ^�� �EA�h]�3 �pb��T0 k� ��5��5(%2't �8t B  ��?    � �8\�\�LE�\iR|�&�� ^�� �EA�h]�3 �pb��T0 k� ��5��5(%2't �8t B  ��?    � �8\�\�MC�XiR|�%�� ^�� �EA�h]�4 �pb��T0 k� ��5��5(%2't �8t B  ��?    � �8\�[�NC�TiR|�%� � ^�� �EA�h]�4 �pb��T0 k� ��5��5(%2't �8t B  ��?    � �8\�Z�OC�TiR|�%� "" ^�� �EA�h]�4 �pb��T0 k� ��6��6(%2't �8t B  ��?    � �8\�Y�OC�PiR|�%��#" ^�� �EA�h]�4 �pb��T0 k� ��6��6(%2't �8t B  ��?    � �8l�Y�PC�LhR|�%��%" ^�� �EA�g]�4 |pb��T0 k� ��6��6(%2't �8t B  ��?    � �8l�X�PK�HhR|�%��&" ^�� �FA� g]�4 |pb��T0 k� ��6��6(%2't �8t B  ��?    � �8l�W�QK�DgR|�%��'" ^�� �FA��g]�4 |pb��T0 k� ��6��6(%2't �8t B  ��?    � �8l�W�QK�@gR|�%��)" ^�� �FA��g]�4 |pb��T0 k� �|6��6(%2't �8t B  ��?    � �8l�V�RK�<fR|�%��*" ^�� �FA��g]�4 |pZ3�T0 k� �|6��6(%2't �8t B  ��?    � �8l�V�RK�8fR} %��," ^�� �FA��g]�4 |pZ3�T0 k� �|6��6(%2't �8t B  ��?    � �8l�V�SK�8fR} %��," ^�� �FA��g]�5 |pZ3�T0 k� �x6�|6(%2't �8t B  ��?    � �8l�V�TK�4eR} %��-" ^�� �FA��g]�5 xpZ3�T0 k� �x6�|6(%2't �8t B  ��?    � �8l�V�TK�0eR} %��." ^�� �EA��g]�6 xpZ3�T0 k� �x6�|6(%2't �8t B  ��?    � �8l�V�UK�0eR} %��/� ^�� �EA��g]�6 xpZ3�T0 k� �t6�x6(%2't �8t B  ��?    � �8l�V�UK�0fR} %��/� ^�� �EA��g]�7 xpZ3�T0 k� �t7�x7(%2't �8t B  ��?    � �8l�V�UK�,fR}%��0� ^�� �EA��f]�7 xpZ3�T0 k� �t7�x7(%2't �8t B  ��?    � �8l�U�UK�(fR}%��1� ^�� �EA��f]�7 xpZ3�T0 k� �p7�t7(%2't �8t B  ��?    � �8l�U�UK�(fR}%��2� ^�� �EA��f]�8 xpZ3�T0 k� �p7�t7(%2't �8t B  ��?    � �8l�U�UL$fR}%��3� ^�� �EA��f]�8 xpZ3�T0 k� �p7�t7(%2't �8t B  ��?   � �8l�U�UL$gR�%��4� ^�� �DA��f]�9 tpbs�T0 k� �l7�p7(%2't �8t B  ��?   � �8l�U�UL gR�%��5� ^�� �DA��f]�9 tpbs�T0 k� �l7�p7(%2't �8t B  ��?    � �8l�T�UL gR�%��6� ^�� �DA��f]�9 tpbs�T0 k� �p7�t7(%2't �8t B  ��?    � �8l�T�ULgR�%��7� ^�� �DA��f]�: tpbs�T0 k� �p7�t7(%2't �8t B  ��?    � �8l�T�ULgR�%��9� ^�� �DA��f]�: tpbs�T0 k� �p7�t7(%2't �8t B  ��?    � �8l�T�ULgR�%��9!� ^�� �DA��f]|; tpbs�T0 k� �p7�t7(%2't �8t B  ��?    � �8l�T�ULhR�%��:!� ^�� �DA��f]x; tpbs�T0 k� �p7�t7(%2't �8t B  ��?    � �8l�S�ULhR�%��;!� ^�� �DA��f]t; tpbs�T0 k� �p8�t8(%2't �8t B  ��?    � �8l�S �ULhR�%ݼ<!� ^�� �CA��f]t< tpbs�T0 k� �p8�t8(%2't �8t B  ��?    � �8l�S �ULhUm%ݸ=!� ^�� �CA��f]p< ppbs�T0 k� �p8�t8(%2't �8t B  ��?    � �8l�S �ULhUm%�?!� ^�� �CA��f]l= ppbs�T0 k� �p8�t8(%2't �8t B  ��?    � �8l�S �ULiUm%�@!� ^�� �CA��e]h= ppZ3�T0 k� �p8�t8(%2't �8t B  ��?    � �8l�S �ULiUm%�A!� ^�� �CA��e]h= ppZ3�T0 k� �p8�t8(%2't �8t B  ��?    � �8l�R �ULiUm%�B!� ^�� �CA��e]d> ppZ3�T0 k� �p8�t8(%2't �8t B  ��?    � �8l�RULiUm%�C!� ^�� �CA��e]`> ppZ3�T0 k� �p8�t8(%2't �8t B  ��?    � �8l�RULiUm%�D!� ^�� �CA��e]`> ppZ3�T0 k� �t8�x8(%2't �8t B  ��?    � �8l�RULiUm%�E� ^�� �CA��e]\? ppZ3�T0 k� �t8�x8(%2't �8t B  ��?    � �8l�RULiUm%�F� ^�� �BA��e]\? ppZ3�T0 k� �t8�x8(%2't �8t B  ��?    � �8l�RUL jA�%��F� ^�� �BA��e]X? ppZ3�T0 k� �t8�x8(%2't �8t B  ��?    � �8l�Q]UL jA�%��G� ^�� �BA��e]T? lpZ3�T0 k� �t8�x8(%2't �8t B  ��?    � �8l�Q]UL jA�%��H� ^�� �BA��e]P@ lpZ3�T0 k� �t9�x9(%2't �8t B  ��?    � �8l�Q]UL�jA�%��H� ^�� �BA��e]P@ lpZ3�T0 k� �t9�x9(%2't �8t B  ��?    � �8l�Q]UL�jA�%��I� ^�� �BA��e]L@ lpZ3�T0 k� �t9�x9(%2't �8t B  ��?    � �8l�Q]UL�jA�%��J� ^�� �BA��e]L@ lpZ3�T0 k� �t9�x9(%2't �8t B  ��?    � �8l�Q�UL�jA�%�|K� ^�� �BA��e]HA lpZ3�T0 k� �t9�x9(%2't �8t B  ��?    � �8l�Q�UL�kA�%�xL� ^�� �BA��e]DA lpZ3�T0 k� �t9�x9(%2't �8t B  ��?    � �8\�P�UL�kA�%�tM� ^�� �BA��d]DA lpZ3�T0 k� �t9�x9(%2't �8t B  ��?    � �8\�P�UL�kA�%�lN� ^�� �BA��d]@A lpZ3�T0 k� �t9�x9(%2't �8t B  ��?    � �8\�P�UL�kA�%�hN� ^�� �AA��d]<B hpZ3�T0 k� �x9�|9(%2't �8t B  ��?    � �8\�P�UL�kA�%hN� ^�� �AA��d]<B hpZ3�T0 k� �x9�|9(%2't �8t B  ��?    � �8\�P�UL�kA�%dO� ^�� �AA��d]<B hpZ3�T0 k� �x9�|9(%2't �8t B  ��?    � �8\�P�UL�kA�%`P� ^�� �AA��d]<B hqZ3�T0 k� �x9�|9(%2't �8t B  ��?    � �8��P�UL�lA�%`P� ^�� �AA��d]<B hqZ3�T0 k� �x9�|9(%2't �8t B  ��?    � �8��O�UL�lA�%\Q� ^�� �AA��d]<C hqZ3�T0 k� �x9�|9(%2't �8t B  ��?    � �8��O�UL�lA�%	�XR� ^�� �AA��c]<C hqZ3�T0 k� �x:�|:(%2't �8t B  ��?    � �8��O�UL�lA�%	�TR� ^�� �AA��c]8C dqZ3�T0 k� �x:�|:(%2't �8t B  ��?    � �8��N�UL�lA�%	�LS� ^�� �AA��c]8C dqZ3�T0 k� �x:�|:(%2't �8t B  ��?    � �8�N]UL�lA�%	�LS� ^�� �AA��c]8C dqZ3�T0 k� �x:�|:(%2't �8t B  ��?    � �8�M]UL�lA�%	�LT� ^�� �AA��c]8C dqZ3�T0 k� �x:�|:(%2't �8t B  ��?    � �8�M]UL�lA�%	�LT� ^�� �@A��c]8C dqZ3�T0 k� �x:�|:(%2't �8t B  ��?    � �8�L]UK��lA�%	�HT� ^�� �@A��c]4D dqZ3�T0 k� �x:�|:(%2't �8t B  ��?    � �8�L]UK��mA�%	�HU� ^�� �@A��c]4D dqZ3�T0 k� �|:��:(%2't �8t B  ��?    � �8�K]UK��mA�%	�HU� ^�� �@A��c]4D dqZ3�T0 k� �|:��:(%2't �8t B  ��?    � �8��K]UK��mA�%	�HU� ^�� �@A��c]4D `qZ3�T0 k� �|:��:(%2't �8t B  ��?    � �8��J] UK��mA�%�HU� ^�� �@A��b]4D `qZ3�T0 k� �|:��:(%2't �8t B  ��?    � �8��J] UK��mA�%�HU� ^�� �@A��b]4D `qZ3�T0 k� �|:��:(%2't �8t B  ��?   � �8��I] UC��mL=%�HU� ^�� �@A��b]4D `rZ3�T0 k� �|:��:(%2't �8t B  ��?   � �8��H] UC��mL=%�DU� ^�� �@A��b]0D `rZ3�T0 k� �|:��:(%2't �8t B  ��?    � �8]P��E��DM,	l���Xw,�C�����~lZ3�T0 k� �dy�hy(%2't �8t B  ��    � #�8]P��E��DM( l���Xy��C�����~lZ3�T0 k� �dy�hy(%2't �8t B  ��    � $�8]P��E}�DM$ l���X{��C�����~lZ3�T0 k� �dy�hy(%2't �8t B  ��    � %�8]P~�E}�DM  l���X}��C�����~hZ3�T0 k� �dz�hz(%2't �8t B  ��    � &�8]L~�E}�DM l���\��C�����~hZ3�T0 k� �d{�h{(%2't �8t B  ��    � '�8]L~#�E}�DM����\���C�����~d"Z3�T0 k� �d~�h~(%2't �8t B  ��    � (�8]H ~'�D��DM����\���C�����~d#Z3�T0 k� �h|�l|(%2't �8t B  ��    � )�8]H ~+�D��D]����`���C�����N`$Z3�T0 k� �h|�l|(%2't �8t B  ��    � *�8�H ~/�D��D]�����`���C�����N`&Z3�T0 k� �pw�tw(%2't �8t B  ��    � +�8�D!~7�D��!D] �����h���
C�����N\)Z3�T0 k� �xs�|s(%2't �8t B  ��    � ,�8�D!~;�I��"D\������h���C�����N\*Z3�T0 k� �|p��p(%2't �8t B  ��    � -�8�@"~?�I��$D\������l��C�����NX,Z3�T0 k� �|m��m(%2't �8t B  ��    � .�8]@"~C�I��&E������p~��C�����NX-Z3�T0 k� ��k��k(%2't �8t B  ��    � /�8]<"nG�I��'E������p~��C�����NX/Z3�T0 k� ��j��j(%2't �8t B  ��    � 0�8]<#nK�I��(E������t}��C�����NT1Z3�T0 k� ��h��h(%2't �8t B  ��    � 1�8]8#nS�I��+E��"���|||��C�����NT4Z3�T0 k� ��e��e(%2't �8t B  ��    � 2�8]8#nW�I� -El�#��|�{��C΄�� NP6Z3�T0 k� ��c��c(%2't �8t B  ��    � 3�8]8$n[�I�.El�$��|�z��C΀��^P7Z3�T0 k� ��b��b(%2't �8t B  ��    � 4�8]4$n[�I�/El�&��|�y��C�|��^P9Z3�T0 k� ��a��a(%2't �8t B  ��    � 5�8]4$n_�I�1El�'��|�x��C�x��^P;Z3�T0 k� ��`��`(%2't �8t B  ��    � 6�8]0%>c�E~3E\�)��|�v��C�l��^L?Z3�T0 k� ��^��^(%2't �8t B  ��    � 7�8]0%>c�E~5E\�+��|�t��C�h��	.L@Z3�T0 k� ��\��\(%2't �8t B  ��    � 8�8],%>g�E~6E\�,��|�s��C�d>�
.LBZ3�T0 k� ��[��[(%2't �8t B  ��    � 9�8],&>k�E~6E\�/  �|�q̼C�\>�.LFZ3�T0 k� ��X��X(%2't �8t B  ��    � :�8](&nk�E~7E\�0  �l�o̸C�T>�.LHZ3�T0 k� ��Y��Y(%2't �8t B  ��    � ;�8]('nk�E~9E\�1� �l�n̴C�P>�.LJZ3�T0 k� ��X��X(%2't �8t B  ��    � <�8]('no�E~:E\�2� �l�l̰C�L��.LLZ3�T0 k� ��X��X(%2't �8t B  ��    � <�8]$'no�E~>E\�5� �l�j̨"C�@
��.PPZ3�T0 k� ��V��V(%2't �8t B  ��    � <�8]$(no�I�?E\�6� �l�h̤$C�8	���PRZ3�T0 k� ��U��U(%2't �8t B  ��    � <�8]$(no�I�AE\�7� �l�g̜%C�4���PTZ3�T0 k� ��T��T(%2't �8t B  ��    � <�8] (no�I�BE\x8���l�eܘ'C�,���PVZ3�T0 k� �|R��R(%2't �8t B  ��    � <�8] (no�I�EE\l:���l�b܌*C� ���TZZ3�T0 k� �|O��O(%2't �8t B  ��    � <�8])no�I�GELd;���l�`܈,C���.X\Z3�T0 k� �|N��N(%2't �8t B  ��    � <�8])^o�I�HEL\<���l�_܄-C���.X^Z3�T0 k� �|L��L(%2't �8t B  ��    � <�8])^k�I�IELT=���l�]�|/C� ��.X`Z3�T0 k� �|J��J(%2't �8t B  ��    � <�8]*^k�I�LELD?��	�\�Z�p1C����.\dZ3�T0 k� ��N��N(%2't �8t B  ��    � <�8]*^k�I�MEL<@��
�\�X�h3C�����.`fZ3�T0 k� ��Q��Q(%2't �8t B  ��    � <�8]*^g�I�NEL4A���\�V�d4C�����.`hZ3�T0 k� ��S��S(%2't �8t B  ��    � <�8]*^g�I�OEL,A���\�U�\6C�����.djZ3�T0 k� ��T��T(%2't �8t B  ��    � <�8]+^c�I�QEL B����R�\6E�����hnZ3�T0 k� ��K��K(%2't �8t B  ��    � <�8]+�_�I�RELC����P�X7E�����hpZ3�T0 k� �|E��E(%2't �8t B  ��    � <�8]+�[�I�RELD����N�P8E�����lrZ3�T0 k� �|@��@(%2't �8t B  ��    � <�8]+�[�I�SELD����M�H9E�����lsZ3�T0 k� �x=�|=(%2't �8t B  ��    � <�8�,�S�I�UE;�F����I�<;E�����twZ3�T0 k� �t7�x7(%2't �8t B  ��    � <�8�,�O�I�VE;�F����G�4<Eݻ���xyZ3�T0 k� �t4�x4(%2't �8t B  ��    � <�8�,�K�I�VE;�F����E�,=Eݳ���x{Z3�T0 k� �p1�t1(%2't �8t B  ��    � <�8�,�G�I�WE;�G����D�$>C����||Z3�T0 k� �l/�p/(%2't �8t B  ��    � <�8�,�C�I�WE;�G����B�>C�����~Z3�T0 k� �l,�p,(%2't �8t B  ��    � <�8�,�;�I�XE;�G����>�?C������Z3�T0 k� �d(�h((%2't �8t B  ��    � <�8� ,�7�I�YE;�G����<�@C���|��Z3�T0 k� �`&�d&(%2't �8t B  ��    � <�8� ,�3�I�YE;�H	|����:��@I����x���Z3�T0 k� �h$�l$(%2't �8t B  ��    � <�8��+�/�I�ZE;�G	|���|8��AI����x���Z3�T0 k� �p"�t"(%2't �8t B  ��    � <�8��+�+�I�ZE;�G	|���|6��AI���t���Z3�T0 k� �t �x (%2't �8t B  ��    � <�8<�+�#�I�ZE;�G	|���x4��AI�{��t��Z3�T0 k� �x�|(%2't �8t B  ��    � <�8<�*��I�[E+�G	|���t2��AI�s��p��Z3�T0 k� �|��(%2't �8t B  ��    � <�8<�*^�I�[E+�G	|� ��t0��AI�o��p
��~Z3�T0 k� �|��(%2't �8t B  ��    � <�8<�*^�I�[E+�G	�� ��p.��BI�k��l	��}Z3�T0 k� �|��(%2't �8t B  ��    � <�8<�*^�I�[E+�F	�� ��l-��BI�c��l��}Z3�T0 k� �|��(%2't �8t B  ��    � <�8<�*^�I�[E+|F	��!��h)��BI�[��h��|Z3�T0 k� �t�x(%2't �8t B  ��    � <�8<�*]��I�[E+xE	��!��d'��BI�W��d~�{Z3�T0 k� �t�x(%2't �8t B  ��    � <�8<�*]��I�[E+pE	|�!�d%��BI�S��d~�zZ3�T0 k� �x�|(%2't �8t B  ��    � <�8<�*M�I�[E+lE	|�!�`#��AI�O��`~�yZ3�T0 k� ����(%2't �8t B  ��    � <�8<�*M�I�[E+hD	|�"�`!�AI�K��` ~�xZ3�T0 k� ����(%2't �8t B  ��    � <�8<�)MߊBN[E+hC	|�"�\�@I�G��_���wZ3�T0 k� ����(%2't �8t B  ��    � <�8L�)M׉BN[EhC%��"�\\�?I�C��[���vZ3�T0 k� �|	��	(%2't �8t B  ��    � <�8L�(MψBN[EdB%��#�\X�>I�?��[���uZ3�T0 k� �x�|(%2't �8t B  ��    � <�8L�(MˇBN[EdB%��#�\\�>I�;��W���tZ3�T0 k� �t�x(%2't �8t B  ��    � <�8L�'M��BN[EdB%��#�\\˨<I�7��S���rZ3�T0 k� �t�x(%2't �8t B  ��    � <�8��&M��@[U�dB%��$|'l\˨<E�3��S���qZ3�T0 k� �t�x(%2't �8t B  ��    � ;�8��&���@[U�dA%��$|'l`˨;E�/��S���pZ3�T0 k� �t�x(%2't �8t B  ��    � :�8��%���@[U�d@%��$|'l`˨;E�+��O���nZ3�T0 k� �{���(%2't �8t B  ��    � 9�8��%���@[U�d@%��$|'l`˨:E�'��O���mZ3�T0 k� �{���(%2't �8t B  ��    � 8�8��%���@[U�d?%��$|
'l`˨:E�#��K���lZ3�T0 k� �{���(%2't �8t B  ��    � 7�8��%���@n[U�h?%��%|	'|`
˨9E]��K���kZ3�T0 k� �{���(%2't �8t B  ��    � 6�8��$���@n[U�h>%�|%|'|d˨8E]��G��hZ3�T0 k� �����(%2't �8t B  ��    � 5�8��#M{�@n[U�h=%�x%| '|d˨8E]�	�G��gZ3�T0 k� �����(%2't �8t B  ��    � 4�8��#Ms�@n[U�h=%�x&| '|d˨7E]�	�C��eZ3�T0 k� �����(%2't �8t B  ��    � 3�8��"Mk�@n[U�h<%�t&| '|dˬ6EM�	�C��dZ3�T0 k� �����(%2't �8t B  ��    � 2�8��"Mc�@�[U�h<%�p&| '|hˬ6EM�	�C��cZ3�T0 k� �����(%2't �8t B  ��    � 1�8��!M[�@�[U�h;%�p&| '�k�ˬ5EL��	�C��aZ3�T0 k� ������(%2't �8t B  ��    � 0�8�� MS�@�[U�l;%�l&| '�k�ˬ5EL��	�C�`Z3�T0 k� ������(%2't �8t B  ��    � /�8��MC�@�[U�l:%�h'|#�'�k�ˬ4EL��	�?�]Z3�T0 k� ������(%2't �8t B  ��    � .�8��=?�CNZU�l9%�d'|#�'�o�ˬ3EL��	�?� [Z3�T0 k� ������(%2't �8t B  ��    � -�8��=7�CNZU�p9%�d'|#�'�o�˰3EL��	�?�$ZZ3�T0 k� ������(%2't �8t B  ��    � ,�8��=/�CNZU�p9%�`'|#�'�o�˰3EL��	�?�(XZ3�T0 k� ������(%2't �8t B  ��    � +�8��='�CNYU�p8%�`'|#�'�o�˰2E<��	�?�,VZ3�T0 k� ������(%2't �8t B  ��    � *�8��=�CNYU�p8%�\(|#�'�o�˰2E<��	�?�,UZ3�T0 k� ������(%2't �8t B  ��    � )�8�M�CNWU�p8%�X(|#�'|s�˰1E<��	�?�4QZ3�T0 k� ������(%2't �8t B  ��    � (�8�M�CNWU�p7%�T(�#�'|s�˴0E<��	�?�4PZ3�T0 k� ������(%2't �8t B  ��    � '�8�M�C^VU�p7�T(�#�'|s�˴0E<��	�?�o8NZ3�T0 k� ������(%2't �8t B  ��    � &�8�L��C^UU�p7�P(�#�'|s�˴/E<��	�?�o<LZ3�T0 k� ������(%2't �8t B  ��    � %�8�L��C^TU�t6�P)�#�'|s�˴/E<��	�?�o<JZ3�T0 k� ������(%2't �8t B  ��    � $�8�L�C^RU�t6�H)�#�'|w�˴.E<��	�?�o@GZ3�T0 k� ������(%2't �8t B  ��    � "�8܈L�C^QU�t5�D)�#�'lw�˴.E<��	�?�oDEZ3�T0 k� ������(%2't �8t B  ��    �  �8܈\ߊC^PU�t5�D)�#�'lw�˸-E<��	�?�oDCZ3�T0 k� ������(%2't �8t B  ��    � �8܈\׋C^OU�t4�@)�#�'lw�˸-E,��	�?�oHBZ3�T0 k� ������(%2't �8t B  ��    � �8܈\όC^NU�x4�<)�#�'lw�˸,E,��	�?�oH@Z3�T0 k� ������(%2't �8t B  ��    � �8܈	\ÍC^KU�x3�4)�#�'l{�˸,E,��	�?�oL<Z3�T0 k� ������(%2't �8t B  �� 
   � �8�\��CnJU�x3�0)�#�'l{�˸+E,���?�oL:Z3�T0 k� ������(%2't �8t B  �� 
   � �8�\��CnIU�x3�,)�#�{�˸+B����?�oL8Z3�T0 k� ������(%2't �8t B  �� 
   � �8�\��CnGU�x2�((�#�{�˼*B����?�_L7Z3�T0 k� ������(%2't �8t B  �� 
   � �8�\��CnFU�|2�((�#��˼*B���?�_L5Z3�T0 k� ������(%2't �8t B  �� 
   � �8�\��CnCU�|1� '�#��˼)B�{�C�_P1Z3�T0 k� ������(%2't �8t B  �� 
   � �8��l��CnAU�|1�'�#����)E�w�C�_L/Z3�T0 k� ������(%2't �8t B  �� 
   � �8��l��Cn@B�|1�&�#����(E�s�C�_L.Z3�T0 k� ������(%2't �8t B  �� 
   � �8��l��Cn>B�|1�&�#����(E�s�C�_L,Z3�T0 k� ������(%2't �8t B  �� 
   � �8��l��Cn;B��0�%�#����'E�k�G�_L)Z3�T0 k� ������(%2't �8t B  ��    � �8ܓ�l��C~9B��0$�#�����'E�k�G�_L'Z3�T0 k� ������(%2't �8t B  ��    � �8ܗ�l�C~7B��/$�#������&E�g�K�_H&Z3�T0 k� ������(%2't �8t B  ��    � �8ܗ�l�C~5B��/#�#������&E�c�K�_H$Z3�T0 k� ������(%2't �8t B  ��    � 
�8ܛ�l�C~3B��/#�#������%E�_�O�_H"Z3�T0 k� ������(%2't �8t B  ��    � �8ܟ�lw�C~/B��."�#������%CLW��S�ODZ3�T0 k� ������(%2't �8t B  ��    � �8ܟ�|w�C~-B��.!�#������%CLW��S�O@Z3�T0 k� ������(%2't �8t B  ��    � �8���|w�C~+B��. �#������$CLS��W�O@Z3�T0 k� ������(%2't �8t B  ��    � �8���|s�C~'B��.�#������$CLK��[�O<Z3�T0 k� ������(%2't �8t B  ��    � �8���|s�C~%B��.��#������$E,G��_��8Z3�T0 k� ������(%2't �8t B  ��    ����8���<s�CN"B��.��#������$E,C��c��8Z3�T0 k� ������(%2't �8t B  ��    ����8|��<o�CN B��.��#������#E,?��g��4Z3�T0 k� ������(%2't �8t B  ��    ����8|��<k�CNB��.��#������#E,;��o��0Z3�T0 k� ������(%2't �8t B  ��    ����8|��<k�CNB��.��#������#E,7��s��,Z3�T0 k� ������(%2't �8t B  ��    ����8|��<k�CNB��.��#������$E,7��w��(Z3�T0 k� ������(%2't �8t B  ��    ����8|��,k�CNB��.��#������$E3����(Z3�T0 k� ������(%2't �8t B  ��    ����8|��,k�CNB��.��#��߿�$E/����� Z3�T0 k� ������(%2't �8t B  ��    ����8|��,k�CNB˴.��#� |��$E+�����Z3�T0 k� �����(%2't �8t B  ��    ����8|��,g�CNB˴.��#� |��$E+�����Z3�T0 k� ����(%2't �8t B  ��    ����8|���g�E�	B˸/� �#� |��%E+�����Z3�T0 k� ����(%2't �8t B  ��    ����8|���g�E�B��/�$�#� |���%E'�����Z3�T0 k� ����(%2't �8t B  ��    ����9|���g�E�B��/�(�#����&E�'�����Z3�T0 k� ���#�(%2't �8t B  ��    ����:|���g�E� B��/�,
�#����&E�'�����Z3�T0 k� �'��+�(%2't �8t B  ��    ����;����k�E��B��/�,	�#����'E�'����OZ3�T0 k� �/��3�(%2't �8t B  ��    ����<����k�E��B��/�4�#��#��(E�'����N�
Z3�T0 k� �?��C�(%2't �8t B  ��&    ����=����k�E>�B��/�8�#��+��$(D�'��ÖN�
bs�T0 k� �G��K�(%2't �8t B  ��&    ����>����k�E>�B��/�8�#��/��()D�'��˕N�	bs�T0 k� �O��S�(%2't �8t B  ��&    ����?���o�E>�B��/�<�#��7��0)D�'��ϕN�	bs�T0 k� �S��W�(%2't �8t B  ��&    ����@���o�E>�B��/�G��#��G��8+D�+��۔N�	bs�T0 k� �W��[�(%2't �8t B  ��&    ����A���s�E>�B��/�G�#��O��@,D�+���N�bs�T0 k� �W��[�(%2't �8t B  ��&    ����B��s�E>�e /�K�#��W��D-D�+���>�bs�T0 k� �W��[�(%2't �8t B  ��&    ����C��w�E.�e/�O�#��_��H.D�/���>�bs�T0 k� �[��_�(%2't �8t B  ��&    ����D��{�E.�e/|W�#��k�<T/D�3����>�bs�T0 k� �c��g�(%2't �8t B  ��&    ����E��{�E.�e0|[�#��s�<X/D�3����>�bs�T0 k� �g��k�(%2't �8t B  ��&    ����F����E.�e0|_�#��{�<\0D�7���N�Z3�T0 k� �g��k�(%2't �8t B  �&    ����E�����E.#�e1|c�#��<d0D�7���N�Z3�T0 k� �c��g�(%2't �8t B  ��/    ����D�����E.#�e1|g�#���<h1D�;���N�	Z3�T0 k� �_��c�(%2't �8t B  ��O    ����C�����E.#�e$2o�#���<p2D�?���N�	Z3�T0 k� �[��_�(%2't �8t B ��O    ����B�����E.#�e(2s�|���<x2D�C���δ	Z3�T0 k� �W��[�(%2't �8t B ��O    ����A	����E.'�e,3w�|���<|2D�G��#�ΰ
Z3�T0 k� �W��[�(%2't �8t B ��O    ����@	����E.'�e03{�|���<�3D�G��'�Ψ
Z3�T0 k� �S��W�(%2't �8t B ��O    ����?	����E.'�e44��|���<�3D�K��+�Τ
Z3�T0 k� �S��W�(%2't �8t B ��O    ����>	����E+�e84��|���<�4D�O��/�ΠZ3�T0 k� �O��S�(%2't �8t B ��O    ����=	����E+�e,@5��|���<�4D�S��3�ΜZ3�T0 k� �K��O�(%2't �8t B ��O    ����<	����E/�e,H6��|#�÷<�5D�[��7�ސb��T0 k� �G��K�(%2't �8t B ��O    ����;	��,��E3�e,L6��|#�-˷<�6E�_��;�ތb��T0 k� �G��K�(%2't �8t B ��O    ����:	��,��E7�e,P6��|#�-Ϸ<�6E�c��?�ވb��T0 k� �@�D(%2't �8t B ��O    ����9	��,��E7�e,T7��|#�-׷<�6E�g��?�ހb��T0 k� �<�@(%2't �8t B ��O    ����8	��,��E;�e,X7���!�#�-۷<�7E�k��C��|b��T0 k� �<
�@
(%2't �8t B ��O    ����8	��,��E?�e,\8���!�#�-߷<�7E�o��C��tb��T0 k� �8�<(%2't �8t B ��O    ����8	��,��EC�e,`8���!�#�-�<�8E�s��G��pb��T0 k� �4�8(%2't �8t B ��O    ����8	��,ñEG�e,d8���!�#�-�<�8E�w��G��lb��T0 k� �4�8(%2't �8t B ��O    ����8	��,ǲEK�eh9���!�#�-�<�8E���G��db��T0 k� �0�4(%2't �8t B  ��O    ����8	��,ϳE�O�el9���!�  -��<�9E����K�N`b��T0 k� �0�4(%2't �8t B  ��O    ����8	��,׵E�W�et:���!� -��<�9E����K�NTZ3�T0 k� �(%�,%(%2't �8t B  /�O    ����8	��,۷E�[�ex:���!� .�<�:E|���K�NLZ3�T0 k� �()�,)(%2't �8t B  ��O    ����8	��,߸E�_�e|;���!� .�<�:E|���K�NDZ3�T0 k� �$,�(,(%2't �8t B  ��O    ����8	��,�E�c�e�;���!� .�<�:E|���K�N@Z3�T0 k� �$0�(0(%2't �8t B  ��O    ����8	��,�E�g�e�;���!� .�<�;E|���K�N8Z3�T0 k� � 4�$4(%2't �8t B  ��O    ����8	��,�E�o�e�<���!� .�<�;E|���K�N4Z3�T0 k� �8� 8(%2't �8t B  ��O    ����8	��,��E�s�e�<���!� .�<�;E|���K�N,Z3�T0 k� �<� <(%2't �8t B  ��O    ����8	��-�E��e,�=���� 	.'�<�<E|���K�N Z3�T0 k� �C�C(%2't �8t B  ��O    ����8	��-�E���e,�=��� 
.+�<�<E|���G��Z3�T0 k� �G�G(%2't �8t B  ��O    ����8	��-�E���e,�=��� 
./�<�=E|���G��Z3�T0 k� �K�K(%2't �8t B  ��O    ����8M�-�E~��e,�>��� �3�<�=D����C��Z3�T0 k� �N�N(%2't �8t B  ��G    ����8M��E~��e,�>��� �7�<�=D�û�C��Z3�T0 k� ��N� N(%2't �8t B  ��G    ����8M�#�E~��e,�?�#�� �?�<�>D�˾�?�M�Z3�T0 k� ��N� N(%2't �8t B  ��G    ����8M�+�E~��e,�?�+�� �C�<�>D����;�M�Z3�T0 k� ��O� O(%2't �8t B  ��G    ����8M�3�D���e,�?�/�� �G�<�?D����7�M�Z3�T0 k� ��O� O(%2't �8t B  ��G    ����8 �7�D���E��@�7�� �K���?D����3�M�Z3�T0 k� ��P��P(%2't �8t B  ��G    ����8 �?�D���E��@�?�� �O���?D����3�M�Z3�T0 k� ��R��R(%2't �8t B  ��G    ����8 �O�D���E��@�K�� �W�� @D���O+�M�Z3�T0 k� ��S� S(%2't �8t B  ��G    �  �8 �S�D���E��@ mO�� �[��AD���O'�M�Z3�T0 k� ��T��T(%2't �8t B  ��G    � �8 �[�D�×E��@ mW�� �[��AD���O#�M�Z3�T0 k� ��S��S(%2't �8t B  ��G    � �8 m�c�D�˗E��@ m[�� �_��BD���O�M� Z3�T0 k� ��S��S(%2't �8t B  ��G    � �8 m��k�D�ϖE��@ mc�� �c��CD���O�M�!Z3�T0 k� ��R��R(%2't �8t B  ��G    � �8 m��{�D�זE��@ mo�� �g��DD���O�=�#Z3�T0 k� ��S��S(%2't �8t B  ��G    � �8 m����D�ۗE��@ ms�� �g��ED�����=�$Z3�T0 k� ��S� S(%2't �8t B  ��G    � �8 m����D�ߗE��@ mw�� �k��FD�����=�%Z3�T0 k� ��P��P(%2't �8t B  ��G    � �8 �����D��E��? m�� �k��GD����=�&Z3�T0 k� ��N��N(%2't �8t B  ��G    � �8 �����D��E��? m��� �o��HD�����=�(Z3�T0 k� ��M��M(%2't �8t B  ��G    � 	�8 �����D��E��> m��� �o��ID�����=�*Z3�T0 k� ��K��K(%2't �8t B  ��G    � 
�8 �����D��E��> m��� �o��JD�����=x+Z3�T0 k� ��K��K(%2't �8t B  ��G    � �8M����D���E��= m��� �o��JD�����=t,Z3�T0 k� ��K��K(%2't �8t B  ��G    � �8M��ýD���E��= m��� �o��KD�����=l.Z3�T0 k� ��K��K(%2't �8t B  ��G    � �8M��ӽD��E��; m��� �o��LD�����=`0Z3�T0 k� ��F��F(%2't �8t B  ��G    � �8                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��er ]�#�#� � �� H�N   Y Y  	   ��+O<     It[�*�    ��              C Z�8�          �`�     ���  8	(          U��     
	  ��@X�     U���@w�      ��               !	 Z�8                 ���   @
"          m�7  9 9     �7]I     m���7�5    �r�#              S Z�8         ��   	  ���   
	'	           %/�  � �
  �Gmt     %0��GX    ��C              k Z�8          �P�     ���  8		           U��   > >      .�Q�|     U���R    ��k   	              Z�8          ��     ���  X

          �*  ��     B��;     �*��;                             ���?              �  ���    00            ����         V��v    ������t5                          �          �     ��@   0
           @MI         j�=�     @`��=#�    ���F                 ��C          (�     ��H   8�          b��        ~� ��     b�W� ��    ���               		 ^�b         �  �  ��B   (

           D�5         ��L��     D͇�M�    ���                    �         	 �      ��@   (
            r^           ���h     rm���     ��e                	    �         
  �0     ��@   P
B          ��
	      � ��{      ��{                              ���_              �  ��@    8	 1	                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          :��  ��        ���p�     :ި��^�                       x                j  �   �   �                          :    ��        ���       :  ��           "                                                �                         �+�@�7�G�Q����=� �L� �������  	  
             
  L    � �� �c�C       $ ``� � a�  a� Ƅ �c@ Ǆ  d@ �� d� �� d� �  d����< ����J ����X � �� \� �� 0\� �  ]  �D ]`���. ����< ����J ����X � ;� `o� <� p� <� p� <�  p� � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }`���� � �  b  �$ �e� �$ f� �D f� �d g  Є g  Ф g@ �D @w@ �� @w� �� @c@ �$ c� �D  c� �� d  �� 0d@ �  d� �D d� �� @[� �$ \@ �D  \` �� \� �� 0\� �  ]  �D ]` �d 0^@ �� 0^� �$ _  �D  _  ��  _` �� �r@ �� s@ �$  }` �d  }����� � 
�� W� 
�\ W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����8�� �� �  ������  
�fD
��L���"����D" � j  "  B   J jF�"     "�j  " ��
��
��"    B�j l �  B �
� �  �  
�  ,��  ��     ��  �    %��  ��     ��G       @    ��     ��=          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �?�      �� � �  ���        � �  ���        �        ��        �        ��        �     ��    � ) Rq        ��                         T�) ,  ���                                     �                 ����            0�� ���%��   �8��               89 Alexnder Mogilny                                                                                 1  1      �B �A �� �� � CB �
CC �" CI �
CJ �	c�R �
k~B k�R �B�( �KG � KO � K? �cj  �B�4 � B�< �K �K" � K$ � K% �K& �c�# � c�+ �C.4 � C4D pcV � � c^ � �"� � � "� � "� � �!*� �""� � #"�- �$� �%
�&&�} '�~8 (*DoP )*CwX **GX  *K_P  *RwH -*P_P .*OwX  *H_P 0*OwX  *H_X  *H_X  *K_ �4��8 5*DoP 6*CwX 7*GX  *K_X 9*H_X  *G8 ;*IoH <*P_X =*H_X  *GX  *K\                                                                                                                                                                                                                         �� R         �    @ 
        �     Z P E [  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    �sO�� ��������������������������������������������������������   �4, 8    ��@-@N��U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           >    &    ��  4�J      �                             ������������������������������������������������������                                                                                                                                      �  ��              �          ��               	 
     ������ ���������� �� �������������� ������ ���� ����� � �������  ���������������� ��� ������ ����������������������� ����������� ��������� ���� ������� �����������  ��� �������������������������� ������������������� ���                                 +    2    ��  L�J        	                           ������������������������������������������������������                                                                                                            
                            �    ��              �          ��                 	 	 ������������ � ��� � �������� ��� ����� ���������������������� � ������ ������������� ��������������� ���� ������������� ��������������������������� ������������������������������������������ �� ���������� �����������                                                                                                                                                                                                                                                                                                                             �             


             �   }�                     '�                       '�                 'v                         ������������  'r  '|����������������������������    ��������������������      ������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" ) J >                                 � #�} �`�                                                                                                                                                                                                                                                                                         	�)n�  "E        e                        m      e            m                                                                                                                                                                                                                                                                                                                                                                                                          0   >�  2�  2�  :#�  EZmp �̎�K��(����
�� �N D��� m���X����������        6  �� � : X
	         �   & AG� �   �              ���                                                                                                                                                                                                                                                                                                                                        N I   �     	                !�� !��                                                                                                                                                                                                                        Y   �� �� ����      �� e      ������ ���������� �� �������������� ������ ���� ����� � �������  ���������������� ��� ������ ����������������������� ����������� ��������� ���� ������� �����������  ��� �������������������������� ������������������� ��������������� � ��� � �������� ��� ����� ���������������������� � ������ ������������� ��������������� ���� ������������� ��������������������������� ������������������������������������������ �� ���������� �����������   ��      $����������������˪�������������������������������������f��ff��ff�������̺�ff�fffffffffffffffffff����ƹ��ffʻfff�fffjffffffffffff��������������������ʺ��l���f˪������������������������������������������������������������������fff�fff�fff�ffk�ffi�ff��ff��ff�ffffffff�fff�x�����w��xx�������wfffffff�ffff�fffww��ww�x����wx��fk��ff��ff��ffʹffj��fʪ�f�ˊ�k������������ʚ��������������������������������������������˫��ʫ��ff��fl��fl��ff̫fff�ffʬ�f���f�����������wu���w��l������f����W��������xww��Wy�l����x������k���W�fi���j���j���f����˘�����y�y�y����������������������������������������������������ʻ����ʫɚ�����l���ƨ�lƘ�j���k���̜i���j���kxx���wx������wx������������ƈx����������������wW����w�������������������������z����������˫��̺������������������������������������������������������������ʺ������k������������������������������������������x�j���˙�x�˘��̩�x������x���xx�x������x������wx���˫��ʫ����������˪�����ʻ��������������������������������������ʻ�ʻ�����ʪ̫����˺��������������������˪�����f���k��f��fǶW�g���k���̻���f������������������x�������˩f̺�����uw�����w��x�wXx��˪�����������l����l���i��ƹx�f�������������������ʫUW��UUU�UUUX      1      :   %�  :                       8     �  ����������      ��     8      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �t� � ���t� � �$ ^$    ���        ��   �   �    >     �f ��        p���� ��     �  �  $� >�������� J  $� �  �  $�   )   �   �    >������   �    v����     �  �� * ���2�������� Jk=   �  �� *       �  e� `� $ �� `� $ �$  �4 ��� �        �  ��   )�������2����   g���  �     f ^�         �� .       )      ��e����2�������J���`���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  "  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��  DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰ wwwywww�www�www�www�www�www�www����������!��������������������a��������݈����������a������������(-�a������!�-���www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�www�������������������������������������!�����!�-����������!-�����������!������www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�www������m����������݈����������������a݈�����m����!�����������a�-������www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�wwwy-��������!�����������������������������������!��������                                          �      �  a r!   f�"""""*��**"*�"�""�""v""*f   "  ""- ��"�"*"-""z"""""����            n   �  "  q  ��                          �  �                                 � gv"!g�vg�vggfvv|�b��r""gb"�vr�rgb��v���g���v���***�*q!q�"!a�!vwfqqr~� qw��q�~~q�����~~~�w~~w�w            �   ~   ��  ~~  �w      v    �                ggj�vvggvvgg!vg�g֪vvg�r�r��⢪rq**gjb�v�q*gjj*vv��gg�z�/�"!�"�*�""*z����qw�~q~ww��q~qwvq�w�`� ��� �w �~p w�p  ��                    �                        lggz�v��g        �       ggbvvrgggavvvqggav� �      ���w!z�w"""�!""*�"! ��        q� q�        `               �        �                      wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                               s   D   O   w   w   v   u   f   T   �   �              3@  DDp ��4 ��tp��wpO�tpdfwGfeTwfeWwfUFwdUFweTfp�DDp���p���@�w�p   C   D   O   D   w   u   U   U  F  d  f   f   D   �   �   �DD ���7���uP��e`O�V ffg ffG Ufw UU� FUN dFw ffp DDp ��p ��@ w�p  C4 4D@O�C���O�Dt�GVfeVfdFfdFfdUfffUfffwFff�DDD���� ���                    0   G   W   W   U   E   E   w   �   �   @    fg D� O�� �� w�}�w��}����������M���M���M��������y�                    �   �   �   �   �   �   �   �   ~   w       ���w���w���~���~�DMw�������������y�                        w���w}��wt��wt��w}M�����������   M   M   ~�  p�  p   p   p      �   �   �   �               vd  eVp ffpw�Op���w���G���M�}�                                     v   ub  ub  f   `   P               "  f  U` wfP        p   p   p   p   p   p   p   p                               C4 �y�                              f  vU`vf`D�O������p}�w�  ?�  ?�  ?�  33  3#                                      f  Ug���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            "! "   "      ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                              "! "   "      ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "! ""! " ""  "!  "! " ""            """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                              
      �  �  ��  �� �� �� 	�� D� EH EZ  DZ 4J 34Z3EH�T��ʄ
����ܩ���� ""�""�""�"/� �� �  ��� ̽� ��� �w� ��� ��� ��� ˻���ܚ��ة��ی����˻ݼˍ�ۻ���Ѕ" �" R�  B      ��  ��  �     �            � �� �   �       �   �   �"  "�  ���        �                                   ��.�  .                 ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                          ����     �   "  "     "   "   �                           ��   ��                  .  .  "  " ��                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��                      .   .   �        �  ��� ��� ��p �r`
wg`�ww   �   w  p  p  w   w  �  �   �  �                                                �                                ����                               ���                          ����                  �   �� �       �  �  "�  "   "              �  �                                                  ��	����ɪ�ܙ����ݼ "-� "� J.��#��C>Z�C U�D �Z�#�U"�C"�� ���                �  �˰ ̻� �wp �&  �vp �w� ɪ� ��� ��� �ۙ ��� �
� �" 0�" 0.�@ "�            ����˰ + �"  "" "  � �     .  .  "   "                   �   �   ��  �"" �""  ""   "                 �   ��   �                            � "�"                  .  ".  "               �                                           � ��                  �  �˰ ��� �wp �& ��� ���  �"  " ��"�""��"! � �  �   �   �   �                                                                                                            �w
���̩ۚ,���+��   �   �   �   �  �  9  D3  D2 T2 DB DB �@ ��  ��  ��  �  "" ""�"!��" ��       �                w�  ��� ��� ��� ˼����ɀ�؊�˽ـ��˰��̰�̻@"���"+H�"$X�"$�@"E� U� E� D� ,˸  ��  ��  ,� "" �"" """�"!���� � �              �         �           �       �                                      "  ."  �"    �          �� ̻� ��� ww� &'� vvw    �   �     �     �  �  "   "   "   "�  �                !��� �                                                                                                                                                                                          � 
��	�˽���w��rb��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            .  .     �   �           ��U %�P UX� ��  ��� ��� �̿ �/�""/�""/ ����    �            �/  ��  �                          �   � � /  �"" �"  �          �        �   �     �       �       "       .      �                    �"  �""� "�                   � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                                         �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �                      	   	   	   	�" �!  �  �� �   �                �  �� Ș ��  ��  �      �     �                                      � ����ݼ� ����                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��                        �          �   � � /  �"" �"  �    P � U  D  ���  ��  ̚  ��  
�  �"" �"" "/ �"����                  �             �   �     ���                            ��� ���  �"  " ��"�""��"! � �  �   �   �   �             ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                          �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �               0   0   �   �" �""��        "   "   "   �   �   ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �  �   �   �   �  �  �  �  �    ��                                 � "�"  �    � � �  ��  �   �    �          �         �                                                                                            �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���                          �    � .� .  �� 	  
  �  ",  ""  �"   "                      �"  �"  �          ��"� �"� ����            �   �   �   D   E�  U�  UO                         "  "  "                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��                        �          �   � � /  �"" �"  �                       �   �                      �".��".  ���    �                            � ��       "   "   "�  �                            �   ���                            �   "                                                                                                    �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �   �   �   ˰  ˙  ɪ  ��� ټ� �̰ �̰ ��� ��  ��                              ��                  �                        ��"� �"� ����          �   �   �   �  �  �  �  �                                                                                                                                                                                                          �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ����))������؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� ����"  �". �.  �                                        �� ��                  �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                          2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=LL����������D����3333DDDD    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����������A������ x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx""""�������I�I������ w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww""""�������I��D���I�������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(�D�M�D���M������3333DDDD �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""�����AMAD������ M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M""""������������������ � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�fFfFDfFFfFffdFffff3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DDFFDfFFfdFffff3333DDDD 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5""""wwwwwwwGGD x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x""""wwwwwwqwAqwAwA w w x y�������H���������������������������������H������yxww""""wwwwqwqAwAqAqAq  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(A�A�A�A��LD�����3333DDDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,�A�LDL�L�D�L�����3333DDDD +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+""""wwwwwwDGAD 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5""""wwwwqqDAAq =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=""""wwwwwwwGGwGGwGwGw     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( UQUUQUUQUUQUUUDUUUUU3333DDDD � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � �DEQQUUDUTEUUUU3333DDDD � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � �""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqB �A �� �� � CB �
CC �" CI �
CJ �	c�R �
k~B k�R �B�( �KG � KO � K? �cj  �B�4 � B�< �K �K" � K$ � K% �K& �c�# � c�+ �C.4 � C4D pcV � � c^ � �"� � � "� � "� � �!*� �""� � #"�- �$� �%
�&&�} '�~8 (*DoP )*CwX **GX  *K_P  *RwH -*P_P .*OwX  *H_P 0*OwX  *H_X  *H_X  *K_ �4��8 5*DoP 6*CwX 7*GX  *K_X 9*H_X  *G8 ;*IoH <*P_X =*H_X  *GX  *K\3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� � � � � � � � � � � � � � � � � � � � ����������������������������������������������������<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ���������������������������������������������������� � � � � � � � � � � � � � � � � � � � ���������������������������������������������������� � � � � � � � � � � � � � � � � � � � �����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3����������������������������������������� ��<�Z�K�\�K��<�S�O�Z�N� � � � � � � � � �-�2�3����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�2�3� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������,�-��.�/�0�1�2������������������������� �!�"�3�4�#�#�#�#�#�#�#�#�$������������������%�&�'�(�)�)�)�)�)�)�)�)�)�)�*�+������������������5�6���7�8�9�:�;�<�=�>�?�������������������� �!�"�#�#�#�#�#�#�#�@�4�#�$������������������%�A�B�C�D�E�F�G�H�I�J�K�L�M�N�O�����������������P�Q�R�S�T�U�V�W�X�Y�W�Z�[�\�]�^��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            