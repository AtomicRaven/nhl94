GST@�                                                           �`�                                                      �                    	      ���������	 J�������̸��X�������        �g      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"    B�j�
�  B ��
                                                                                 ����������������������������������      ��    bb= QQ0 4 111 44              		 

                     ��� �   � �                 nnE ))         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                ,i  �   O  �   @  #   �   �                                                                                '     )n)nE  �    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ���@�K� �� S� l�b|?�A�#�����0����3� T0 k� ��#;P e1�t B�1	�"q ��/    ����8���@�K� �� S� l�b|?�A�#������0����3� T0 k� ��#;P e1�t B�1	�"q ��/    ����8���@�K� �� S� l�b|?�Em#������0����3� T0 k� ��#;P e1�t B�1	�"q ��/    ����8���@�K� �� S� l�b|?�Em#������0����3� T0 k� ��#;P e1�t B�1	�"q ��/    ����8���@�K� �� S� l�b|?�Em#������0����3� T0 k� ��#[P e1�t B�1	�"q ��/    ����8���@�K� �� S� l�b|?�Em#������0����3� T0 k� ��#[P e1�t B�1	�"q ��/    ����8���@�K� �� S� l�Z<?�Em#������0����3� T0 k� ��#[P e1�t B�1	�"q ��/    ����8���@�K� �� S� l�Z<?�Em#������0����3� T0 k� ��#[P e1�t B�1	�"q ��/    ����8���@�O� �� S� l�Z<?�Em#������0����3� T0 k� ��#[P e1�t B�1	�"q ��/    ����8���@�O� �� S� l�Z<?�Em#������0����3� T0 k� ��#kP e1�t B�1	�"q ��/    ����8���@�O� �� S� l�Z<?�Em������0����3� T0 k� ��#kP e1�t B�1	�"q ��/    ����8���@�O� �� S� l�Z<?�Em������0����3� T0 k� ��#kP e1�t B�1	�"q ��/    ����8���@�O� �� S� l�Z<?�Em������0����3� T0 k� ��#kP e1�t B�1	�"q ��/    ����8���@�O� �� S� l�Z<?�Em������0����3� T0 k� ��#kP e1�t B�1	�"q ��/    ����8���@�O� �� S� l�Z<?�E]������0����3� T0 k� ��#{P e1�t B�1	�"q ��/    ����8���@�O� �� S� l�Z<?�E]�����0����3� T0 k� ��#{P e1�t B�1	�"q ��/    ����8���@�O� �� S� l�Z<?�E]�����0����3� T0 k� ��#{P e1�t B�1	�"q ��/    ����8���@�O� �� S� l�b�?�E]�����0����3� T0 k� ��#{P e1�t B�1	�"q ��/    ����8���@�O� �� S� l�b�?�E]�����0����3� T0 k� ��#{P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�b�?�C������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�b�?�C������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�b�?�C������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�b�?�C������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�b�?�C������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�b�?�C������0��]�3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�b�?�C������0��]�3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�b�?�C������0��]�3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�b�?�C������0��]�3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�Z<?�C������0��]�3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�Z<?�C������0��]�3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�Z<?�C������0��]�3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�S� �� S� l�Z<?�C������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�C������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�C������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�C������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�C������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A]�����0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A]�����0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A]�����0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A]�����0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A]�����0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A]�����0����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A]�����0����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A]�����0����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A]�����0����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A������0����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A������0����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�W� �� S� l�Z<?�A������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�[� �� S� l�Z<?�A������0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�[� �� S� l�Z<?�A������0���3� T0 k� ��$P e1�t B�1	�"q ��/    ����8���@�[� �� S� l�Z<?�A������0���3� T0 k� ��$P e1�t B�1	�"q ��/    ����8���@�[� �� S� l�Z<?�A������0���3� T0 k� ��$P e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A������0���3� T0 k� ��$P e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A������0���3� T0 k� ��$P e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A������/���3� T0 k� ��#;P e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A������/���3� T0 k� ��#;P e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A�������/���3� T0 k� ��#;P e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A�������/���3� T0 k� ��#;P e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A�������/���3� T0 k� ��#;P e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A�������/���3� T0 k� ��#KP e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A�������/���3� T0 k� ��#KP e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A�������/���3� T0 k� ��#KP e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A������/���3� T0 k� ��#KP e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A������/���3� T0 k� ��#KP e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A������/���3� T0 k� ��#kP e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A������/���3� T0 k� ��#kP e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A������/���3� T0 k� ��#kP e1�t B�1	�"q ��/    ����8���@�[� �� O� l�Z<?�A������/���3� T0 k� ��#kP e1�t B�1	�"q ��/    ����8���@�_� �� O� l�Z<?�A������/���3� T0 k� ��#kP e1�t B�1	�"q ��/    ����8���@�_� �� O� l�Z<?�A������/���3� T0 k� ��#{P e1�t B�1	�"q ��/    ����8���@�_� �� O� l�Z<?�A������/���3� T0 k� ��#{P e1�t B�1	�"q ��/    ����8��2A��� � O8# o;�Y| A�+��(2P<  ����#3� T0 k� �  � e1�t B�1	�"q  ��/    �   2��2A��� � O8# o;�a� A�+��(2P<  ����#"s� T0 k� �  � e1�t B�1	�"q  /�/    �   3��2A��� � O8# o;�a� A�+��(2P<  ����#"s� T0 k� ����e1�t B�1	�"q ��/    �   4��2A��� � O8# o;�a� A�+��(2P<  ����#"s� T0 k� ����e1�t B�1	�"q ��/    �   5��2A��� � O8# o;�a� A�+��(2P<  ����#"s� T0 k� ����e1�t B�1	�"q ��/    �   6��2A��� � O8# o;�a�  A�+��(2P<  ����#"s� T0 k� ����e1�t B�1	�"q ��/    �   7��2A��� � O8# o;�a�  A�+��(2P<  ����#"s� T0 k� ����e1�t B�1	�"q ��/    �   8��2A��� � O8# o;�a�  A�+��(2P<  ����#"s� T0 k� ����e1�t B�1	�"q ��/    �   9O�2D��� � �8# o;�a�$ D�+� (2P< P����#"s� T0 k� ����e1�t B�1	�"q ��/    �   :O�2D��� � �8" ;�Y|$ D�+� (2P< P����#3� T0 k� ���#�e1�t B�1	�"q ��/    �   ;O�2D��� � �8" ;�Y|$ D�+� (2P< P����"3� T0 k� ���#�e1�t B�1	�"q ��/    �   <O�2D��� � �8! ;�Y|$ D�+� (2P< P����"3� T0 k� �#��'�e1�t B�1	�"q ��/    �   =O�2D��� � �8! ;�Y|( D�+� (2P< P����"3� T0 k� �'��+�e1�t B�1	�"q ��/    ��� = �2D��� � �8  ;�Y|( D�+� `(2P< �����"3� T0 k� �'��+�e1�t B�1	�"q ��&    ��� = �2D��� � �8 O;�Y|( A�+� `(2P< �����"3� T0 k� �#��'�e1�t B�1	�"q ��&    ��� = �2E��� � �8O;�Y|( A�+� `(2P< �����!3� T0 k� ���#�e1�t B�1	�"q ��&    ��� = �2E��� � �8O;�Y|( A�+� `(2 < �����!3� T0 k� ���#�e1�t B�1	�"q ��&    ��� = �2E��� � �8O;�Y|( A�+� `(2 < ����� 3� T0 k� ���#�e1�t B�1	�"q ��&    ��� = o�2E��� � �8O;�Y|( A�+�@(2 < ����� 3� T0 k� ���#�e1�t B�1	�"q ��&    ��� = o�2E��� � �8�;�Y|( A�+�@(2 < �����3� T0 k� ���#�e1�t B�1	�"q ��&    ��� = o�2E�� � �8�;�a�( A�+�@(3 < �����"�� T0 k� ���#�e1�t B�1	�"q  ��&    ��� = o�2E�� � �8�;�a�( A�+�@(3 �< �����"�� T0 k� ���#�e1�t B�1	�"q  ��&    ��� = o�2E�� � �8�;�a�( A�+�@(3 �<����"�� T0 k� ���#�e1�t B�1	�"q  ��&    ��� =O�2E�� � �8�;�a�( A�/��(4 �<�� �"�� T0 k� ���#�e1�t B�1	�"q  ��&    ��� =O�2E�� � �8�;�a�( A�/��(4 �<�� �"�� T0 k� ���#�e1�t B�1	�"q  /�&    ��� <O�3Eo�� � �8�;�a�( A�/��(5 �<�� �"�� T0 k� ���#�e1�t B�1	�"q  ��&    ��� ;O�3Eo�� � �8�;�a�( A�/��(5@<�� �"�� T0 k� ���#�e1�t B�1	�"q  ��&    ��� :O�3Eo�� � �8�;�a�( A�/��(6@<�� �"�� T0 k� ���#�e1�t B�1	�"q  ��&    ��� 9O�4Eo�� � 8�;�a�( A�3��(6@<����"�� T0 k� �#��'�e1�t B�1	�"q  ��&    ��� 8O�4Eo�� � 8;�a�( A�3��(7@<����"�� T0 k� �#��'�e1�t B�1	�"q  ��&    ��� 7O�6E��� � 8;�a�( A�3��$8@<����"�� T0 k� �#��'�e1�t B�1	�"q  ��&    ��� 6O�6E��� � 8;�Y|( A�3��$9@<����3� T0 k� �#��'�e1�t B�1	�"q  ��&    ��� 5_�7E��� � 8;�Y|( A�3��$:@<����3� T0 k� �#��'�e1�t B�1	�"q  ��&    ��� 4_�8E��� � 8
o;�Y|( A�3��$;P<����3� T0 k� �#��'�e1�t B�1	�"q  ��&    ��� 3_�9E��� � 8	o;�Y|( A�7�� <P<����3� T0 k� �'��+�e1�t B�1	�"q  ��&    ��� 2_�:E��� � 8o;�Y|( A�7�� =P< ��p�3� T0 k� �'��+�e1�t B�1	�"q  ��&    ��� 1_�:E��� � 8o;�Y|( A�7�� >P< ��p�3� T0 k� �'��+�e1�t B�1	�"q  ��&    ��� 0_�<E��� � o8o;�Y|( A�7��@P<	 ��p�3� T0 k� �'��+�e1�t B�1	�"q  ��&    ��� ./�=E��� � o8 o7�Y|( A�7��AP<
 ��p�3� T0 k� �'��+�e1�t B�1	�"q  ��&    ��� ,/�?E��� � o;�_7�Y|( A�7��BP<
з�p�3� T0 k� �+��/�e1�t B�1	�"q  ��&    ��� */�@F�� � o;�_7�Y|( A�;��BP<
з�p�3� T0 k� �+��/�e1�t B�1	�"q  ��&    ��� )/�AF�� � o;�_3�Y|( A�;��CP<
з�p�3� T0 k� �+��/�e1�t B�1	�"q  ��&    ��� '/�BF�� � o7�_3�Y|( A�;��DP<
л�p�3� T0 k� �+��/�e1�t B�1	�"q  ��&    ��� %/�BF�� �o7�/�Y|( A�;��D`<
п�p�3� T0 k� �+��/�e1�t B�1	�"q  ��&    ��� #/�CF�� �o3�/�Y|( A�;��E`<
п�p�3� T0 k� �+��/�e1�t B�1	�"q  ��&    ��� !/�CE��� �o3�+�Y|( A�;��F`<���p�3� T0 k� �+��/�e1�t B�1	�"q  ��&    ��� /�DE��� �o/�+�Y|( A�;��H`<���p�3� T0 k� �/��3�e1�t B�1	�"q  ��&    ��� ��FE��� �_+�'�Y|( A�?��J`<���`�3� T0 k� �/��3�e1�t B�1	�"q  ��&    ��� ��HE��� �_'�'�Y|( A�?��L�<���`� 3� T0 k� �/��3�e1�t B�1	�"q  ��&    ��� ��IE�� �_'�'�Y|( A�?��M�<���`��3� T0 k� �/��3�e1�t B�1	�"q  ��&    ��� ��JE�� �_#�#�Y|( A�?��O�<���`��3� T0 k� �/��3�e1�t B�1	�"q  ��&    ��� ��JE�� �_��#�Y|( A�?��R�<���`��3� T0 k� �/��3�e1�t B�1	�"q  ��&    ��� ��LE�� �_���Y|( A�?��S�8 ���`��3� T0 k� �3��7�e1�t B�1	�"q  ��&    ��� ��MI��� �_���Y|( A�C��U�8!���`��3� T0 k� �3��7�e1�t B�1	�"q  ��&    ��� ��NI�� �_���Y|( A�C��V�8#���`��3� T0 k� �3��7�e1�t B�1	�"q  ��&    ��� ��PI�   �_���Y|( A�C��X�4$���`��3� T0 k� �3��7�e1�t B�1	�"q  ��&    ��� ��PI� �	_��Y|( A�C��[�4(���`��3� T0 k� �3��7�e1�t B�1	�"q  ��&    ��� 	�QI� �	^���Y|( A�C��]�0)���P��3� T0 k� �3��7�e1�t B�1	�"q  ��&    ��� �SI� �
N���Y|( A�C��^�0+���P��3� T0 k� �3��7�e1�t B�1	�"q  ��&    ��� �UI� �
N���Y|( A�C��`�,,���P��3� T0 k� �3��7�e1�t B�1	�"q  ��&    ��� �XI� �N���Y|( A�G��c�(0 ��P��3� T0 k� �7��;�e1�t B�1	�"q  ��&    ��� /�YI� �N��
�Y|( A�G�� d�$1 ��P��3� T0 k� �7��;�e1�t B�1	�"q  ��&    �����/�YI� ����
�Y|( A�G�� f� 3 ��P��3� T0 k� �7��;�e1�t B�1	�"q  ��&    �����/�ZI� ����
�Y|( A�G���g� 4 ��P��3� T0 k� �7��;�e1�t B�1	�"q  ��&    �����/�\I�	 ����
�Y|( A�G���i�6 ��P��3� T0 k� �7��;�e1�t B�1	�"q  ��&    �����/�]I�	 ����
��Y|( A�G���k�7 ��P��3� T0 k� �7��;�e1�t B�1	�"q  ��&    �����/�]I�
 ����
��Y|( A�G���n�: ��P��3� T0 k� �7��;�e1�t B�1	�"q  ��&    ������^I� ����
��Y|( A�G���p�< ��P��3� T0 k� �7��;�e1�t B�1	�"q  ��&    ������`I� ����
��Y|( A�G���q�= ��@��3� T0 k� �7��;�e1�t B�1	�"q  ��&    ������aI� ����
��Y|( A�G���s�> ��@��3� T0 k� �;��?�e1�t B�1	�"q  ��&    ������bI� ����
��Y|( A�K���t� @ ��@��3� T0 k� �;��?�e1�t B�1	�"q  ��&    ������dI� ����
��Y|( A�K���v��A ��@��3� T0 k� �;��?�e1�t B�1	�"q  ��&    ������eI� ����
.��Y|( A�K���x��B ��@��3� T0 k� �;��?�e1�t B�1	�"q  ��&    ������fI� ����
.ۿY|( A�K���y��C ��@��3� T0 k� �;��?�e1�t B�1	�"q  ��&    ������hI� ��{�
.ϾY|( A�K���|��E ��@��3� T0 k� �;��?�e1�t B�1	�"q  ��&    ������jI� ��s�
.˾Y|( A�K���}��F ��@��3� T0 k� �;��?�e1�t B�1	�"q  ��&    ������kI� ��k�
.ǽY|( A�K�����G ��@��3� T0 k� �;��?�e1�t B�1	�"q  ��&    �������lI� ��g�
.��Y|( A�K��̀��H ��@��3� T0 k� �;��?�e1�t B�1	�"q  ��&    �������mI� ��_�
.��Y|( A�K��Ȁ��I ��0��3� T0 k� �;��?�e1�t B�1	�"q  ��&    �������nI� ��W�
.��Y|( A�K��Ā��J ��0��3� T0 k� �;��?�e1�t B�1	�"q  ��&    �������oB@ ��O�
.��Y|( A�K�����K ��0��3� T0 k� �?��C�e1�t B�1	�"q  ��&    �������pB@ ��G�
.��Y|( A�O�߼��K ��0��3� T0 k� �?��C�e1�t B�1	�"q  ��&    �������qB@ ��?�
��Y|( A�O�ߴ��L ��0��3� T0 k� �?��C�e1�t B�1	�"q  ��&    �������qB@ ��7�
��Y|( A�O�߰~��L ��0��3� T0 k� �?��C�e1�t B�1	�"q  ��&    �������rB@ ��/�
��Y|( A�O�߬~��M ��0��3� T0 k� �?��C�e1�t B�1	�"q  ��&    �������s@ ��'�
��Y|( A�O��~��M ��0��3� T0 k� �?��C�e1�t B�1	�"q  ��&    �������s@ ���
��Y|( A�O��}��M �� ��3� T0 k� �?��C�e1�t B�1	�"q  ��&    �������t@ ���
��Y|( A�O��}��N0�� ��3� T0 k� �?��C�e1�t B�1	�"q  ��&    �������t@ ���
�Y|( A�O��|��N0�� ��3� T0 k� �?��C�e1�t B�1	�"q  ��&    �������u@ ���
{�Y|( A�O��|��N0�� ��3� T0 k� �?��C�e1�t B�1	�"q  ��&    ������u@` ����
k�Y|( A�O��{��N0�� ��3� T0 k� �?��C�e1�t B�1	�"q  ��&    ������v@` ����
g�Y|( A�O��|z��N0�� ��3� T0 k� �?��C�e1�t B�1	�"q  ��&    ������v@` ����
>_�Y|( A�O��tz��N ����3� T0 k� �?��C�e1�t B�1	�"q  ��&    ������v@` ����
>W�Y|( A�O��py��N ����3� T0 k� �C��G�e1�t B�1	�"q  ��&    ������v@` ����
>O�Y|( A�O�?hx��N ����3� T0 k� �C��G�e1�t B�1	�"q  ��&    ������vE� ����
>K�Y|( A�S�?`w�|M ����3� T0 k� �C��G�e1�t B�1	�"q  ��&    ������vE�
 ����
>C�Y|( A�S�?\w�xM ����3� T0 k� �C��G�e1�t B�1	�"q  ��&    ������ vE�
 �ͻ�
>;�Y|( A�S�?Tv�tM
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    ������(vE�	 �ͳ�
>3�Y|( A�S�?Pu�pL
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����p,vE� �ͫ�
>+�Y|( A�S�	�Hu�lL
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����p0vE  �ͣ�
>#�Y|( A�S�	�Dt�hK
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����p8vE  �͓�
>�Y|( A�S�	�8s�`J
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����p<uE   �M��
�Y|( A�S�	�4s�\J
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����pDuE $ �M��
�Y|( A�S�	�0r�XI
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����pHtE $ �M{�
��Y|( A�S�	�(r�XH
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����pLtE ( �Ms�
��Y|( A�S�	�$q�TH
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����pPsE , �Mk�
�Y|( A�S�	� q�PG
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����pTsE, �Mc�
�Y|( A�S�	�q�LF
������3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����pXrE0  �M[�
�Y|( A�S��p�HE
�����3� T0 k� �C��G�e1�t B�1	�"q  ��&    �����p\qE4  �MS�
ۯY|( A�S��p�DD
�����3� T0 k� �G��K�e1�t B�1	�"q  ��&    �����``qE7� �MK�
ӯY|( A�S��p�@C
�����3� T0 k� �G��K�e1�t B�1	�"q  ��&    �����`dpE;� �MC�
˯Y|( A�S��o�@B
�����3� T0 k� �G��K�e1�t B�1	�"q  ��&    �����`lnE?� �=3�
��Y|( A�W��n�8@
�����3� T0 k� �G��K�e1�t B�1	�"q  �&    �����`lmE?� �=+����Y|( A�W�� n�4?
�� ��3� T0 k� �G��K�e1�t B�1	�"q  �&    ������plE?� �=#����Y|( A�W���n�0>
�� ��3� T0 k� �G��K�e1�t B�1	�"q  ��&    ������tkE?� �=����Y|( A�W���m�0=
�� ��3� T0 k� �G��K�e1�t B�1	�"q  ��&    ������xjEC� �=����Y|( A�W���m�,<
�� ��3� T0 k� �G��K�e1�t B�1	�"q  ��&    ������|iE�C� �=����Y|( A�W���l�(;
�� ��3� T0 k� �G��K�e1�t B�1	�"q  ��&    ������|hE�G� �=����Y|( A�[���l�$:
�#� ��3� T0 k� �K��O�e1�t B�1	�"q  ��&   �������gE�G� �<�����Y|( A�[���l�$9
�'� ��3� T0 k� �K��O�e1�t B�1	�"q  ��&    �������fE�K� �<�����Y|( A�[���k� 8
�'� ��3� T0 k� �K��O�e1�t B�1	�"q  ��&    �������dE�K� �<�����Y|( A�[���k�7
�+� ��3� T0 k� �K��O�e1�t B�1	�"q  $�&    �������cE�O� �,�����Y|( A�[���j�6
�/� ��3� T0 k�  O��S�e1�t B�1	�"q  ��&   �������bE�O� �,����Y|( A�_���j�5
�/� ��3� T0 k�  O��S�e1�t B�1	�"q  ��&    �������`E�O� �,���{�Y|( A�_���j�4
�3� ��3� T0 k�  O��S�e1�t B�1	�"q  ��&    �������_E�O� �,���w�Y|( A�_���i�3
�7� ��3� T0 k�  O��S�e1�t B�1	�"q  ��&    �������]E�S� �,� �s�Y|( A�_���i�2
�7� ��3� T0 k�  S��W�e1�t B�1	�"q  ��&    �������\E�S� �,��o�Y|( A�_���i�2
�;� ��3� T0 k� �S��W�e1�t B�1	�"q  ��&   �������ZE�S� �,��k�Y|( A�c���h�1
�?� ��3� T0 k� �S��W�e1�t B�1	�"q  ��&    �������XE�S� �,��g�Y|( A�c���h�0
�?� ��3� T0 k� �S��W�e1�t B�1	�"q  ��&    �������WE�S� �,��g�Y|( A�c���h�/
�C� ��3� T0 k� �W��[�e1�t B�1	�"q  ��&   �������UE�S� �,��c�Y|( A�c���g�.
�C� ��3� T0 k� �W��[�e1�t B�1	�"q  ��&    �������SE�W� �,�	�c�Y|( A�g���g� -
�G� ��3� T0 k� �W��[�e1�t B�1	�"q  ��&    �������RC�W� ����_�Y|( A�g���g� -
�G� ��3� T0 k� �W��[�e1�t B�1	�"q  ��&    �������PC�S� ����_�Y|( A�g���f��,
�K� ��3� T0 k� �W��[�e1�t B�1	�"q  ��&    �������NC�S� ����[�Y|( A�g���f��+
�O� ��3� T0 k� �[��_�e1�t B�1	�"q  ��&    �������LC�S� ����[�Y|( A�g���f��*
�O� ��3� T0 k� �[��_�e1�t B�1	�"q  ��&    �������JC�S� ����[�Y|( A�k���e��*
�S� ��3� T0 k� �[��_�e1�t B�1	�"q  ��&    �������IC�S� ����W�Y|( A�k���e��)
�S� ��3� T0 k� �[��_�e1�t B�1	�"q  ��&    �������GC�O� ����W�Y|( A�k���e��(
�W� ��3� T0 k� �[��_�e1�t B�1	�"q  ��&    �����`�EK�O� |���W�Y|( A�k���d��(
�W� ��3� T0 k� �_��c�e1�t B�1	�"q  ��&    �����`�CK�O� |���W�Y|( A�k���d��'
�[� ��3� T0 k� �_��c�e1�t B�1	�"q  ��&    �����`�AK�O� |���W�Y|( A�o���d��&
�[� ��3� T0 k� �_��c�e1�t B�1	�"q  �&    �����`�?K�K� |���W�Y|( A�o���d��&
�_� ��3� T0 k�  c��g�e1�t B�1	�"q  ��/    �����`�=K�K� |���W�Y|( A�o���c��%
�_� ��3� T0 k�  g��k�e1�t B�1	�"q ��/    �����`�;K�K� |���W�Y|( A�o���c��$
�c� ��3� T0 k�  k��o�e1�t B�1	�"q ��/    �����0�9K�K� |���W�Y|( A�o���c��$
�c� ��3� T0 k�  o��s�e1�t B�1	�"q ��/    �����0�7K�G� |̀�[�Y|( A�s���c��#
�c� ��3� T0 k�  s��w�e1�t B�1	�"q ��/    �����0�5K�G� |�| �[�Y|( A�s���b��#
�g� ��3� T0 k�  w��{�e1�t B�1	�"q ��/    �����0�3K�G� |�|!�[�Y|( A�s���b��"
�g� ��3� T0 k� �{���e1�t B�1	�"q ��/    �����0�1K�G� |�x"�[�Y|( A�s���b��!
�k� ��3� T0 k� �����e1�t B�1	�"q ��/   �����0�/K�G� |�t$�_�Y|( A�s���b��!
�k� ��3� T0 k� ������e1�t B�1	�"q ��/    �����0�-K�C� |�p%�_�Y|( A�w��|a�� 
�o� ��3� T0 k� ������e1�t B�1	�"q ��/    �����0�+K�C� | �p&�c�Y|( A�w��|a�� 
�o� ��3� T0 k� ������e1�t B�1	�"q ��/    �����0�)L C� | �l'�c�Y|( A�w��xa��
�o� ��3� T0 k� 0�����e1�t B�1	�"q ��/    �����0�'L C� | �h(�g�Y|( A�w��xa��
�s� ��3� T0 k� 0�����e1�t B�1	�"q ��/    �����0�%L C� | �h)�g�Y|( A�w��ta��
�s� ��3� T0 k� 0�����e1�t B�1	�"q ��/    �����0�#L ?� | �d*�k�Y|( A�w��t`��
�w� ��3� T0 k� 0�����e1�t B�1	�"q ��/    �����@� L ?� | �`+�k�Y|( A�{��p`��
�w� ��3� T0 k� 0�����e1�t B�1	�"q ��/    �����@�L ?� | �`,�o�Y|( A�{��l`��
�w� ��3� T0 k� ������e1�t B�1	�"q ��/    �����@�L ?� x �\.�s�Y|( A�{��l`��
�{� ��3� T0 k� ������e1�t B�1	�"q ��/    �����@�L ?� x �X/�w�Y|( A�{��h_��
�{� ��3� T0 k� ������e1�t B�1	�"q ��/    �����@�L ;� x �X0�w�Y|( A�{��h_��
�{� ��3� T0 k� ������e1�t B�1	�"q ��/    �����@�L ;� x �T1�{�Y|( A�{��d_��
�� ��3� T0 k� ������e1�t B�1	�"q ��/    �����@�L ;� x!�T2��Y|( A�{��d_��
�� ��3� T0 k�  � �� e1�t B�1	�"q ��/    �����@�L ;� x!�P2���Y|( A���`_��
�� ��3� T0 k�  � �� e1�t B�1	�"q ��/    �����@�L ;� x!�L3���Y|( A���`_��
у� ��3� T0 k�  ���e1�t B�1	�"q ��/    �����@�L 7� x!�L4���Y|( A���\^��
у� ��3� T0 k�  ���e1�t B�1	�"q ��/    �����@�L 7� x!�H5���Y|( A���\^��
у� ��3� T0 k�  ���e1�t B�1	�"q ��/    �����P�
L 7� x!�H6���Y|( A���\^��
ч� ��3� T0 k� ����e1�t B�1	�"q ��/    �����P�L 7��x!�D7���Y|( A���X^��
ч� ��3� T0 k� ����e1�t B�1	�"q ��/    �����P�L 7��x!�D8���Y|( A���X^��
ч� ��3� T0 k� ����e1�t B�1	�"q ��/    �����P�L 7��x!�@9���Y|( A����T]��
ы� ��3� T0 k� ����e1�t B�1	�"q ��/    �����P�L 7��x!�@:���Y|( A����T]��
ы� ��3� T0 k� ����e1�t B�1	�"q ��/    �����P��L 3��x!�<;���Y|( A����P]��
ы� ��3� T0 k� @���e1�t B�1	�"q ��/    �����P��L 3��x!�<;���Y|( A����P]��
я� ��3� T0 k� @�	��	e1�t B�1	�"q ��/    �����P��L 3��x!�8<���Y|( A����P]��
я� ��3� T0 k� @�
��
e1�t B�1	�"q ��/    �����P��L 3��x!�8=���Y|( A����L]��
я� ��3� T0 k� @���e1�t B�1	�"q ��/    �����P�L 3��x"�4>���Y|( A����L]��
я� ��3� T0 k� @���e1�t B�1	�"q ��/    �����P{�L 3��x"�4?���Y|( A����H\��
ѓ� ��3� T0 k� ����e1�t B�1	�"q ��/    �����`w�L 3��x"�0?�ǢY|( A����H\��
ѓ� ��3� T0 k� ����e1�t B�1	�"q ��/    �����`w�L /��x"�0@�ˢY|( A����H\��
ѓ� ��3� T0 k� ����e1�t B�1	�"q ��/    �����`s�L /��x"�,A�ӢY|( A����D\��
ї� ��3� T0 k� ��� e1�t B�1	�"q ��/    �����`o�L /��x"�,B�עY|( A����D\��
ї� ��3� T0 k� � �e1�t B�1	�"q ��/    �����`k�L /��x"�(B�ۢY|( A����D\��
ї� ��3� T0 k� !�e1�t B�1	�"q ��/    �����`g�L /��x"�(C��Y|( A����@\��
ї� ��3� T0 k� !�e1�t B�1	�"q ��/    �����`c�L /��x"�(D��Y|( A����@[��
ћ� ��3� T0 k� !�e1�t B�1	�"q ��/    �����`_�L /��x"�$D��Y|( A����<[��
ћ� ��3� T0 k� !�e1�t B�1	�"q ��/   �����`_�L +��x"�$E��Y|( A����<[��
ћ� �3� T0 k� !�e1�t B�1	�"q ��/    �����`_�L '��x"� F���Y|( A����<[��
ћ� �3� T0 k� ��e1�t B�1	�"q ��/   �����`_�L '��t"� F���Y|( A����8[��
џ� �3� T0 k� �� e1�t B�1	�"q ��/    �����0[�L #��t"� G��Y|( A����8[��
џ� �3� T0 k� � �$e1�t B�1	�"q  ��/    �����0[�L ��t"�H��Y|( A����8[��
џ� �3� T0 k� �$�(e1�t B�1	�"q  -�/    �����0[�L ��t"�H��Y|( A����8[��
џ� �3� T0 k� �(�,e1�t B�1	�"q  ��/    �����0W�L ��t#I��Y|( A����4Z��
џ� �3� T0 k� 1,�0e1�t B�1	�"q  ��/    �����0W�K���t#I��Y|( A����4Z��
ѣ� �3� T0 k� 10�4e1�t B�1	�"q  ��/    �����0S�K���t#J�'�Y|( A����4Z��
ѣ� �3� T0 k� 14�8e1�t B�1	�"q ��/    �����0O�K���t#K�/�Y|( A����0Z��
ѣ� �3� T0 k� 18�<e1�t B�1	�"q ��/    �����0O�K���t#K�7�Y|( A����0Z��
ѣ� �3� T0 k� 1<�@e1�t B�1	�"q ��/    �����0O�K���t#L�;�Y|( A����0Z��
ѣ� �3� T0 k� �@�De1�t B�1	�"q ��/    �����0O�K���t#�L�C�Y|( A����,Z��
ѧ� �3� T0 k� �D�He1�t B�1	�"q ��/    �����0K�C���t#�M�K�Y|( A����,Z��
ѧ� �3� T0 k� �H�Le1�t B�1	�"q ��/    �����0G�C���t#�M�S�Y|( A����,Z��
ѧ� �3� T0 k� �L �P e1�t B�1	�"q ��/    �����@G�C���t#�M�[�Y|( A����,Y��
ѧ� �3� T0 k� �P!�T!e1�t B�1	�"q ��/    �����@C�C����t#�N�_�Y|( A����(Y��
ѧ� �3� T0 k� !T!�X!e1�t B�1	�"q ��/    �����@?�C����t#�N�g�Y|( A����(Y��
ѫ� �3� T0 k� !X"�\"e1�t B�1	�"q ��/    �����@?�C����t#�N�o�Y|( A����(Y��
ѫ� �3� T0 k� !\#�`#e1�t B�1	�"q ��/    �����@;�C����t#� N�w�Y|( A����(Y��
ѫ� �3� T0 k� !`$�d$e1�t B�1	�"q ��/    �����@7�C����t#� O��Y|( A����$Y��
ѫ� �3� T0 k� !d%�h%e1�t B�1	�"q ��/    �����@3�EO���t#� O���Y|( A����$Y��
ѫ� �3� T0 k� �h&�l&e1�t B�1	�"q ��/    �����@/�EO���t#�$O���Y|( A����$Y��
ѯ� �3� T0 k� �l&�p&e1�t B�1	�"q ��/    �����@/�EO���t#�$O���Y|( A����$Y��
ѯ� �3� T0 k� �p'�t'e1�t B�1	�"q ��/    �����@+�EO���t#�(O���Y|( A���� Y��

ѯ� �3� T0 k� �t(�x(e1�t B�1	�"q  ��/    �����@'�EO���t#�(O���Y|( A��� Y��

ѯ� �3� T0 k� �x)�|)e1�t B�1	�"q  ��/    �����P#�E?׿�t#�,N���Y|( A��� X��

ѯ� �3� T0 k� A|*��*e1�t B�1	�"q  ��/    �����P�E?Ӿ�t$�0N���Y|( A��� X��

ѯ� �3� T0 k� A�+��+e1�t B�1	�"q  ��/    �����P�E?ϼ�t$�0N���Y|( A��� X��

ѳ� �3� T0 k� A�+��+e1�t B�1	�"q  /�/    �����P�E?˻�t$�4N���Y|( A���X��	
ѳ� �3� T0 k� A�,��,e1�t B�1	�"q  ��/    �����P�E?˹�t$�8M�àY|( A���X��	
ѳ� �3� T0 k� A�-��-e1�t B�1	�"q  ��/    �����P�COǸ�t$�<M�ˠY|( A���X��	
ѳ� �3� T0 k� �.��.e1�t B�1	�"q  ��/    �����0�COö�t$�<M�ӠY|( A���X��	
ѳ� �3� T0 k� �/��/e1�t B�1	�"q  ��/    �����0�CO���t$�@L�נY|( A���X��	
ѳ� �3� T0 k� �0��0e1�t B�1	�"q  ��/    �����0�CO���t$�DL�ߠY|( A���X��	
ѳ� �3� T0 k� �0��0e1�t B�1	�"q  ��/    �����0�CO���t$�HK��Y|( A���X��
ѷ� �3� T0 k� �1��1e1�t B�1	�"q  ��/    �����0�I_���t$�LK��Y|( A���X��
ѷ� �3� T0 k� �2��2e1�t B�1	�"q  ��/    �����?��I_���t$�PJ��Y|( A���X��
ѷ� �3� T0 k� �3��3e1�t B�1	�"q  ��/    �����?��I_���t$�TJ���Y|( A���X��
ѷ� �3� T0 k� �4��4e1�t B�1	�"q  ��/    �����?��I_���t$�XI���Y|( A���W��
ѷ� �3� T0 k� �4��4e1�t B�1	�"q  ��/    �����?�I_���t$�\H���Y|( A���W��
ѷ� �3� T0 k� �5��5e1�t B�1	�"q  ��/    �����?�Io���t$�`H��Y|( A���W��
ѷ� �3� T0 k� �6��6e1�t B�1	�"q  ��/    �����?�Io���t$�dG��Y|( A���W��
ѷ� �3� T0 k� �7��7e1�t B�1	�"q  ��/    �����?�Io�� t$�hF��Y|( A���W��
ѻ� �3� T0 k� ��8��8e1�t B�1	�"q  ��/    �����?�Io�� t$�lE��Y|( A���W��
ѻ� �3� T0 k� ��9��9e1�t B�1	�"q  ��/    �����?�Io�� t$�tD��Y|( A���W��
ѻ� �3� T0 k� ��9��9e1�t B�1	�"q  ��/    �����O�I_�� t$�xD��Y|( A���W��
ѻ� �3� T0 k� ��:��:e1�t B�1	�"q  ��/    �����O�I_�� t$�|C�'�Y|( A���W��
ѻ� �3� T0 k� ��;��;e1�t B�1	�"q  ��/    �����OߢI_�� t$��B�+�Y|( A���W��
ѻ� �3� T0 k� ��<��<e1�t B�1	�"q  ��/    �����O۠I_�� t$��A�/�Y|( A���W��
ѻ� �3� T0 k� ��=��=e1�t B�1	�"q  ��/    �����O۟I_�� t$�@�3�Y|( A���W��
ѻ� �3� T0 k� ��=��=e1�t B�1	�"q  ��/    �����OמIo�� t$�?�7�Y|( A���W��
ѿ� �3� T0 k� ��>��>e1�t B�1	�"q  ��/    �����OלIo�� t$�>�;�Y|( A���W��
ѿ� �3� T0 k� ��?��?e1�t B�1	�"q  ��/    �����OӛIo�� t$�=�C�Y|( A���W��
ѿ� �3� T0 k� ��@��@e1�t B�1	�"q  ��/    �����OӚIo�� t$�<�G�Y|( A���W��
ѿ� �3� T0 k� ��A��Ae1�t B�1	�"q  ��/    �����OϘIo�� t%�;�K�Y|( A���W��
ѿ� �3� T0 k� ��A��Ae1�t B�1	�"q  ��/    �����OϗI_�� t%�9�O�Y|( A���W��
ѿ� �3� T0 k� ��B��Be1�t B�1	�"q  ��/    �����O˖I_�� t%�8�S�Y|( A���V��
ѿ� �3� T0 k� ��C��Ce1�t B�1	�"q  ��/    �����O˕I_�� t%�7�W�Y|( A���V��
ѿ� �3� T0 k� ��D��De1�t B�1	�"q  ��/    �����OǔI_�� t%�6�W�Y|( A���V��
ѿ� �3� T0 k� ��D� De1�t B�1	�"q  ��/    �����OǓI_�� t%|�5�W�Y|( A���V��
�ü �3� T0 k� � E�Ee1�t B�1	�"q  ��/    �����OÑIo�� t%|�3�W�Y|( A���V��
�ü �3� T0 k� �F�Fe1�t B�1	�"q  ��/    �����OÐIo�� t%|�2�[�Y|( A���V��
�ü �3� T0 k� �G�Ge1�t B�1	�"q  ��/    �����O��Io�� t%|�1�[�Y|( A���V��
�ü �3� T0 k� �H�He1�t B�1	�"q  ��/    �����O��Io�� t%|�0�_�Y|( A���V��
�ü �3� T0 k� �H�He1�t B�1	�"q  ��/    �����O��Io�� t%|�/�_�Y|( A���V��
�ü �3� T0 k� �I�Ie1�t B�1	�"q  ��/    �����O��I_�� t%|�.�_�Y|( A���V��
�ü �3� T0 k� �J�Je1�t B�1	�"q  ��/    �����O��I_�� t%|�-�c�Y|( A���V��
�ü �3� T0 k� �K� Ke1�t B�1	�"q  ��/    �����O��I_�� t%|�,�c�Y|( A���V��
�ü �3� T0 k� �L� Le1�t B�1	�"q  ��/    �����O��I_�� t%|�+�c�Y|( A���V��
�ü �3� T0 k� � L�$Le1�t B�1	�"q  ��/    �����O��Io�� t%} )�c�Y|( A���V��
�Ǽ �3� T0 k� �(N�,Ne1�t B�1	�"q  ��/    �����O��Io�� t%}(�g�Y|( A���V��
�Ǽ �3� T0 k� �,O�0Oe1�t B�1	�"q  ��/    �����O��Io�� t%}'�g�a�( A���V��
�Ǽ �"�� T0 k� �0O�4Oe1�t B�1	�"q  ��/    �����O��Io�� t%�&�g�a�( A���V��
�Ǽ #�"�� T0 k� �4P�8Pe1�t B�1	�"q  ��/   �����O��Io�� t%�%�g�a�( A���V��
�Ǽ #�"�� T0 k� �8Q�<Qe1�t B�1	�"q  ��/    �����O��Kߧ� t%�$�g�a�( A���V��
�Ǽ #�"�� T0 k� �<R�@Re1�t B�1	�"q  ��/    �����O��K߫� t%�#�g�a�( A��� V��
�Ǽ #�"�� T0 k� �@R�DRe1�t B�1	�"q  ��/    �����O��K߫� t%� "�g�a�( A��� V��
�Ǽ #�"�� T0 k� �DS�HSe1�t B�1	�"q  ��/    �����O��K߫� t%�$!�g�a�( A��� V��
�Ǽ #�"�� T0 k� �DT�HTe1�t B�1	�"q  ��/    �����O��K߫� t%�( �k�a�( A��� V��
�Ǽ #�"�� T0 k� �HU�LUe1�t B�1	�"q  ��/    �����O��K߫� t%�,�k�a�( A��� V��
�Ǽ #�"�� T0 k� �LU�PUe1�t B�1	�"q  ��/    �����O��K߯� t%�0�k�a�( A��� V��
�Ǽ #�"�� T0 k� �PV�TVe1�t B�1	�"q  ��/    �����O��K߯� t%�4�k�a�( A��� V��
�Ǽ #�"�� T0 k� �TW�XWe1�t B�1	�"q  ��/    �����O��K߯� t%�8�o�Y|( A��� U��
�˼ #�3� T0 k� �XX�\Xe1�t B�1	�"q  ��/    �����O��K߯� t%�<�o�Y|( A��� U��
�˼ #�3� T0 k� �\Y�`Ye1�t B�1	�"q  ��/    �����O��K߯� t%�@�s�Y|( A��� U��
�˼ #�3� T0 k� �`Y�dYe1�t B�1	�"q  ��/    �����?��Kﳢ t%�D�s�Y|( A��� U��
�˼ #�3� T0 k� �dZ�hZe1�t B�1	�"q  ��/    �����?��Kﳢ t%�H�w�Y|( A��� U��
�˼ #�3� T0 k� �h[�l[e1�t B�1	�"q  ��/    �����?��Kﳢ t%�L�w�Y|( A����U��
�˼ #�3� T0 k� �h\�l\e1�t B�1	�"q  ��/    �����?��Kﳢ t%�P�w�Y|( A����U��
�˼ #�3� T0 k� �l\�p\e1�t B�1	�"q  ��/   �����?��Kﳢ t%�T�w�Y|( A����U��
�˼ #�3� T0 k� �p]�t]e1�t B�1	�"q  ��/    �����?��K﷢ t%�X�{�Y|( A����U��
�˼ '�3� T0 k� �t^�x^e1�t B�1	�"q  ��/   �����o��K﷣ t%�\�{�Y|( A����U��
�˼ '�3� T0 k� �x_�|_e1�t B�1	�"q  ��/    �����o��K﷣ t&�`��Y|( A����U��
�˼ '�3� T0 k� �|_��_e1�t B�1	�"q  ��/    �����o��Kﻣ t&�d��a�( A����U��
�˼ '�"s� T0 k� �`��`e1�t B�1	�"q  ��/    �����o��Kﻣ t&�h���a�( A����U��
�˼ '�"s� T0 k� �a��ae1�t B�1	�"q  ��/    �����o��Kﻣ t&�h���a�( A����U��
�˼ '�"s� T0 k� �a��ae1�t B�1	�"q  ��/    �����_��K￣ t&�l���a�( A����U��
�˼ '�"s� T0 k� �b��be1�t B�1	�"q  ��/    �����_��K￣ t&�p���a�( A����U��
�˼ '�"s� T0 k� �c��ce1�t B�1	�"q  ��/    �����_��K�ã t&�t���a�( A����U��
�ϼ '�"s� T0 k� �d��de1�t B�1	�"q  ��/    �����_��K�ã t&�x���a�( A����U��
�ϼ '�"s� T0 k� �d��de1�t B�1	�"q  ��/    �����_��K�ä t&�x���a�( A����U��
�ϼ '�"s� T0 k� �e��ee1�t B�1	�"q  ��/    �����_�K�Ǥ t&�|���a�( A����U��
�ϼ '�"s� T0 k� �f��fe1�t B�1	�"q  ��/    �����O{�K�Ǥ t&�����a�( A����U��
�ϼ '�"s� T0 k� �g��ge1�t B�1	�"q  ��/    �����Ow�K�Ǥ t&�����a�( A����U��
�ϼ '�"s� T0 k� �g��ge1�t B�1	�"q  ��/    �����Os�K�ˤ t&�����Y|( A����U��
�ϼ '�3� T0 k� �h��he1�t B�1	�"q  ��/    �����Os�K�ˤ t&�����Y|( A����U��
�ϼ '�3� T0 k� �i��ie1�t B�1	�"q  ��/    �����Oo�K�Ϥ t&�����Y|( A����U��
�ϼ '�3� T0 k� �j��je1�t B�1	�"q  ��/    �����Ok�K�ϥ t&�����Y|( A����U��
�ϼ '�3� T0 k� �j��je1�t B�1	�"q  ��/    �����Og�K�ӥ t&�����Y|( A����U�|
�ϼ '�3� T0 k� �k��ke1�t B�1	�"q  ��/    �����Oc�K�ӥ t&��
���Y|( A����U�|
�ϼ '�3� T0 k� �l��le1�t B�1	�"q  ��/    �����?_�K�ӥ t&��
���Y|( A����U�|
�ϼ '�3� T0 k� �l��le1�t B�1	�"q  ��/    �����?[�K�ץ t&��	���Y|( A����U�|
�ϼ '�3� T0 k� �m��me1�t B�1	�"q  ��/    �����?W�K�צ�t&��	���Y|( A����U�| 
�ϼ '�3� T0 k� ��n��ne1�t B�1	�"q  ��/    �����?S�K�ۦ�t&}����Y|( A����U�| 
�ϼ '�3� T0 k� ��o��oe1�t B�1	�"q  ��/    �����?O�K�ۦ�t&}����Y|( A����U�| 
�ϼ +�3� T0 k� ��o��oe1�t B�1	�"q  ��/    �����?K�K�ۦ�t&}����Y|( A����U�| 
�ϼ +�3� T0 k� ��p��pe1�t B�1	�"q  ��/    �����?G�K�ߦ�t&}����Y|( A����U�| 
�ϼ +�3� T0 k� ��q��qe1�t B�1	�"q  ��/    �����?C�K�ߦ�t&}�ϯ�Y|( A����U�| 
�ϼ +�3� T0 k� ��q��qe1�t B�1	�"q  ��/    �����??�K�ߦ�t&}�ϳ�Y|( A����U�| 
�Ӽ +�3� T0 k� ��r��re1�t B�1	�"q  ��/    �����/;�K���t&ݬϳ�Y|( A����U�| 
�Ӽ +�3� T0 k� ��s��se1�t B�1	�"q  ��/    �����/7�K���t&ݰϷ�Y|( A����U�| 
�Ӽ +�3� T0 k� ��t��te1�t B�1	�"q  ��/    �����/7�K���t&ݰϷ�Y|( A����U�| 
�Ӽ +�3� T0 k� ��t��te1�t B�1	�"q  ��/    �����/3�K���t&ݴϻ�Y|( A����U�| 
�Ӽ +�3� T0 k� ��u��ue1�t B�1	�"q  ��/    �����//�K���t&ݸϻ�Y|( A����U�| 
�Ӽ +�3� T0 k� ��v��ve1�t B�1	�"q  ��/    �����//�K���t&ݼϿ�Y|( A����U�| 
�Ӽ +�3� T0 k� ��v��ve1�t B�1	�"q  ��/    �����/+�K���t&��Ͽ�Y|( A����U�| 
�Ӽ +�3� T0 k� ��w��we1�t B�1	�"q  ��/    �����/+�K���t&���ÛY|( A����U�| 
�Ӽ +�3� T0 k� ��x��xe1�t B�1	�"q  ��/    �����/+�K���t&�� �ÛY|( A����U�| 
�Ӽ +�3� T0 k� ��x��xe1�t B�1	�"q  ��/    �����/'�K���t&����ÛY|( A����U�| 
�Ӽ +�3� T0 k� ��y��ye1�t B�1	�"q  ��/    �����/'�K���t&����ǛY|( A����U�| 
�Ӽ +�3� T0 k� ��z��ze1�t B�1	�"q  ��/    �����'�K���t&����ǛY|( A����U�| 
�Ӽ +�3� T0 k� ��{� {e1�t B�1	�"q  ��/    �����'�K���t&����˛Y|( A����U�| 
�Ӽ +�3� T0 k� � {�{e1�t B�1	�"q  ��/    �����#�K���t&����˛Y|( A����U�| 
�Ӽ +�3� T0 k� �|�|e1�t B�1	�"q  ��/    �����#�K���t&����˛Y|( A����U�| 
�Ӽ +�3� T0 k� �}�}e1�t B�1	�"q  ��/    �����#�K���t&����˛Y|( A����U�| 
�Ӽ +�3� T0 k� �}�}e1�t B�1	�"q  ��/    ������#�K���t&����˛Y|( A����U�| 
�Ӽ +�3� T0 k� �~�~e1�t B�1	�"q  ��/    ������#�K����t&����˛Y|( A����U�| 
�Ӽ +�3� T0 k� ��e1�t B�1	�"q  ��/    ������#�K����t&����ϚY|( A����U�| 
�Ӽ +�3� T0 k� ��e1�t B�1	�"q  ��/    �������K����t&����ϚY|( A����U��
�Ӽ +�3� T0 k� ����e1�t B�1	�"q  ��/    �������K����t&����ϚY|( A����U��
�Ӽ +�3� T0 k� ����e1�t B�1	�"q  ��/    �������A���t&����ӚY|( A����U��
�Ӽ +�3� T0 k� ��� �e1�t B�1	�"q  ��/    �������A���t&���ӚY|( A����U��
�Ӽ +�3� T0 k� � ��$�e1�t B�1	�"q  ��/    �������A���t&���ӚY|( A����U��
�Ӽ +�3� T0 k� �$��(�e1�t B�1	�"q  ��/    �������A���t&���ӚY|( A����U��
�Ӽ +�3� T0 k� �(��,�e1�t B�1	�"q  ��/    �������A���t&���ךY|( A����T��
�׼ +�3� T0 k� �(��,�e1�t B�1	�"q  ��/    �������A_���t&���ךY|( A����T��
�׼ +�3� T0 k� �,��0�e1�t B�1	�"q  ��/    �������A_���t&���ךY|( A����T��
�׼ +�3� T0 k� �0��4�e1�t B�1	�"q  ��/    �������A_���t&�'��ۚY|( A����T��
�׼ +�3� T0 k� �4��8�e1�t B�1	�"q  ��/    �������A_���t&�+��ۚY|( A����T��
�׼ /�3� T0 k� �8��<�e1�t B�1	�"q  ��/    �������A_���t&�/��ۚY|( A����T�{�
�׼ /�3� T0 k� �8��<�e1�t B�1	�"q  ��/    �������K���t&�7��ۚY|( A����T�{�
�׼ /�3� T0 k� �<��@�e1�t B�1	�"q  ��/    �������K��t&�;��ۚY|( A����T�{�
�׼ /�3� T0 k� �@��D�e1�t B�1	�"q  ��/    �������K��t&�C��ۚY|( A����T�{�
�׼ /�3� T0 k� �D��H�e1�t B�1	�"q  ��/    �������K��t&G��ۚY|( A����T�{�
�׼ /�3� T0 k� �D��H�e1�t B�1	�"q  ��/    �������K��t&O��ۚY|( A����T�{�
�׼ /�3� T0 k� �H��L�e1�t B�1	�"q  ��/    �������K?��t&W��ߚY|( A����T�{�
�׼ /�3� T0 k� �L��P�e1�t B�1	�"q  ��/    �������K?��t&[��ߚY|( A����T�{�
�׼ /�3� T0 k� �P��T�e1�t B�1	�"q  ��/    �������K?��t&c��ߚY|( A����T�{�
�׼ /�3� T0 k� �P��T�e1�t B�1	�"q  ��/    �������K?��t&g��ߙY|( A����T�{�
�׼ /�3� T0 k� �T��X�e1�t B�1	�"q  ��/    �������K?��t&o��ߙY|( A����T�{�
�׼ /�3� T0 k� �X��\�e1�t B�1	�"q  ��/    �������Ko��t&s���Y|( A����T�{�
�׼ /�3� T0 k� �\��`�e1�t B�1	�"q  ��/    �������Ko��t&{���Y|( A����T�{�
�׼ /�3� T0 k� �\��`�e1�t B�1	�"q  ��/    �������Ko��t&����Y|( A����T�{�
�׼ /�3� T0 k� �`�de1�t B�1	�"q  ��/    �������Ko��t&����Y|( A����T�{�
�׼ /�3� T0 k� �d�he1�t B�1	�"q  ��/    �������Ko��t&�� o�Y|( A����T�{�
�׼ /�3� T0 k� �h�le1�t B�1	�"q  ��/    �������J��t&�� o�Y|( A����T�{�
�׼ /�3� T0 k� �h�le1�t B�1	�"q  ��/    �������J��t&�� o�Y|( A����T�{�
�׼ /�3� T0 k� �l�pe1�t B�1	�"q  ��/    �������J��t&�� o�Y|( A����T�{�
�׼ /�3� T0 k� �p�te1�t B�1	�"q  ��/    �������J��t&�� o�Y|( A����T�{�
�׼ /�3� T0 k� �t�xe1�t B�1	�"q  ��/    �������J��t&�����Y|( A����T�{�
�׼ /�3� T0 k� �t~�x~e1�t B�1	�"q  ��/    �������J��t&�����Y|( A����T�{�
�׼ /�3� T0 k� �x~�|~e1�t B�1	�"q  ��/    �������J��t&�����Y|( A����T�{�
�׼ /�3� T0 k� �|~��~e1�t B�1	�"q  ��/    �������J��t&�����Y|( A����T�{�
�׼ /�3� T0 k� �~��~e1�t B�1	�"q  ��/    �������K�� t&�����Y|( A����T�{�
�׼ /�3� T0 k� �~��~e1�t B�1	�"q  ��/    �������K�� t&�����Y|( A����T�{�
�׼ /�3� T0 k� �~��~e1�t B�1	�"q  ��/    ��������@�?� �� W� l�Z<?�Lm�����1���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�?� �� W� l�Z<?�Lm�,����1���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�?� �� W� l�Z<?�Lm�,����1���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�?� �� W� l�Z<?�Lm�,����1���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�?� �� W� l�Z<?�Lm�,����1���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�?� �� W� l�Z<?�Lm�,����1���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�C� �� W� l�Z<?�Lm� �����0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�C� �� W� l�Z<?�Lm� �����0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�C� �� W� l�Z<?�Lm� �����0���3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�C� �� W� l�Z<?�Lm� �����0����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�C� �� W� l�Z<?�Lm� �����0�����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�C� �� W� l�Z<?�Lm� �����0�����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�C� �� W� l�Z<?�Lm� �����0�����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�G� �� W� l�Z<?�Lm� �����0�����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�G� �� W� l�Z<?�L]� �����0�����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�G� �� W� l�Z<?�L]� �����0�����3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�G� �� S� l�Z<?�L]� �����0����#�3� T0 k� ��#�P e1�t B�1	�"q ��/    ����8���@�G� �� S� l�Z<?�L]�����0����#�3� T0 k� ��$P e1�t B�1	�"q ��/    ����8���@�G� �� S� l�b|?�L]�����0���]#�3� T0 k� ��$P e1�t B�1	�"q ��/    ����8���@�G� �� S� l�b|?�L]�����0���]�3� T0 k� ��$P e1�t B�1	�"q ��/    ����8���@�G� �� S� l�b|?�A�#�����0���]�3� T0 k� ��$P e1�t B�1	�"q ��/    ����8���@�G� �� S� l�b|?�A�#�����0���]�3� T0 k� ��$P e1�t B�1	�"q ��/    ����8���@�K� �� S� l�b|?�A�#�����0���]�3� T0 k� ��#;P e1�t B�1	�"q ��/    ����8                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \���$ ]�)�)� � �#����   � �
     ���֨    ��Z�����    
�	�              ����           ��    ���   0		 
 
         ��2�  � �
   ���|C    ��A���    ���          P����           ��     ���  (	 
           &��          ��&�     &����&�                   p �����         �     ���  8�         �Ġd   * *	     ��i�    ���w����    �h   	           5  ����           ��   
  ���  (
	         ��{   \ [     .����    �������h    KZ             ����          ��     ��� P
B            �� ��     B�
'?      ���
'?                             ���P         @    m  ���    81
           ��Z�       V (�8    ��] (��    �� $                 �8         �     ��H   8	           T�	    	    j�|��     T�	�|��      ��                 l ;         ��     ��@   0	          ��F�          ~����    ��I�����    ����             �� D               ��@   8
	          ���V  � �	     � u�p    ���V u�C       ]               �� �         	 �@
`     ��P   @

	(		         ���          � K��    ��� K��       H                  �         
  ��     ��@   H
	 		           K> ��
	      � ��      K> ��                             ���o              m  ��@    8

 '                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          ~h  ��        � ��     ~C� ��    ��+                  x                j  �   �   �                          ~    ��        � �       ~   �           "                                                �                         �����������
 (�|�� u K ��� � �       	    
      
    "{. X�D       � �c@ � d@ � d` �d  _����. ����< ����J ����X � �  _� �D _� �� ]`��� ����  ����. ����< ����J ����X � � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� � }`���� � � }`���� � xD �o� yD  p� y� 0q  y� q` �d �^@ �d _@  � �m@ � n@ �d �[� �d \� � �j� � k� �D }@ � }` � �c@ � d@ �� �`� �� a� � a����� � �� _� � �m@ �  n@ �� �j� �� k� 
� V� 
�< V� 
�\ W  
�\ W� 
�� W� 
�\ W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ������������   ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"    B�j
��  B �
� �  �  
� ��    ��     �   �    &    ��     ���      ��    ��     � (          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �/�      ��T ���        �/T ���        �        ��        �        ��        �    ��     v 7 ��        ��                         I:  # 
����                                    �                 ����            �� ���%��  ������               13 Mats Sundin lik     0:14                                                                        3  2      �IcjTa crL'c~ �< c� �C �) C" � C# �B� � �	C$ �	
J� � �J� � �J� � �	C. � �C4 � �C6 � �kV � � k^ � xc� � Lc� � l c� � D c� �
"�
 "�1 �"� �*�* �"� � � "� � �� � � 
� � �� � � 
� � �  "� � �!� � � 
� � �#� � � 
� � � 
� � � &"� � �'� � � 
� � � 
� � � 
� � � 
� � � 
� � 
� �X  "K �X  "H �X  "K �X  "K �X  "G rP 3"C zX 4"G rX  "K � � 6b� ~ � 7b� ~ �8b` � � b^ � �  b� � �  b� � � <b� � � =b� � � >b� � � bt �                                                                                                                                                                                                                         t� P         �    @ 
        "     c P E g  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    �{T�� ��������������������������������������������������������   �4, P� 0 5� ���� ���� A*�������&���                                                                                                                                                                                                                                                                                                                          ��
�@;"@z�p�                                                                                                                                                                                                                                   	 " +    � �  L�J       (                             �������������������������������������������������������                                                                    	                                                                  �    ��             �   !      �   �             	 	 ������ ������� ������������ ���������� �� ����� ���� ������������������� ��� � �������������  ������������������������ ����� � � ����������������������� ���������������� ������  �������� ������������������� ��������������������                      	     A  
  %     �  9<�J      ��                             ������������������������������������������������������                                                                                                                                           �  6�                  9 P    ��                   ���������� ������������������������ ������� ��������������������������� ������� ���� ����������� ������ ������ ����������� ���������������������� ��������������� �������� ������ ������������������ ������ ���� ��� ���������������� ��            �                                                                                                                                                                                                                                         
                                                                     �             


             �  }�                    R�                                                       'v            ������������  +������������������������������������       ��������������������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" " L ?                                 � E��_ �`�                                                                                                                                                                                                                                                                                          )n)nE  �                d      m      k                                                                                                                                                                                                                                                                                                                                                                                                                                        > �  
>�  
�  2�  2�  EZmk ��� r�������H�n����{�̞� �N I�����8����;a        6   }�> :��		         �   & AG� �   �              �4�                                                                                                                                                                                                                                                                                                                                        I G   �                     !��                                                                                                                                                                                                                            Y   �� �� Ѱ��      �� 4      ������ ������� ������������ ���������� �� ����� ���� ������������������� ��� � �������������  ������������������������ ����� � � ����������������������� ���������������� ������  �������� ������������������� ������������������������������ ������������������������ ������� ��������������������������� ������� ���� ����������� ������ ������ ����������� ���������������������� ��������������� �������� ������ ������������������ ������ ���� ��� ���������������� ��     �     $�l�������l����������������������l��������������f���f���f��ff���f������ffffflffffffffffffffffffff����ff��lfflffffffffffffffffffffl��l��̼���l����l��lf���ll��������l�����ll������l�����������������l���������������l��������������fff�lff�ll��l���li��f���l���f��ffffffffffff��������������������fffffff�ffl��̻�����������������f�l���l�llll�l�̦ll̜f�̊�l̊���l����������������������������������������������������������������f���f���f���f���f���f��ɜ�����������������������̺��ƹ��li��fiy��������������˩�ff��fl��fk��fj���f̈�f̈�f̈�f̈�fl�{ʜ�����������l����������������̼��������������������������������������̼̼��������j���ˊ��̗��̸���ʈ���Ɉ��i���������������������������y��fj���k���̨��̹��l���̹��lɹ��ʘ�����ɬ��ȼ�������l���̘��̈���������̼����̼������̼�����̼��������������̼���������̼���̼̼���k�̼̈��̈��ˈ��˘̼����˘��̘�Ɉ����������������ˈ�����������k��ɫ��ɫ����ff��ɶ��ɻ�ll���������̉��ˈ��̈��̙��ˈ�̼���l�����������������̼����˼�̶���̻�������������˨̩��������������������ʈ����������|����i����Ʒi��i��������������������������j���f��������̹�̼���̘�fʘ��ɉ����̊�̼��ȸ�{�Ɉ��h�����l���j���h��fȹ����̈xx�������������f���l��l�������    6      6   �� ~                       4     �   �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$    `d  �@���6 ��  �@���6 �$ ^$ �s@  �@  �s@   o 
�� ��   o 
   ���   ����  ��   ����  �$ ^$�� �   �         �   /       H `� ބ �� `� ބ **� �  �� �       �  ��   l�����������J   g��� 
        f ^�         �� ��      l      �����������J���J������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  "!  " ! " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "! ""! " ""  "!  "! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  "!  " ! " ""  !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                       ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .   ��  �   ��  �                    �     �                              �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                             "  "(��ȩ�ܚ��ۊ����� ��  �   �   �   �   �� ��� ̻� ˽� ��� �w� �������������������������� �̻ ���         �   �       �   �   "" �+� Ȼ� ɫ� ɨ� ��                �� �I��3 ��D 
UD 
UD TD  T�  ˸  ��  �� ̰ �+ ��"/ �"/  ����  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �                    �               �  �  ��  �   �   �                    �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                    �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   ��  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �   �   �                .                        �   �      ��   �  ��  �  �  �         � �������������  �              � � ��      �                                                                                                                                  
      �  �  ��  �� �� �� 	�� D� EH EZ  DZ 4J 34Z3EH�T��ʄ
����ܩ���� ""�""�""�"/� �� �  ��� ̽� ��� �w� ��� ��� ��� ˻���ܚ��ة��ی����˻ݼˍ�ۻ���Ѕ" �" R�  B      ��  ��  �     �            � �� �   �       �   ��  ��  ��  ���        �                                      �                             ���                         �  ��                    �����                                                                                                                                                                                                                                    
  �  ̈ �� ,�  ""   "                       �������݅]̻�U�˅U3�U\�BU\�3 "��",�"��"��� ��  �             ݽ���۹����" ��" ��"��".�  �"  �/� .���" � ��              �   .   �   � � �� �� ��                    ��  ��  ���            � ˹ Y�����
�ڛ��٩ �� �̽���ݪ۽w�}�֪�vv���p���             "   "   "       �         �        �   �     �       �   �   �   �   �      �                    ��� ���� ��             �  �˰ ��� �wp ���                                                                                                                                                                                         �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                   �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �   �   "   "   "  !�    ��                ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                                                                                                                                                                    �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                   � ��                  �  �˰ ��� �wp ��� �   �   �   �                               �    �    ��                        �  �  �                                                                 �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �  "������"    /   �  �   ��                                �   �                      �������  ���    � �� �  �  �      �   �                       ���                     �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                          ̻  ��  rb  wg 
�w ���
���ɛ������̽�̪��̙���̻̽̽���٘"#3 ""DR�U� T� �� 	��  ��  ,� "� "� ""��""�������� �  ��   �   p   z   ��  ��  ��� �̹ �ؚ �ک ��������������32"�D2" UR" EU@ EU@ 4U@ K˰ 
�� ��  �   "   ""  "" ��"/���� �� �     ��  ��  ��  ��  ��  ��  �                             �� ̽��  ��  �   �                        �  ��� ̻� ��� rbp wgz�               �������  ���    �                       � ��                  �  �˰ ��� �wp ���      � ���� ��   � � �                                                                                                                                    �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �    �   ��  �  ��  �             �  �   �   ��  �                                        ��                  �                        ���� ��� ����                               � ��                  �  �˰ ��� �wp ��� �   �   �   �                               �    �    ��                        �  �  �                                                                         �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��                  �          �         �   �  �  �   �               �   �                     �                        �         �  �� �  �� ��                                                                                                                                                   �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""������������������""""������������������������""""������������������������""""������ADAIA�A""""�������I�A�A�A""""�����DD�I""""�������DAADAI""""������IDA��""""��������DD��I�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD������������������������3333DDDD�A�AM�M�DM��M334CDDDD�A�AM�M�DDM����3333DDDDDM����DD�����3333DDDDMAM��D�DDM�����3333DDDDDD����M��DM�����3333DDDD������������DD������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ADA�LL��L�D����3333DDDD x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(XxLL����������D����3333DDDD w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""����������A������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(""""�������I�I������ �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�""""�������I��D���I������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`�D�M�D���M������3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(MD�M�A�����MD�����3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(�""""�����AMAD������ � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(�""""������������������ � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqIcjTa crL'c~ �< c� �C �B� � �B� � �B� � �	C$ �	
J� � �J� � �J� � �	C. � �C4 � �C6 � �kV � � k^ � xc� � Lc� � l c� � D c� �
"�
 "�1 �"� �*�* �"� � � "� � �� � � 
� � �� � � 
� � �  "� � �!� � � 
� � �#� � � 
� � � 
� � � &"� � �'� � � 
� � � 
� � � 
� � � 
� � � 
� � 
� �X  "K �X  "H �X  "K �X  "K �X  "G rP 3"C zX 4"G rX  "K � � 6b� ~ � 7b� ~ �8b` � � b^ � �  b� � �  b� � � <b� � � =b� � � >b� � � bt �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0�������������������������������������������;�O�I�N�G�X�J��<�S�K�N�R�O�Q� � � � � �,�>�0�������������������������������������������7�G�Z�Y��<�[�T�J�O�T� � � � � � � � � �:�>�/�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������:�>�/� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������,�>�0� �� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            