GST@�                                                            \     �                                                ���                        ����e ��	 J���������������~���        h     #    ~���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    
 �j,� B ��
                                                                                 ����������������������������������      ��    ooo  gog    +      '       ���                  	 7 V 	                 ��          8:8�����������������������������������������������������������������������������������������������������������������������������o=  0  o4   1  +      '           �                    	�  7�  V�  	�                  n  	          : �����������������������������������������������������������������������������                                ��  k   �  $�   @  #   �   �                                                                                '     ��  	n    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E s �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    D�p��D������{�|;�D��E��C��.JBߩ>�3��T0 k� �'��+�%�0d  851t"Q  ��G    �����D�p��D��m���w�|;�D��E�C��-@�ߩ>ې3��T0 k� �'��+�%�0d  851t"Q  ��G    �����D�q���D��m���o�|;�C��E�C��-@�ߩ>א3��T0 k� �'��+�%�0d  851t"Q  ��G    �����D�q��D��m���k�|;�C�w�E�C��,@�ߩ>Ӑ3��T0 k� �#��'�%�0d  851t"Q  ��G    �����D�q��D��m���g�|;�C�o�E�EO�+@�ߩ>ˏ3��T0 k� �#��'�%�0d  851t"Q  ��G    �����D�r��D��m���_�|;�C�g�E�EO�*@�ߩ>Ǐ3��T0 k� �#��'�%�0d  851t"Q  ��G    �����D�r�ۈD��m���[�|;�C�_�E�EO�)Aߩ>Î3��T0 k� �#��'�%�0d  851t"Q  ��G    �����D�r�ψD��m��W�|;�C�W�B�EO�(Aߩ3��T0 k� ����%�0d  851t"Q  ��G    �����Dxs@ǉD����O�|;�C�O�B�EO�'Aߩ3��T0 k� ����%�0d  851t"Q  ��G    �����Dht@��D����G�|;�C�?�B�EO�%Aߩ3��T0 k� ����%�0d  851t"Q  ��G    �����D`t@��D����C�|;�C�;�B�EOx$ARߩ3��T0 k� ����%�0d  851t"Q  ��G    �����DXt@��D����?�|;�C�3�E�EOp$ARߩ3��T0 k� ����%�0d  851t"Q  ��G    �����DPu@��D����;�|;�C�+�E�EOh#ARߩ3��T0 k� ����%�0d  851t"Q  ��G    �����DHu@��C����7�|;�C�#�E�E?`"ARߩ3��T0 k� ����%�0d  851t"Q  ��G    �����D@u@��C����3�|;�C��E�E?X!ARߩ3��T0 k� ����%�0d  851t"Q  ��G    �����C�8v@��C�w���3�|;�C��E�E?PD2ߪ���3��T0 k� ����%�0d  851t"Q  ��G    �����C�0v�{�C�o���/�|;�C��Eo�E?HD2ߪ�{�3��T0 k� ����%�0d  851t"Q  ��G    �����C�(v�s�C�c�����+�|;�C��Eo�E?@D2۪�w�3��T0 k� ������%�0d  851t"Q  ��G    �����C�w�c�C�S��{��'�|;�EO�Eo�E?4D2۪�k�3��T0 k� ������%�0d  851t"Q  ��G    �����C�w�[�C�K��w��#�|;�EO�Eo�E?,C�۪�c�3��T0 k� ������%�0d  851t"Q  ��G    �����C�w�O�C�C��s��#�|;�EO�A��E?$C�ת�_�3��T0 k� ������%�0d  851t"Q  ��G    �����C� x�G�C�;��s��#�|;�EO۴A��COC�׫�_�3��T0 k� ������%�0d  851t"Q  ��G    �����C��x�?�C�/��o���|;�EOӴA���COC�׫�[�3��T0 k� ������%�0d  851t"Q  ��G    �����C��x�7�C�'��k���|;�C�˴A���COC�ӫ�[�3��T0 k� ������%�0d  851t"Q  ��G    �����C��y�/�C���k���|;�C�ôA���COC�ӫ�W�3��T0 k� ������%�0d  851t"Q  ��G    �����C��y��C���g���|;�C���En��I^�C�ӫS�3��T0 k� ������%�0d  851t"Q  ��G    �����C��y��C���g���|;�C���En�I^�C�ϫO�3��T0 k� ������%�0d  851t"Q  ��G    �����C��z��C����c���|;�EO��En�I^�C�ϬO�3��T0 k� ������%�0d  851t"Q  ��G    �����C��z��C����c���|;�EO��En�I^�C�ϬO�3��T0 k� ������%�0d  851t"Q  ��G    ����C�z���C����c���|;�EO��En��I^�
C�ˬK�3��T0 k� ������%�0d  851t"Q  ��G    ����~C�{��C����_���|;�EO��En��I^�	C�ˬK�3��T0 k� ������%�0d  851t"Q  �G    ����C�{��C����_���|;�EO�E^��In�C�ˬG�3��T0 k� .�����%�0d  851t"Q ��O    �����C�{�ۑE����_���|;�EOw�E^��In�C�ǬG�3��T0 k� .�����%�0d  851t"Q ��O    �����C�|�ϑE޿��_���|;�EOo�E^��In�C�ǬC�3��T0 k� .�����%�0d  851t"Q ��O    �����C��|�ǑE޷��_����|;�E?g�E^��In�C�íC�3��T0 k� .�����%�0d  851t"Q ��O    �����C��|߿�Eޯ��_����!�;�E?_�E^��In�C�íNC�3��T0 k� .�����%�0d  851t"Q ��O    �����D ||߷�Eާ��[����!�;�E?W�E���E>�C�NC�3��T0 k� .�����%�0d  851t"Q ��O    �����D x}﯒Eޟ��[����!�;�E?S�E���E>�C�N?�3��T0 k� ������%�0d  851t"Q ��O    �����D h}Eދ��[����!�;�I_C�E���E>��C�N?�3��T0 k� ������%�0d  851t"Q ��O    �����D `}Eރ��[����!�;�I_?�E���E>��D�� ?�3��T0 k� ������%�0d  851t"Q ��O    �����D X}E�{��[����!�;�I_7�E��E>��D�� ?�3��T0 k� ������%�0d  851t"Q ��O    �����D P~O��E�s� m[����!�;�I_3�E��E>��D�� ?�3��T0 k� >�����%�0d  851t"Q ��O    �����D H~O{�I�k� m[����!�;�I_+�E��E>��D�� ?�3��T0 k� >�����%�0d  851t"Q ��O    �����D @~Os�I�c� m[�M��!�;�Io'�E��E>��D�� ?�3��T0 k� >�����%�0d  851t"Q ��O    �����D 8~Ok�I�[� m[�M��!�;�Io#�E��E.��D���?�3��T0 k� >�����%�0d  851t"Q ��O    �����D 0~Oc�I�S� m[�M��|;�Io�D>��E.��D���?�3��T0 k� >�����%�0d  851t"Q ��O    �����D(O[�I�K�M[�M��|;�Io�D>��E.��D���?�3��T0 k� ������%�0d  851t"Q ��O    �����D OS�I�G�M[�M�|;�Io�D>��E.��D���?�3��T0 k� ������%�0d  851t"Q ��O    �����DOC�I�7�M[�M�|;�I_�D>��E.��D���C�3��T0 k� ������%�0d  851t"Q ��O    �����D?;�I�3�M[�M�|;�I_�D>��E.��D���C�3��T0 k� ������%�0d  851t"Q ��O    �����D �?3�I�+�M[�M�|;�I_�D>��E.��D���C�3��T0 k� .�����%�0d  851t"Q ��O    �����D�?+�I�'�M[�M�|;�I_�D>{�E.��D��G�3��T0 k� .�����%�0d  851t"Q ��O    �����D�?#�I��M[���|;�I^��E�w�E.��D{��G�3��T0 k� .�����%�0d  851t"Q ��    �����D�?�I��M[���|;�In��E�o�E.��Ds��K�3��T0 k� .�����%�0d  851t"Q ��    �����E_�?�I���[���|;�In��E�g�E.��Do��K�3��T0 k� .�����%�0d  851t"Q ��    �����E_�~?�I���[���!�;�In��E�_�E��Dg�O�3��T0 k� ������%�0d  851t"Q ��    �����E_�~?�I���[���!�;�In�E�O�E��D_�S�3��T0 k� ������%�0d  851t"Q ��    �����E_�~?�I���[���!�;�A�E�G�E��DW�S�3��T0 k� ������%�0d  851t"Q ��    �����E_�~N��I����[���!�;�A�E�?�E��DO�W�3��T0 k� ������%�0d  851t"Q ��    �����E_�}N��I����[���!�;�A�E�;�E��C�K�[�3��T0 k� N�����%�0d  851t"Q ��    �����E_�}N�I����[���!�;�A�E�3�E��C�C�_�3��T0 k� N�����%�0d  851t"Q ��    �����E_�}N�I����[���!�;�A߰E�3�E��C�;�_�3��T0 k� N�����%�0d  851t"Q ��    �����E_�}N�I����[���!�;�E�߱E�+�B���C�7�c�3��T0 k� N�����%�0d  851t"Q ��    �����E_�|>ߠI����[���!�;�E�۱E�#�B���C�/�g�3��T0 k� N����%�0d  851t"Q ��    �����EO�|>ӡI����W��ߒ!�;�E�ӲE��B���C��o�3��T0 k� ����%�0d  851t"Q ��    �����EO||>ϢI����W��ߓ|;�E�ϳE��B���C��s�3��T0 k� ����%�0d  851t"Q ��    �����EOt|>ˣI����W��ۓ|;�E�ǳEn�B���C��w�3��T0 k� ����%�0d  851t"Q ��    �����EOl{>ˣI����W��۔|;�E�ôEn�E���C��{�3��T0 k� ����%�0d  851t"Q ��    �����EOd{>ǤI����W��ە|;�EEm��E���C���3��T0 k� ����%�0d  851t"Q ��    �����EOTz.ǤI����W��ו|;�EEm��E���C����3��T0 k� /���%�0d  851t"Q ��    �����EOLz.ǤI����W��ז|;�I���E���E���C����3��T0 k� /���%�0d  851t"Q ��    �����EODz.ǥI����W��Ӗ|;�I���E���E���C����3��T0 k� /���%�0d  851t"Q ��    �����EO<y.ǦI����W��Ӗ|;�I���E���E���C�۰��3��T0 k� /���%�0d  851t"Q  ��    �����EO8y.˧I����W��ϖ|;�I���E���E���C�ӱ��3��T0 k� /���%�0d  851t"Q  -�    �����EO0x.˨I����W��ϗ|;�I���E���E���C�˱��3��T0 k� ����%�0d  851t"Q  ��    �����E? w.˪I����W��˗|;�I���E���E���C�.��3��T0 k� ����%�0d  851t"Q  ��    �����E?w.ϪI����W��Ǘ|;�IΛ�E���E���C�.��3��T0 k� ����%�0d  851t"Q  ��    �����E?vϫI����W��Ǘ|;�IΛ�E���E���C�.��3��T0 k� ����%�0d  851t"Q ��    �����E?vӬI����S��×|;�IΛ�E���E���C�.��3��T0 k� ?��#�%�0d  851t"Q ��    �����E?uӭI����S����|;�IΗ�E���E���C�.��3��T0 k� ?��#�%�0d  851t"Q ��    �����E>�t׮I����S����|;�IΗ�F��E���D����3��T0 k� ?#��'�%�0d  851t"Q ��    �����E>�s߯I����S����|;�I���F��E���D����3��T0 k� ?#��'�%�0d  851t"Q ��    �����E>�r��I����L ���|;�I���F��E���D���3��T0 k� �'��+�%�0d  851t"Q ��    �����E>�q��I����H��|;�I���F� E���Dw���3��T0 k� �#��'�%�0d  851t"Q ��    �����E>�p��I����H��|;�I���F�E.��I�o���3��T0 k� �'��+�%�0d  851t"Q ��    �����E.�o���I����H��|;�IΏ�F�E.��I�g���3��T0 k� �'��+�%�0d  851t"Q ��    �����E.�n���I����H��|;�IΏ�F�E.��I�c���3��T0 k� �+��/�%�0d  851t"Q ��    �����E.�m /�I���mD��|;�IΏ�D݄E/�I�[���3��T0 k� /;��?�%�0d  851t"Q ��    �����E.�k /�A���mD��|;�IΏ�D݄E/�I�K���3��T0 k� /O��S�%�0d  851t"Q ��    �����E.�j /�A���mDm��|;�I���D݄E/�I�C�ø3��T0 k� /[��_�%�0d  851t"Q  ��    �����E.�h /�A���m@m��|;�I���D݄	E/�I�;�Ǹ3��T0 k� /c��g�%�0d  851t"Q  ��    �����E.�g /#�A���}@m��|;�I���D݀
E/#�I�3�˹3��T0 k� �o��s�%�0d  851t"Q  ��    �����E.�f /'�A���}@	m��|;�I���D݀E/'�I�+�Ϻ3��T0 k� �{���%�0d  851t"Q  ��    �����E.�e //�A���}@
m�|;�I���D݀E/+�I�#�Ӻ3��T0 k� ������%�0d  851t"Q  /�    �����E.�d /7�A���}<m{�|;�E^��F|E3�C��׻3��T0 k� ������%�0d  851t"Q  ��    �����E.�c ??�A���}<ms�|;�E^��F|E7�C��׼3��T0 k� ������%�0d  851t"Q  ��    �����E.�a ??�A���}<mo�|;�E^��F|E7�C��ۼ3��T0 k� O�����%�0d  851t"Q  �    �����E�_ ?O�BM���8mg�|;�E^��F|EC�C����3��T0 k� O�����%�0d  851t"Q  ��    �����E�^ ?W�BM���8m_�|;�E^��F|EG�C����3��T0 k� O�����%�0d  851t"Q  ��    �����E�] ?c�BM���4m[�|;�EN��F|EO�C���3��T0 k� OǷ�˷%�0d  851t"Q  ��    �����E�[ ?k�BM���4}W�|;�EN��F|EW�C���3��T0 k� �Ϸ�ӷ%�0d  851t"Q  ��    �����E�Z ?s�BM���4}O�|;�EN��F|E[�C�߱��3��T0 k� �׶�۶%�0d  851t"Q  ��    �����B��Y ?{�B����0}K�|;�EN�F|!B�c�C�ױ��3��T0 k� �߶��%�0d  851t"Q  ��    �����B��X ?��B����0}G�|;�EN{�E�|#B�k�C�ϱ���3��T0 k� ����%�0d  851t"Q  ��    �����B��W ?��B����,}?�|;�C�{�E�|%B�o�E�Ǳ���3��T0 k� �����%�0d  851t"Q  ��    �����B��V O��B����,};�|;�C�w�E��&B�w�E࿱���3��T0 k� ������%�0d  851t"Q  ��    �����B��U O��B����(}7�|;�C�s�E��(B��Eෲ��3��T0 k� �����%�0d  851t"Q  ��    �����B��T O��B����(}3�|;�C�o�E��*B���E௲��3��T0 k� ����%�0d  851t"Q  ��    �����B��S O��B����(}/�|;�C�o�E��,B���E৲��3��T0 k� ����%�0d  851t"Q  ��    �����B�|R O��B����$}'�|;�C�k�E��.B���E�����3��T0 k� ����%�0d  851t"Q  �    �����E�|Q��B����$�#�|;�C�g�E��/@��E��� �3��T0 k� ����%�0d  851t"Q  �    �����E�|PǷB����$��|;�C�c�E��1@��E��� �3��T0 k� ����%�0d  851t"Q  ��    �����E��N׶B���� !��|;�C�[�E��4@��E��� #�3��T0 k� ����%�0d  851t"Q  ��    �����E��M߶B���� "��|;�C�[�@�6@��A�{� '�3��T0 k� ����%�0d  851t"Q  ��    �����E��KO�B���� #��|;�C�W�@�8@��A�s� +�3��T0 k� ����%�0d  851t"Q  ��    �����E��JO�B���� $��|;�C�S�@�9@��A�o� /�3��T0 k� ����%�0d  851t"Q  ��    �����E��IO��B���� $��|;�C�O�@�;@��A�g� 3�3��T0 k� �#��'�%�0d  851t"Q  ��    �����E��HO��B���� %��|;�ENG�@�<@��A�_� 7�3��T0 k� �+��/�%�0d  851t"Q  ��    �����E��G@�B���� &��|;�ENC�@�>@��A�W� ;�3��T0 k� �/��3�%�0d  851t"Q  ��    �����E��E0�B���� &��|;�EN?�@�?@��I�S� ?�3��T0 k� �7��;�%�0d  851t"Q  ��    �����E��D0�B���� '��|;�EN;�@�A@��I�S� C�3��T0 k� �;��?�%�0d  851t"Q  �    �����E��C0�E���� '��|;�EN7�@�B@��I�S� G�3��T0 k� �;��?�%�0d  851t"Q  ��    �����E��A0�E���� '��|;�EN3�@�D@��I�S� K�3��T0 k� �;��?�%�0d  851t"Q  ��    �����CN�@0�E����$(��|;�EN/�@�E@��I�S� O�3��T0 k� �;��?�%�0d  851t"Q  ��    �����CN�?0�E����$(���|;�A+�@�G@��J�S� S�3��T0 k� �;��?�%�0d  851t"Q  ��    �����CN�=0�E����$(���|;�A'�@�H@��J�S� W�3��T0 k� �;��?�%�0d  851t"Q  ��    �����CN�<@�E����$(���|;�A#�@�I@�J�S� [�3��T0 k� �;��?�%�0d  851t"Q  ��    �����CN�:@�E����()���|;�A�@�K@�J�S� _�3��T0 k� �;��?�%�0d  851t"Q  ��    �����CN�8@�E���()���|;�A�@�L@�J�S� c�3��T0 k� �;��?�%�0d  851t"Q  ��    �����CN�7@�E���,)���|;�A�@�M@�J�W� c�3��T0 k� �;��?�%�0d  851t"Q  ��    �����CN�5@�E���,)���|;�A�@�O@�J�W� g�3��T0 k� �K��O�%�0d  851t"Q �    �����C^�4P�E���0)���|;�A�@�P@�J�W� k�3��T0 k� �[��_�%�0d  851t"Q ��    �����C^�2P�E���0)��|;�A�@�Q@#�APW� o�3��T0 k� �g��k�%�0d  851t"Q ��    �����C^�0P�B���4)��|;�A�@�R@+�APW� s�3��T0 k� �w��{�%�0d  851t"Q ��    �����C^�/P�B�#��4)��|;�A�@�S@/�APW� w�3��T0 k� ������%�0d  851t"Q ��    �����C^�-P�B�'��8)��|;�A�@�U@3�APW� w�3��T0 k� ����%�0d  851t"Q ��    �����E.�+`�B�/��<(��|;�A�@�V@7�APW� {�3��T0 k� ����%�0d  851t"Q ��    �����E.�)`�B�3��<(��|;�A��@�W@;�A�W� �3��T0 k� ����%�0d  851t"Q ��    �����E.�(`�B�7��@(��|;�A��@�X@;�A�W� ��3��T0 k� �÷�Ƿ%�0d  851t"Q ��    �����E.�&`�B�?��D(��|;�A��@�Y@?�A�[� ��3��T0 k� �ϸ�Ӹ%�0d  851t"Q	 ��    �����E.�$`�B�C��D'��|;�A��@�Z@C�A�[� ��3��T0 k� �߹��%�0d  851t"Q
 ��    �����E.�"`�B�K��H'��|;�A��@�[@G�A�[� ��3��T0 k� ����%�0d  851t"Q ��    �����E.� `�B�O��L&��|;�A��@�\@K�A�[� ��3��T0 k� ������%�0d  851t"Q ��    �����B��`�CW�P&��|;�A��@�]@O�A�[� ��3��T0 k� ����%�0d  851t"Q ��    �����B��`�C[�T&��|;�A��@�^@O�A�[� ��3��T0 k� ����%�0d  851t"Q ��    �����B��`�Cc�X%��|;�A��@�_@S�A�[� ��3��T0 k� �'��+�%�0d  851t"Q ��    �����B��`�Cg�\%��|;�A�@�`@W�A�[� ��3��T0 k� �7��;�%�0d  851t"Q ��    �����B��`�Co�`$��|;�A�@�a@[�A�[� ��3��T0 k� �G��K�%�0d  851t"Q ��    �����B��`�Cs�d#��|;�A߿@�b@_�A�_� ��3��T0 k� �S��W�%�0d  851t"Q ��    �����B��`�C{�h#�߸|;�A۾@�c@c�A�_� ��3��T0 k� �c��g�%�0d  851t"Q ��   �����B��`�C�l"�߸|;�A۾@�d@g�A�[� ��3��T0 k� �s��w�%�0d  851t"Q ��    �����B��`�C��p!�߸|;�A׾@�e@k�A�[� ��3��T0 k� �����%�0d  851t"Q ��    �����B��`�C��t!�߹|;�AӾ@�f@k�E`[� ��3��T0 k� �����%�0d  851t"Q ��    �����B��`�C��x �۹|;�Aӽ@�g@o�E`[� ��3��T0 k� �����%�0d  851t"Q ��    �����B��`�C���|�۹|;�AϽ@�h@s�E`[� ��3��T0 k� �����%�0d  851t"Q ��    �����C�	`�C��݀�۹|;�AϽ@�h@w�E`[� ��3��T0 k� �����%�0d  851t"Q ��    �����C�`�C��݄�ۺ|;�A˽@�i@{�E`W� ��3��T0 k� ������%�0d  851t"Q ��    �����C� �C��݈�׺|;�AǼ@�j@{�EPW� ��3��T0 k� ������%�0d  851t"Q ��    �����C� �C��ݐ�׺|;�AǼ@�k@�EPS� ��3��T0 k� ������%�0d  851t"Q ��    �����C� �C��ݔ�׻|;�Aü@�l@��EPS� ��3��T0 k� ������%�0d  851t"Q ��    �����C�  �C��ݘ�׻|;�Aü@�m@��EPO� ��3��T0 k� ����%�0d  851t"Q ��   �����C�� �C��ݜ�ӻ|;�A��@�m@��EPO� ��3��T0 k� ����%�0d  851t"Q ��    �����C�� �C��ݤ�ӻ|;�A��@�n@��C�K� ��3��T0 k� �#��'�%�0d  851t"Q ��    �����C�� �C��ݨ�Ӽ|;�A��@�o@��C�K� ��3��T0 k� �3��7�%�0d  851t"Q ��    �����C�� �C��ݬ�Ӽ|;�A��@�p@��C�G� ��3��T0 k� �?��C�%�0d  851t"Q ��    �����C�� �C.��ݰ�Ӽ|;�A��@�p@��C�C� ��3��T0 k� �O��S�%�0d  851t"Q ��    �����C�� �C.����ϼ|;�A��@�q@��C�?� ��3��T0 k� �_��c�%�0d  851t"Q ��    �����C�� �C.����Ͻ|;�A��@�r@��C�;� ��3��T0 k� �k��o�%�0d  851t"Q ��    �����C�� �C.�����Ͻ|;�A��@�r@��AP;� ��3��T0 k� �{���%�0d  851t"Q ��    �����C�� �C.�����Ͻ|;�A��@�s@��AP7� ��3��T0 k� �����%�0d  851t"Q ��    �����C�� #�E����Ͻ|;�A��@�t@��AP3� ��3��T0 k� �����%�0d  851t"Q ��    �����C�� #�E����Ͼ|;�A��@�t@��AP/� ��3��T0 k� �����%�0d  851t"Q ��    �����C� #�E����˾|;�A��@�u@��AP+� ��3��T0 k� �����%�0d  851t"Q ��    �����C� #�E����˾|;�A��@�v@��AP+� ��3��T0 k� ������%�0d  851t"Q ��    �����C� #�E'����˾|;�A��@�v@��AP'� ��3��T0 k� ������%�0d  851t"Q ��    �����C� #�E+���	�˿|;�A��@�w@��AP#� ��3��T0 k� ������%�0d  851t"Q ��    �����C� #�E3����˿|;�A��@�x@��AP� ��3��T0 k� ������%�0d  851t"Q ��    �����C/� #�E;����˿|;�A��@�x@��AP� ��3��T0 k� �����%�0d  851t"Q ��    �����C/� #�EC����ǿ|;�A��@�y@��AP� ��3��T0 k� ����%�0d  851t"Q ��    �����C/� #�B�K���ǿ|;�A��@�y@��AP� ��3��T0 k� ���#�%�0d  851t"Q ��    �����C/#� #�B�S�����|;�A��@�z@��AP� ��3��T0 k� �+��/�%�0d  851t"Q ��    �����C/'� #�B�[�����|;�A��@�{@��AP� ��3��T0 k� �;��?�%�0d  851t"Q ��    �����K�+� #�B�c�����|;�A��@�{@��AP� ��3��T0 k� �K��O�%�0d  851t"Q ��    �����K�/� #�B�k������|;�A��@�|@��AP� ��3��T0 k� �W��[�%�0d  851t"Q ��    �����K�3� '�Io��#����|;�A��@�|@��AP� ��3��T0 k� �g��k�%�0d  851t"Q ��    �����K�7� '�Iw��+����|;�A��@�}@��AP� ��3��T0 k� �w��{�%�0d  851t"Q ��   �����K�7� '�I{��/����|;�A��@�}@��AP� ��3��T0 k� �����%�0d  851t"Q ��    �����K�;� '�I���7����|;�A��@�~@��AP� ��3��T0 k� �����%�0d  851t"Q ��    �����K�?� '�I��;����|;�A��@�~@��AP� ��3��T0 k� �����%�0d  851t"Q ��    �����K�C� '�I/��?����|;�A��@�@��A_�� ��3��T0 k� �����%�0d  851t"Q ��    �����K�G� '�I/��G����|;�A��@�@��A_�� ��3��T0 k� �����%�0d  851t"Q ��    �����K�K� '�I/��K����|;�A��@�@��A_�� ��3��T0 k� �� �� %�0d  851t"Q ��    �����K�O� '�I/��S����|;�A��@�@��A_�� ��3��T0 k� ����%�0d  851t"Q $�    �����K�O� '�I/��~W����|;�A��@�@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�S� '�I��~[����|;�A��@�@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�W� '�I��~c����|;�A��@�@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�[� '�I��~g����|;�A��@�@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�_� '�I��~k����|;�A��@�~@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�_� '�I��~s����|;�A��@�~@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�c� '�I/��~w����|;�A��@�~@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�g� '�I/��~{����|;�A��@�~@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�k� '�I/��~����|;�A�@�}@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�k� +�I/��~�����|;�A�@�}@��A_�� ��3��T0 k� ����%�0d  851t"Q $�    �����K�o� +�I/ê������|;�A�@�}@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�s� +�Iê������|;�A�@�}@��A_�� ��3��T0 k� ����%�0d  851t"Q ��    �����K�s� +�IǪ������|;�A{�@�}@��A_�� ��3��T0 k� �� �� %�0d  851t"Q ��    �����K�w� +�IǪ������|;�A{�@�|@��A_�� ��3��T0 k� ������%�0d  851t"Q ��    �����K�{� +�I˪�����|;�A{�@�|@��A_�� ��3��T0 k� ������%�0d  851t"Q ��    �����K�{� +�I˪�����|;�Aw�@�|@��A_�� ��3��T0 k� �����%�0d  851t"Q ��    �����K�� +�I/Ϫ�����|;�Aw�@�|@��A_�� ��3��T0 k� �����%�0d  851t"Q ��    �����Kσ� +�I/Ϫ�����|;�Aw�@�|@��A_�� �3��T0 k� �����%�0d  851t"Q ��    �����Kσ� +�I/Ϫ�����|;�Aw�@�{@��A_�� �3��T0 k� �����%�0d  851t"Q ��    �����Kχ� +�I/Ϫ�����|;�As�@�{@��A_�� �3��T0 k� �����%�0d  851t"Q ��    �����Kχ� +�I/Ϫ����#�|;�As�@�{@��A_�� �3��T0 k� �����%�0d  851t"Q ��    �����Kϋ� +�IӪ����'�|;�As�@�{@��A_�� �3��T0 k� �����%�0d  851t"Q ��    �����KϏ� +�IӪ����/�|;�As�@�{@��A_�� �"���T0 k� �����%�0d  851t"Q ��    �����KϏ� +�IӪ����3�|;�As�@�{@��A_�� �"���T0 k� �����%�0d  851t"Q ��    �����Kϓ� +�IӪ����7�|;�Ao�@�z@��A_�� �"���T0 k� �����%�0d  851t"Q ��    �����Kϓ� +�IӪ����?�|;�Ao�@�z@��A_�� �"���T0 k� �����%�0d  851t"Q
 ��    �����Kϓ��+�@Ӫ����G�|;�Ao�@�z@��A_�� �"���T0 k� �����%�0d  851t"Q
 ��    �����Kϓ��+�@Ӫ����K�|;�Ao�@�z@��A_�� �"���T0 k� �����%�0d  851t"Q	 ��    �����Kϓ��+�@ת����S�|;�Ao�@�z@��A_�� �"���T0 k� �����%�0d  851t"Q	 ��    �����Kϓ��+�@ת����W�|;�Ak�@�z@��A_�� �"���T0 k� �����%�0d  851t"Q ��    �����Kϓ��+�@ת����_�|;�Ak�@�y@��A_�� �"���T0 k� ӿ����%�0d  851t"Q ��    �����Kϗ��+�K�ת����g�|;�Ak�@�y@��A_�� �"���T0 k� ӿ����%�0d  851t"Q ��    �����Kϗ��/�K�ת����o�|;�Ak�@�y@��A_�� �"���T0 k� ӿ����%�0d  851t"Q ��    �����Kϗ��/�K�۪����s�|;�Ak�@�y@��A_�� �3��T0 k� ӿ����%�0d  851t"Q ��    �����Kϗ��/�K�۪����{�|;�Ag�@�y@��A_�� �3��T0 k� ӿ����%�0d  851t"Q ��    �����Kϗ��/�K�۪������|;�Ag�@�y@��A_�� �3��T0 k� ������%�0d  851t"Q ��    �����Kϗ��/�K�۪������|;�Ag�@�y@�A_�� �3��T0 k� ������%�0d  851t"Q ��    �����Kϛ��/�K�۪������|;�Ag�@�x@�A_�� �3��T0 k� ������%�0d  851t"Q ��    �����Kϛ��/�K�ߪ������|;�Ag�@�x@�A_�� �3��T0 k� ������%�0d  851t"Q ��    �����Kϛ��/�K�ߪ������|;�Ac�@�x@�A_�� �3��T0 k� ������%�0d  851t"Q ��    �����Kϛ��/�K�ߪ������|;�Ac�@�x@�A_�� �3��T0 k� ӿ����%�0d  851t"Q ��    �����Kϛ��/�K�ߪ������|;�Ac�@�x@�A_�� �3��T0 k� ӿ����%�0d  851t"Q  ��    �����K����/�K�ߪ������|;�Ac�@�x@�A_�� �3��T0 k� ӿ����%�0d  851t"Q  ,�    �����K����/�K�������|;�Ac�@�x@�A_�� �3��T0 k� ӿ����%�0d  851t"Q  ��    �����K����/�K�������|;�Ac�@�w@�A_�� �"s��T0 k� ӿ����%�0d  851t"Q  ��    �����K����/�K�������|;�A_�@�w@�A_�� �"s��T0 k� �����%�0d  851t"Q ��    �����K����/�K�������|;�A_�@�w@�A_�� �"s��T0 k� �����%�0d  851t"Q ��    �����K����/�K�������!�;�A_�@�w@�A_�� �"s��T0 k� �����%�0d  851t"Q ��    �����B����/�K�������!�;�A_�@�w@�A_�� �"s��T0 k� �����%�0d  851t"Q ��    �����B����/�K�������!�;�A_�@�w@�A_�� �"s��T0 k� �����%�0d  851t"Q ��   �����B����/�K�������!�;�A_�@�w@�A_�� �"s��T0 k� �����%�0d  851t"Q ��    �����B����/�K�����!�;�A_�@�w@�A_�� �"s��T0 k� �����%�0d  851t"Q ��    �����B����/�K�����!�;�A[�@�w@�A_�� �"s��T0 k� �����%�0d  851t"Q ��    �����E/���/�K�����!�;�A[�@�v@�A_�� �"s��T0 k� �����%�0d  851t"Q ��    �����E/�� /�K�����!�;�A[�@�v@�A_�� �"s��T0 k� �����%�0d  851t"Q ��    �����E/�� /�K����'�!�;�A[�@�v@�A_�� �3��T0 k� ÿ����%�0d  851t"Q ��    �����E/�� /�K��#��/�!�;�A[�@ v@�A_�� �3��T0 k� ÿ����%�0d  851t"Q ��    �����E/�� /�K���'��7�!�;�A[�@ v@�A_�� �3��T0 k� ÿ����%�0d  851t"Q ��    �����E�� /�K���'��?�|;�A[�@ v@�A_�� �3��T0 k� ÿ����%�0d  851t"Q ��    �����E�� /�K���+��G�|;�A[�@ v@�A_�� �3��T0 k� ÿ����%�0d  851t"Q ��    �����E�� /�K���/��O�|;�AW�@ v@�A_�� �3��T0 k� ������%�0d  851t"Q ��    �����E�� /�K���3��_�|;�AW�@ v@�A_�� #�3��T0 k� ������%�0d  851t"Q ��    �����E��� /�K���7��k�|;�AW�@ v@�A_�� #�3��T0 k� ������%�0d  851t"Q ��    �����E��� /�K���;��s�|;�AW�@ u@�A_�� #�3��T0 k� ������%�0d  851t"Q ��    �����E�Ô 3�K���?��{�|;�AW�@ u@�A_�� #�3��T0 k� ӿ����%�0d  851t"Q ��    �����E�ǔ 3�K���?����|;�AW�@ u@�A_�� #�3��T0 k� ӿ����%�0d  851t"Q ��    �����E�˔ 3�K���C����|;�AW�@ u@�A_�� #�3��T0 k� ӿ����%�0d  851t"Q ��    �����E�ϓ 3�K���G����|;�AW�@ u@�A_�� #�3��T0 k� ӿ����%�0d  851t"Q ��    �����Eӓ 3�K���K����!�;�AS�@ u@�A_�� #�3��T0 k� ӿ����%�0d  851t"Q ��    �����Eӓ 3�K���O����!�;�AS�@ u@�A_�� '�3��T0 k� �����%�0d  851t"Q ��    �����Eד 3�K���S����!�;�AS�@ u@�A_�� '�3��T0 k� �����%�0d  851t"Q ��    �����Eۓ 3�K���W�޳�!�;�AS�@ u@�A_�� '�3��T0 k� �����%�0d  851t"Q  ��    �����Eߓ 3�K���[�޿�!�;�AS�@u@�A_�� '�3��T0 k� �����%�0d  851t"Q  ��    �����E� 3�K���_����!�;�AS�@u@�A_�� '�3��T0 k� �����%�0d  851t"Q  .�    �����E� 3�K���c����!�;�AS�@u@�A_�� '�3��T0 k� �����%�0d  851t"Q  ��    �����Eo� 3�K����g����!�;�AS�@t@�A_�� '�3��T0 k� �����%�0d  851t"Q  ��    �����Eo� 3�K����g����!�;�AS�@t@�A_�� '�3��T0 k� �����%�0d  851t"Q  ��    �����Eo� 3�K����k����!�;�AS�@t@�A_�� '�3��T0 k� �����%�0d  851t"Q  ��    �����Eo� 3�K����o����!�;�AO�@t@#�A_�� '�3��T0 k� �����%�0d  851t"Q  ��    �����Eo� 3�K����o����|;�AO�@t@#�A_�� +�3��T0 k� ÿ����%�0d  851t"Q  ��    �����D?� 3�K����s����|;�AO�@t@#�A_�� +�3��T0 k� ÿ����%�0d  851t"Q  ��    �����D?�� 3�K����w���|;�AO�@t@#�A_�� +�3��T0 k� ÿ����%�0d  851t"Q  ��    �����D?�� 3�K����w���|;�AO�@t@#�A_�� +�3��T0 k� ÿ����%�0d  851t"Q  ��    �����D?�� 3�K����w���|;�AO�@t@#�A_�� +�3��T0 k� ÿ����%�0d  851t"Q  ��    �����D?�� 3�K����{���|;�AO�@t@#�A_�� +�3��T0 k� ������%�0d  851t"Q  ��    �����Eo�� 3�K����{��'�|;�AO�@t@#�A_�� +�3��T0 k� ������%�0d  851t"Q  ��    �����Eo�� 3�K����{��/�|;�AO�@t@'�A_�� +�3��T0 k� ������%�0d  851t"Q  ��   �����Eo�� 3�K������7�|;�AO�@t@'�A_�� +�3��T0 k� ������%�0d  851t"Q  ��    �����Eo�� 7�K�����?�|;�AO�@t@'�A_�� +�3��T0 k� ������%�0d  851t"Q  ��    �����Eo�� 7�K�����G�|;�AO�@t@'�A_�� +�3��T0 k� ������%�0d  851t"Q  ��    �����E_�� 7�K����O�|;�AO�@t@'�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����E_�� 7�@���O�|;�AK�@t@'�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����E_�� 7�@����S�|;�AK�@s@'�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����E_�� ;�@����W�|;�AK�@s@'�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����E_�� ;�@����_�|;�AK�@s@'�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����E�� ;�@����_�|;�AK�@s@+�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����E�� ;�J����_�|;�AK�@s@+�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����E�� ;�J����c�|;�AK�@s@+�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����E�� ;�J�����c�|;�AK�@s@+�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����E� ?�J�����g�|;�AK�@s@+�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����Ko� ?�J�����k�|;�AK�@s@+�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����Ko� ?�J�����o�|;�AK�@s@+�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����Ko� ?�J����s�|;�AK�@s@+�A_�� /�3��T0 k� ������%�0d  851t"Q  ��    �����Ko� ?�J����s�|;�AK�@s@+�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����Ko� ?�J����w�|;�AK�@s@+�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����E� ?�J����{�|;�AK�@s@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����E� C�J����{�|;�AG�@s@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����E� C�J�O���{�|;�AG�@s@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����E� C�J/�O����|;�AG�@s@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����E� C�J/�O�����|;�AG�@s@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����Eߙ C�J/�O�����|;�AG�@s@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����E/ߙ C�J/�O�����|;�AG�@s@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����E/ۙ C�J/�O�����|;�AG�@s@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����E/י G�J/ߪO�����|;�AG�@s@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����E/י G�J/ߪO�����|;�AG�@s@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����E/ә G�J/ߪO�����|;�AG�@r@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����K�ϙ G�J/ߪO�����|;�AG�@r@/�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����K�˙ G�J/ߪO�����|;�AG�@r@3�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����K�˙ G�J/ߪO�����|;�AG�@r@3�A_�� 3�3��T0 k� ������%�0d  851t"Q  ��    �����K�Ǚ G�J۪O�����|;�AG�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����K�Ù G�J۪ �����|;�AG�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����K�Ù K�J۪ �����|;�AG�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����K��� K�J۪ �����|;�AG�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����K��� K�J۪ �����|;�AG�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����K��� K�Jת �����|;�AG�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����K��� K�Jת �����|;�AG�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����K��� K�Jת �����|;�AG�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����K��� K�JӪ �����|;�AG�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����K��� K�JӪ �����|;�AG�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����Kϫ� K�JϪ �����|;�AC�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����Kϫ� O�J?Ϫ �����|;�AC�@r@3�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����Kϧ� O�J?Ϫ �����|;�AC�@r@7�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����Kϧ� O�J?Ϫ �����|;�AC�@r@7�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����Kϣ� O�J?˪ �����|;�AC�@r@7�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����Kϣ� O�J?˪ �����|;�AC�@r@7�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��   �����Kϟ� O�J?˪ �����|;�AC�@r@7�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����Kϛ� O�J?˪ �����|;�AC�@r@7�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����Kϛ� O�J?˪ �����|;�AC�@r@7�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����Kϗ� O�J?˪ �����|;�AC�@r@7�A_�� 7�3��T0 k� ������%�0d  851t"Q  ��    �����Kϗ� O�J?˪ ����|;�AC�@r@7�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��   �����Kϓ� O�J?˪ ����|;�AC�@r@7�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����Kϓ��S�J˪ ����|;�AC�@r@7�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����KϏ��S�J˪ ��ÿ|;�AC�@r@7�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����KϏ��S�J˪���ÿ|;�AC�@r@7�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����Kϋ��S�J˪���ÿ|;�AC�@r@7�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����Kϋ��S�J˪����ǿ|;�AC�@r@7�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����Kϋ��S�J˪����ǿ|;�AC�@r@7�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����Kχ��S�J˪����˿|;�AC�@r@7�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����Kχ��S�J˪����˿|;�AC�@r@7�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����Kσ��S�J˪����Ͽ|;�AC�@r@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����Kσ��S�J˪���Ͼ|;�AC�@r@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K���S�J˪���Ӿ|;�AC�@r@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K���S�J˪���Ӿ|;�AC�@r@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K���W�J˪���׽|;�AC�@r@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�{��W�J˪���׽|;�AC�@r@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�{��W�J˪���ۼ|;�AC�@r@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�w��W�J˪���oۼ|;�AC�@r@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�w��W�J˪���oۻ|;�AC�@r@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�w��W�J˪���o߻|;�AC�@q@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�s��W�J˪���oߺ|;�AC�@q@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�s��W�J˪���oߺ|;�AC�@q@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�o��W�J˪���o�|;�AC�@q@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�o��W�J˪���o�|;�AC�@q@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�o��W�J˪���o�|;�AC�@q@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�k��W�J˩���o�|;�AC�@q@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�k��W�J˩���?�|;�AC�@q@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�k��W�J˩���?�|;�AC�@q@;�A_�� ;�3��T0 k� ������%�0d  851t"Q  ��    �����K�g��W�J˩���?�|;�AC�@q@;�A_�� ?�3��T0 k� ������%�0d  851t"Q  ��    �����K�g��[�J˩���?�|;�AC�@q@;�A_�� ?�3��T0 k� ������%�0d  851t"Q  ��    �����DD`��Q�/��dG�|C�D��A�E��E3��ᯚc��T0 k� ����%�0d  851t"Q  ��    ��� =DD\��Q�+��`C�|C�D��A�E��E3��ᣚc��T0 k� �ץ�ۥ%�0d  851t"Q  ��G    ��� :DDX��Q�+��\?�|C�D��A�E��E3��ᛙc��T0 k� �ϥ�ӥ%�0d  851t"Q  ��G    ��� 7DTT���U2+��\7�|C�D��A��E��IS��ᓙc��T0 k� �å�ǥ%�0d  851t"Q  ��G    ��� 4DTL���U2'��X/�|C�D��A�E�{�IS����c��T0 k� ����%�0d  851t"Q  ��G    ��� 1DTH���U2'��T'�|C�D��A�E�w�IS���w�c��T0 k� ����%�0d  851t"Q  ��G    ��� .DTD���U2'��P#�|C�D��A׷D�s�IS��k�c��T0 k� ����%�0d  851t"Q  ��G    ��� +DT@���U2#�0L�|C�D{�A϶D�s�Ic{�1c�c��T0 k� ����%�0d  851t"Q  ��G    ��� (DT8 �ÿU2#�0L�|C�Ds�A!öD�o�Ics�1[�c��T0 k� ����%�0d  851t"Q  ��G    ��� %DT4!㻿U2#�0H�|C�Dk�A!��D�h Ico�1O�c��T0 k� ����%�0d  851t"Q  ��G    ��� "DT0"㳾U2�0D�|C�Dc�A!��D�dIck�1G�c��T0 k� �����%�0d  851t"Q  ��G    ��� DT,#㫽U2�0@�|C�D[�A!��I�dIcg�1?�c��T0 k� �w��{�%�0d  851t"Q  ��G    ��� DT($㟼@��0<���|C�DS�A!��I�`E3c�13�c��T0 k� �k��o�%�0d  851t"Q  ��G    ��� Dd'㟼@��04���|C�C�C�A!��I�\E3W�1#�c��T0 k� �W��[�%�0d  851t"Q  ��G    ��� Dd(�@��00 ���|C�C�;�A!��I�\
E3S�1�3��T0 k� �O��S�%�0d  851t"Q  ��G    ��� Dd)�@��0, ���|C�C�3�A!w�I�XE3O�1�3��T0 k� �G��K�%�0d  851t"Q  ��G    ��� Dd+�E��0+����|C�C�+�E�o�I�XE3G�1�3��T0 k� �?��C�%�0d  851t"Q  ��G    ��� Dd,�E��P'����|C�C�'�E�g�I�TE3C�0��3��T0 k� �;��?�%�0d  851t"Q  ��G    ��� 
Ed-�{�E��P#����|C�C��E�[�I�TE3?�@��3��T0 k� �3��7�%�0d  851t"Q  ��G    ��� Ec�/�s�E��P����|C�C��E�S�I�TE#;�@�3��T0 k� �+��/�%�0d  851t"Q  ��G    ��� Ec�1�c�E��P�з�|C�C��E�?�I�PE#3�@ی3��T0 k� ����%�0d  851t"Q  ��G    ��� Ec�3�[�E��P���|C�C���E�7�I�PE#/�@Ӌ3��T0 k� ����%�0d  851t"Q  ��G    �����ES�4�[�E��P���|C�C���E�/�I�PE#+�@Ǌ3��T0 k� ����%�0d  851t"Q  ��G    �����ES�5�[�E��P����|C�C��E�#�I�PE#'�@��3��T0 k� ������%�0d  851t"Q  ��G    �����ES�7S�E��_�����|C�C��E��I�PE##�@��3��T0 k� �����%�0d  851t"Q  ��G    �����ES�8K�E��_���� |C�C�߯E��I�PE#�@��3��T0 k� ����%�0d  851t"Q  ��G    �����ES�9K�E������� |C�C�ׯE��I�PE#�@��3��T0 k� �߯��%�0d  851t"Q  ��G    �����C��:C�C�������| |C�C�ϯE���I�PE#�@��3��T0 k� �ׯ�ۯ%�0d  851t"Q  ��G    �����C��;?�C�������t|C�C�ǯE��I�PE�P��3��T0 k� �Ϯ�Ӯ%�0d  851t"Q  ��G    �����C�>/�C�������d|C�C�E��I�PE�P��3��T0 k� ����%�0d  851t"Q  ��G    �����C�?'�C�������\|C�C�E�׮I�PE�Pw�3��T0 k� ����%�0d  851t"Q  ��G    �����C�@�C�������T|C�C�E�ϮI�LE�Po�3��T0 k� ����%�0d  851t"Q  ��G    �����C�A�C�������L|C�C�E�ǮI�LE��g�3��T0 k� ����%�0d  851t"Q  ��G    �����C�B�C�������@|C�C�E໮I�LE��_�3��T0 k� ����%�0d  851t"Q  ��G    �����C�C�C������8|C�D��E೭EaL E��S�3��T0 k� ������%�0d  851t"Q  ��G    �����C�D�C������0|C�D��EP��EaL!E��K�3��T0 k� ������%�0d  851t"Q  ��G    �����C�E��C������(|C�D�EP��EaH"E��C�3��T0 k� �����%�0d  851t"Q  ��G    �����C�G�C������� |C�Dw�EP��EaH"E��;�3��T0 k� �s��w�%�0d  851t"Q  ��G    �����C�xH�C������� |C�Do�EP��EaD#E���3�3��T0 k� �k��o�%�0d  851t"Q  ��G    �����C�pI�C������� |C�Dg�EP��EQD$E���+�3��T0 k� �_��c�%�0d  851t"Q  ��G    �����C�lJߣC������� |C�D_�EPw�EQ@%E���#�3��T0 k� �W��[�%�0d  851t"Q  ��G    �����C�dJעC�������|C�DW�EPo�EQ@&E����3��T0 k� �K��O�%�0d  851t"Q  ��G    �����C�\KϠC�������|C�DO�EPg�EQ<'E����3��T0 k� �C��G�%�0d  851t"Q  ��G    �����C�XLǟC���w����|C�DG�E@[�EQ8(E����3��T0 k� �;��?�%�0d  851t"Q  ��G    �����C�PM��C���o����|C�D?�E@S�C�8)E���3��T0 k� �/��3�%�0d  851t"Q  ��G    �����C�HNⷝC���g����|C�D7�E@K�C�4)E����3��T0 k� �'��+�%�0d  851t"Q  ��G    �����C�@O⯜D���_����|C�D/�E@?�C�0*E����3��T0 k� ���#�%�0d  851t"Q  ��G    �����C�<P⫛D���[����|C�D+�E@7�C�,+E���3��T0 k� ����%�0d  851t"Q  ��G    �����D4Q⣚D��S����|C�D#�E@/�C�(,E���3��T0 k� ����%�0d  851t"Q  ��G    �����D,R⛙D��K����|C�D�E@'�C�$,E���3��T0 k� ����%�0d  851t"Q  ��G    �����D$SⓘD��C����|C�D�E@�C� -E��ۊ3��T0 k� ������%�0d  851t"Q  ��G    �����DS⋗D��;����|C�D�A �C�.E��׋3��T0 k� �����%�0d  851t"Q  ��G    �����DT⃖D�3����|C�D�A �C�/E��ϋ"s��T0 k� ����%�0d  851t"Q  ��G    �����DU�{�Dw��+����|C�D��A �C�/E��ǋ"s��T0 k� ����%�0d  851t"Q  ��G    �����DV�s�Ds��#����|C�D�A��C�0E��Ë"s��T0 k� �ۗ�ߗ%�0d  851t"Q  ��G    �����D W�o�Dk������|C�D�A��C�1E�ﻌ"s��T0 k� �ӗ�ח%�0d  851t"Q  ��G    �����D�W�g�Dc������|C�C��EO�C�2E�﷌"s��T0 k� �˖�ϖ%�0d  851t"Q  ��G 	   �����D�X�_�D[���o��|C�C�۲EO�EQ 2E߳﯌"s��T0 k� �Õ�Ǖ%�0d  851t"Q  ��G 	   �����D�Y�W�DW���o��|?�C�ӲEOۧEP�3E߲頻"s��T0 k� ������%�0d  851t"Q  ��G 	   �����D�Z�O�DO����o��|?�C�˲EOӧEP�4E߲"s��T0 k� ������%�0d  851t"Q  ��G 	   �����D�Z�G�DG����o��|?�C�òEO˦EP�4E۲"s��T0 k� ������%�0d  851t"Q  ��G 	   �����D�[�?�D?�>��o�|?�CỲEOæEP�5E۱"s��T0 k� ������%�0d  851t"Q  ��G 	   �����D�\�3�D/�>��os�|?�C᫲EO��EP�6Eױ"s��T0 k� ������%�0d  851t"Q  ��G 	   �����D�]�+�D'�>��ok�|?�CᣲEO��E@�7Eױ3��T0 k� ������%�0d  851t"Q  $�G 	   �����D�^�#�D�>��og�|?�CᛲEO��E@�7Eװ3��T0 k� ���%�0d  851t"Q  ��G 	   �����D�^��D�>��o_�|?�CᓲE?��E@�8B�Ӱ��3��T0 k� ���%�0d  851t"Q  ��G 	   �����D�_��D�>��_W�|?�CዲE?��E@�8B�Ӱ�w�3��T0 k� �����%�0d  851t"Q  ��G 	   �����D�`�C��>��_S�|?�C�E?��E@�8B�ӯ�s�3��T0 k� �{���%�0d  851t"Q  ��G 
   �����D�`�C���>��_K�|?�C�{�E?�E@�9B�ӯ�o�3��T0 k� �s��w�%�0d  851t"Q  ��G 
   �����C�a��C���>��_C�|?�C�s�E?w�E@�9B�ӯ�g�3��T0 k� �k��o�%�0d  851t"Q  ��G 
   �����C�b��C���>��_;�|?�C�k�E?w�E@�9B�ӯ�c�3��T0 k� �g��k�%�0d  851t"Q  ��G 
   �����C�b�C���>��_3�|?�C�c�E?o�E@�9B�Ӯ�_�3��T0 k� �c��g�%�0d  851t"Q  ��G 
   �����C�|c�C���N���+�|?�C�[�E?g�E@�9B�Ӯ�_�3��T0 k� �[��_�%�0d  851t"Q  ��G 
   �����C�ldׁC���N����|?�C�K�E?[�C��9JBӮ�W�3��T0 k� �O��S�%�0d  851t"Q  ��G 
   �����C�deρC���N����|?�C�C�E?S�C��9JB׭�O�"���T0 k� �G��K�%�0d  851t"Q  ��G 
   �����C�\eǁC��N{���|;�C�;�E/S�C�|9JB׭�K�"���T0 k� �K��O�%�0d  851t"Q  $�G 
   �����C�Tf��C��^s����;�C�3�E/S�C�t9JB׭�G�"���T0 k� �O��S�%�0d  851t"Q  ��G 
   �����C�Lf��C��^o����;�D/�E/O�C�p9JB׭�?�"���T0 k� �O��S�%�0d  851t"Q  ��G 
   �����C�Dg��C��^g�����;�D'�E/K�C�h9JB׬�;�"���T0 k� �O��S�%�0d  851t"Q  ��G 
   �����C�@g��C��^_�����;�D�E/C�C�`8JB׬�7�"���T0 k� �K��O�%�0d  851t"Q  ��G    �����C�8h��C��^W�����;�D�E/?�C�X8JB׬�3�"���T0 k� �G��K�%�0d  851t"Q  ��G    �����C�0h��C���~S����|;�D�E/;�C�P8JB׬�+�"���T0 k� �C��G�%�0d  851t"Q  ��G    �����C�(i��C��~K����|;�D�E/7�C�H8JB۬�'�"���T0 k� �?��C�%�0d  851t"Q  ��G    �����C� i��C�w�~C����|;�D ��E/7�C�@7JB۫�#�"���T0 k� �?��C�%�0d  851t"Q  ��G    �����C�j{�C�o�~?����|;�D ��E/3�C�87JB۫��"���T0 k� �;��?�%�0d  851t"Q  ��G    �����C�js�C�g�~7����|;�D �E//�C�06JB۫��3��T0 k� �7��;�%�0d  851t"Q  ��G    �����C�kk�C�_�~3����|;�D �E+�C�(6JB۫��3��T0 k� �3��7�%�0d  851t"Q  ��G    �����C� kc�C�W�~+����|;�D ߴE'�C� 5JB۫��3��T0 k� �/��3�%�0d  851t"Q  ��G    �����C��l�W�C�K�~'����|;�D״E'�C�5JB۪��3��T0 k� �/��3�%�0d  851t"Q  ��G    �����C��l�O�D C�~����|;�DϴE#�C�4JB۪��3��T0 k� �+��/�%�0d  851t"Q  ��G    �����C��m�G�D ;������|;�DǴE�C�3JB۪��3��T0 k� �'��+�%�0d  851t"Q  ��G    �����D�m�?�D 3������|;�D��E�C� 3JBߪ���3��T0 k� �'��+�%�0d  851t"Q  ��G    �����D�n�/�D #������|;�D��E��C��1JBߪ>��3��T0 k� �'��+�%�0d  851t"Q  ��G    �����D�n�'�D ������|;�D��E��C��1JBߪ>�3��T0 k� �+��/�%�0d  851t"Q  ��G    �����D�o��D �������|;�D��E��C��0JBߩ>�3��T0 k� �'��+�%�0d  851t"Q  ��G    �����D�o��D �������|;�D��E��C��/JBߩ>�3��T0 k� �'��+�%�0d  851t"Q  ��G    �����                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \���2 ]�">"= 0 ����|�  � �
	   ��ٖ�    ��u����     d�$   
          g����          ���     ���   0
% 
          ���   � �
	    � �    ��� �]     Y �               �����          n�  �  ���   0
 	         ��s"  � �        ��	�    ������%�    ����           $
	����          �
`     ���   8

          ��6   � �
     ��$    ��6��$                       	����           _�    ���   8         ���   C C     .���     ��ll���K    �: �   	            ����          � �     ���  P
		         ���i  ��	      B�r    ���i�r                             ���l              �  ���    P             ��8�       V�P�    ��9�P
�    ����                
  � 8         ��     ��B    
8

            q�x         j����     q�d���.    �� B                ���          �p  �  ��@   0
          �Ԗ*        ~ N�*    �ԓ N�#     / �             
      @�               ��@   0          ��ma        ���z�    ��L���la    � �                    �         	 �0     ��@   8	'	           ��I�          � g    ��Ee �     B v                    :         
  ��     ��@   0
         ���J ��
	      � ���    ���J ���                                �              A  ��H   		 5              �2  ��      �b�      �2b�                                                               �                               ��        ���          ��                                                                 �                         ����  ��        � ���    ���� ���         "                  x                j  �       �                         ��    ��        � �      ��   �           "                                                �                         �� ��������P�� N��  ��� � �  
         	      
     n4� ���B       (� `e� )D  f� �� _` � _� �$  _� �$  _����J ����X � 
�\ V  
�| W� 
�� W� 
�\ W����. ����< ����J ����X � Hd n` H� n� 
�� V� 
�\ W  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0� ���� � � }`���� ����� � 
�\ V� 
�� V� 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ������������   ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"     
�j,� B �
� �  �  
� ��   ��     � �      ����  ��     �       ��   ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  � 5 5      ��  �  ���        �8 �  ��        �        ��        �        ��        �    ��     G�� _��        ��                         �$ ( ! ���                                    �                ����           �� ����%��  ���� 
 F � $          11 Evgeny Davydov      1:57                                                                        1  1     � �
�+ �J� � � J� � � J� � �J� � � J� � � J� � �C � �	C  � �
C$ � �k� � k� �K � �C. � �C4 � �c� �B� � �B� � � B� � � B� � �B� � qk~ �"� � � "� � �"� � �*� � � "  | � "J � "  |8!� |`  "O �@ "2 |` !"@ |` ": �` ": �` ": �`  "O �@&"2 |` ": � � ("J �)"  |`  "K �X  "K �& ,"G �^  "P �[  "P �	  "P � �0"* |  "P � 2"G �>  "P � � 4"F � �5" � �6!� |  "E � � 8"G � � 9"P � � :"F � �;" � �<!� |
  "E � �>!� |  "E �                                                                                                                                                                                                                         |� R        �     @ 
        �     V P E d  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��    �^R�� ��������������������������������������������������������   �4, R� @'�@6��@[�Y                                                                                                                                                                                                                                                                                                                                                 @X�                                                                                                                                                                                                                                         
    N    /    ��   D�J    	  �  	                           ������������������������������������������������������                                                                                                                                       �     '      �        �        � F?          	  
 	 
 	 	 ��������� ������������ ������������ ���� ������� ��������������������� ����� ���������������������� ����� �����  ��� � � ��� ���������������������������������� �� ������������������� ��� ��� ���� ��� ����������  �������������                                   ,     ��  K
�J                                     ������������������������������������������������������                                                                        	                                                           	       �      �              ��      ��             	 	 
  	 
 
 ����� �������������������� ��������������� ���� ���� �������� �� ������������������ ������� ������������������ ������������������������������������ ��������������� �� � �� ������  ������� ����� ������ ��������������������� ��������             F                                                                                                                                                                                                                                                  
                                                             �             


             �  }�                                                                   '�     '�               ����������������  '|����������������������������   &    ������������     '�����������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" % K ?               	                  � � � �\        �c�b7.P�1sc$                                                                                                                                                                                                                                                           ��  	n                                      m            l                                                                                                                                                                                                                                                                                                                                                                                                        	( �  (�  
(�  (�   `  EZmm ������)��p �N G��8����� p��d�j��d�t����2j        6  ���� %��         	 �   & AG� �   �   
           	A\�                                                                                                                                                                                                                                                                                                                                        B F   �     
   
      "         !��                                                                                                                                                                                                                        Y��   �� �� �      �� A 	     ��������� ������������ ������������ ���� ������� ��������������������� ����� ���������������������� ����� �����  ��� � � ��� ���������������������������������� �� ������������������� ��� ��� ���� ��� ����������  ������������� ����� �������������������� ��������������� ���� ���� �������� �� ������������������ ������� ������������������ ������������������������������������ ��������������� �� � �� ������  ������� ����� ������ ��������������������� ��������      �     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    @      <     ��                       B     �   �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ��[�  �    � �$ ^$    ����  �}  ޢ  ��  �1   �    >     �f ��        p���� ��   p���� �$      ���l�����D�������� J  ��  �h       � �N ^$   �   ;���    �z � �N ^$    ;  ��             2�           � ��� �� � ��� �$  � �#��#  �      �   d   ����� e�����  g���        f ^�         �� !��      �      �������2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  " ! " "" """ "!   " ""                                                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "! ""! " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  " ! " "" """ "!   " ""                                                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                       "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��             �  �˰ ��� �wp ���                                                                                                                                                                         �  �  �   �        �� +  �"/��"/����� � ��       ""� "/� ��                      ݼ w|
�wz����������˹�������̽��� ��� ��� ��� I��
D��T33�TCDDTCDET0DED0DDD0��K���  ̘  ��        �  ઠ ઌ ��̐��٠�ˊ��������н�"� ""� "J�  J�  J�  U�  U�  EP  L�  ɀ ��  �� �+" �                                                  �� �� ��               �  �  �     �   �  �  �                ��� �  ��     �                                    �  �� �                         ����     �   �  �  �  ��  �   �                           ��   ��                  �  �  �� � ���                                       �   �   �   �   w  �� ɪ�̚��ə���̚���ɭ�̼��̻��̻���+���(�� H� �C3 UC3
TDCTD0�C 	�� 
�� ���� ���"/� ��   ���   ��  ��  ��  w�  wp  ��� ��� ��̰��̀�͹���ڀ��ذ��� �̰ �̰ ̸� ��� ��3 333�3330�C3: TD3�C��ݸ�	��  ����̲����"/����                  /   /�  �          �      	  *  ,  +   "   � ��  ��  �                            �   �    �   �       �   �   �                .  �   �  ���� �   �             �   ��  ��  ��  �  �   ��  ��                            ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                   ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .      �����                       ���� �                                                                                                                                                                                        ̰ ˻����wݩk}�gz� w�� �  �  � ^� UNMTNL�DB,��2"ʪ����� � �" ""/ ���    �    �   ��  ��  ��� ��� ��� ��� ���0۹�0؊�3���3˻�3���C��X��U��T�����  ��  �   �  "��" �"                  �"  ��  ��  �                                         �   �   ��  ��  ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����            �����                         �     �                                                                                                                                                                                          �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �      �  �  �  �  �  �   �                                                                                                                                                                                                                                                                                 �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �   �� ��� ��                      "   "   "  �� ��                   ����������                                ��  ��  ���  �  �  �   �   ��  �                            �   ���                            �   �                                                                                                    �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   ��  ��  ��  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ��� ���                                                                                                                                                                                              �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �              "      �           �  �   �   ��  �                                        ��  ����   �       �                                   �    ���  ��                    ��  ��  ���                         ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �      �  �                         	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                       �  ��  ��  ww  ��  vv  w"   "   "  �� ��                   ����������                                �    � �  ��                  ���                                                                                                                                                                            �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �              "      �           �  �   �   ��  �            ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                                                                                                                                                                                                                                        �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��    ��    �                              �   �  �  �   �               �   �                               � ����ݼ� ����                                                                                                                                                                             �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""���������������������""""������II������""""������IIII""""������DI�I�""""������DI�I�""""�����IIDIIIA""""��������DD""""������IADD�A��""""��������I���I�������I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ADA�LL��L�D����3333DDDD x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(XxLL����������D����3333DDDD w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""����������A������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(""""�������I�I������ �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�""""�������I��D���I������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`�D�M�D���M������3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(MD�M�A�����MD�����3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(�""""�����AMAD������ � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(�""""������������������ � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
�+ �J� � � J� � � J� � �J� � � J� � � J� � �C � �	C  � �
C$ � �k� � k� �K � �C. � �C4 � �c� �B� � �B� � � B� � � B� � �B� � qk~ �"� � � "� � �"� � �*� � � "  | � "J � "  |8!� |`  "O �@ "2 |` !"@ |` ": �` ": �` ": �`  "O �@&"2 |` ": � � ("J �)"  |`  "K �X  "K �& ,"G �^  "P �[  "P �	  "P � �0"* |  "P � 2"G �>  "P � � 4"F � �5" � �6!� |  "E � � 8"G � � 9"P � � :"F � �;" � �<!� |
  "E � �>!� |  "E �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.�������������������������������������������/�\�M�K�T�_��.�G�\�_�J�U�\� � � � � � �@�9�1�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������@�9�1� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            