GST@�                                                           ~      �       	                                         ��              a         ��  � j� ��         ���    ����        �     %    ����                                d0<|    � �?     uC� ��.�̈�ff"                                                                                                                                                   ����������������������������������������������������������������������������������������������������������������������������������������                               �����                                                                                   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                         �   @  &   �   �                                                                                 'w w                             �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� ��   �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    � � �  �  �                                            ^L��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ���  ��.   ����ff"                                                                                                                                                                                                                                ��                                                                                                              ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �E6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �  � �  �  ��  �  ��  �  ��  �  ��  �  ��  ������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �� �'   Cu  ` � �'   ��  ` �j     � ��     � �$ ^h                  a         �� � �j ��        ���   ` � z�  w                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �                            ����                            ����                            ����                            ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   � � � � � � � ��    �                                                                                   �   �   �   �   �   �   �   ��  �  �  �  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   � � � � � � � �                �     ������  � � � �   �� ���      � �   �� ��  ��� �    �� �� �� �� ��  ��  �� ��������  �  �  �  �  �  �  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �   �                        ��������   ���  � �� �  ��          �    �   �  �� �� �� ��  ���  �  � �� �  �                      �����  ��         ����                        ��������������   �           � � � � �� �� �� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������������
        �  �          �  �  �  ��  ��  ��  ��  ��         �  �  �  �  �  ���������                                    �   �   �   �   �� �� �� �� �� �� �� �� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������  � � � � � � �  � �          ��  ��  �� �� �� �� ��  ���  �  �  �  �  �  �  �  ����       �  �  ����    ��  ��   �                            �   � ��������������������� �� �� �� �� �� �� �� �                       �  �  �   �   �             �   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         � ������  ��  �     �       ��     ����
�      �  ��  �   �   �        �   � ��  �  �        �   �   �  �   �   �                � ��� ��  ��                                       ���  ��  �  �             � �� �� �  �  �  �  �  �          �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �  �  �  � � ��
 ��  ��  �� �� �� �� �� �� �� �� �� ��������������        ���������     ��  �� �� �� �� �� ������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ��  ��  ��  ��  ��� ��� �����       �         ����������� �� ��� �� �� �� �� ��  ���������������������������������� � �     �� �������������������������������������������� �� �� �� �� �� �� �� �����������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���        ��� � �����    ��� ��  �                        ���������    ������� ������  ��������������   ������ ����� ����     ����    ���� ��������� ������� ��������� ���������������������    �� ���������    ���� �������    ������������  ���  ��� �  �������  ��� � ���������     ����������    ������������    �   �����           ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��������� � �    �  �      ����� �       �  �  ��  ��  ��  ��  ����� ��  �� �� �� �� �� ���� �� � �� �     �  �  � �    � � � � ����������    � � ��� �  �   �   �  �  ��  ��  ��  �  �� �� �� �� �� �� �� �� ���������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������������������������������������   �      �  �  ����������������� ��  �   �   �   �   �  �  � �� � � � � � �       �  ��  ��  ��  �   � ��� � 
��
����� �����   ��  ��  �  �  �  �   �   � � � � � � �      ����������������                              �                            �                ��  ������ ��  �  �                              �                       �   �  �                     �   �                                                                                                                                                                                                                                                                                                                                               �����������������  �  �        � � �� ��������������q�q ������ ��� ��� ��� ��       �q     � ��     ��   �   �        ��   �   � �� �� �� ���������quW  �         �  ��U ��U��UU�UUU�           ��� UUU UUU U�U U�U   � U UX UX �UX UZ��U� �U� � ����  ��  ��� � U � U�U�U          �  U  �U UU Z� X       �U� UU� UUP UUP U�P ��P                                                                                                                                                                                                                                                                                                                                                                                                                                                     ���������                ����������������            ��������������������          ����������������� ���       �   �   �   Z   U  UU �UU�   �   � ��� ��� �  ��   �  �  ����� ��� ��� ��� ��� ���  �X �ZX UUP UUP UUPUUP
UU UU   �       �  �  ��  �� �  ��         ����������������                ����������������   �           ���������������������      �   �������������������������  ��  ��������������������� �        �������� ��� ����               ��� ���������  �                   �   ����������������           �  �������� �������      �  U� U� U� �Z U� �UX�UUPUUUPUUU UUU �UP �U� UX        �  � �  �  ��  ��    ��Z�UZ�UUUX UUP UZ  UP �Z �Z UUUUUUUU UU UUU �UZ U� U�U� UU UUUUUU� UZ� UZ��U���U���UU��UU��UU��XU������������X��� �� ��Z�U�U�U�U�U U�Z UUP UU  �UP �UP �UP �UX �UX �U�  U�� U��                 �   �  U  �Z                                                                                                                                                                                                                                                                                                                                                                                                  ����������� ��� ��� ��� �� ��������������������������������������������������������������������  ��  �   �   �  �  
   U  U UZZU���U� UZU UXU U�U U�X UUX   �  � �� �� �� �� ��� ������ ���������������������������� UX       ��������������������   ��  �� ��� ��  ��  ��� ��� ���             �� ����� �   �         � ������������ �   �   �      � ��� � �  �   �  U�  U������������� �� �   �P  �P  ��� ��  � � �� ��  ��   �  � �    UU UUU UUXUUXUUUUU��UZ��U    U   U   U   �   �P  UP  UP  �������������� ��� ��� ��� �����������������������������  ��   �ZP UX  U�  U�  U�  U� U� U�                           � U�� U�� U�� U�� U�� U�� U�� UZ �U �U �U �U  U �U �U ����� ��� ��P �ZP �X� ��  ��  ��U���U���U���U�U�U�U�U�U U�X UXX����U��Z��P��P�P� ��U ��UUU  UU  UZ  ZP  ZP X� �  �   UX� UP� UX��UZ���Z���UU�UX�UX
X  ��  U   U   X   �                                                                                                                                                                                                                                                                                                                                                                                                             ��  �  �   �   �   �      ��������������������������������������� ��� ��� ��� ��� ��������  
U  �U UU UU �UU �U   �   UUX UUX UU� UU� UU� UU  UU  UU   ��� ��� ��� ��� ��� ���������������������������� ��� ��� ��  �   ��� ���� ��         UP  UX  ��  ����������  ��  �  � �   �  U  U  �U U� 
U� UUU UUU�  �U  �X �X ��P � P� P� P�  U  UU UUU UUU UUUUUUUUUUUUUUP  �P  �P  �P  �P  �P  ��  ��  �   U  U U U U� U� U� U�������������������������UU�UUXU�  U   �P  �P  U   U      �   � ��� ��� ��� ����������� ��������  ��  �� �� �� �� ��  ��� U� U� UU UZ UU UU UU UU    �  � �� ��� ��� ��  �   �  �� U � U�  U�  U   U �U�U
�UU �U  �U  UU UU�XU�PUUU UUU �  �X  �   �  �  �  ��  �  �  UZP U�  U�  U�  U�  U� U� ZX  ��U � U � U � U � X � P �  � �  U   U   U                   �UX�    �                                                                                                                                                                                                                                                                                                                                                                                                                                    �  �������� � ��         �   �   ��   �   �   ���������������  ��  ��       ���������������� ��� ������������  �  �   �  �  
�  �  �  UU  UU  UZ  UX  UX  UX  UP  UX  �������������������� ��� ��  �   �  
   U   U  U  UU 
UUUP UP UUP UUP UUP UUP ZU� UU       � �� U� U�U �   �� UUU�UUUX�UX�U� U� 
U� U�  ���������U������������������ �UZ UUUUUU�UU� U�� U��U��UU�UU� �� �� � ��� ��� ��� �   � � U� �U  UX U� U� U� �U� �U�UUUX�UUPUX� U   X  �  �    � �� �� ����  ��    �  U  Z������� ��     X U� U��UU�UU� �   ��  �  ��  �P  �U� �UP �UU UU �UU UZ�UZPUZX
UUUUUU      � ��� UUUUUXUUPUUX UX  ZX������U  ��  �   �   
  �  �UUX UUP UX  U   U   U   �        �  �  �   ��  ��  �   �   UU �UU �UP  U�  U   U  �   �                                                                                                                                                                                                                                                                                                                                                                                                              � �� ��  �     � �        ��� ��� � �� � �  �   �                �   U   U UZ UU ��    �  �U  �U  �U   U  U ��   �   �   �  �  �� U  �U UU �   U� �U� UUP UUP UU� ZU� ZU  ���������� ��� ��� ����������  �  ��  U�  U�  U�  U�  U   UU�  Z�  Z�  X   X  �  �  �  ��� ��� ��� ��  ��  �� ��  ���  �UU UUUU�U�U�UUX�UU� U�  U  UUU� UU  UU� UU� UU� UU� UU�UU� ��� ��� ��� ��� ��� ���������  U�  U� U� U� �U���U��U��U��UP �U �P �P UP �U  �U  �P  ��UU�UU�UU��UU��UU��UU �U� �U�   �  U� ��PUZPUXP�UPUUX UUP ��U�X�UU �UU�UU��UU��U� �UX �UZ�  �  �     �  ���UUUUUUUUUX 
�U X����U �U� �X  U�  �       �UU��UUU UUU  �U  U  X�� ���� U� �U  �U  �X  �P  �   �        UUU UUU UUU U�� U �   ��  ��  U�  U   P                         �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  U  U  U     U �UUUUUUUUUUZ�UXUUU�UUUUP UUX�UUUUUUZ�UUU�UUU�UUUUUUUUU  � � � � � P � P�X����U���X U� �U�UUUUUUUUUUUUUU��UX�UPU �U ��Z � X � �� ��
 ��Z ��X UU UUUUXU�UP�UZ�UZ��U� ��� ��UU� UX  UX  UX  UX  UX  UP  UP  �������� �� ���������������   U   U  U  U  
U  U� �U� �U�  ��  ��  ��  �Z  X  X �X ���� ��������������� �� �  
�    U�  U�  U�  U�� U�� U�� U�� UUU�UU�UU �UU��UU��UU�UU 
UU�������  ��U�� U���U ��Z �UP �UP ��U��UU�UUU�UUU�UZP�UZ��UU��UU�P  �P  ��  �   �   �   �  �  � UU� UUU �UU �UU �UU �UU  U   U UU� UX  U  U  P  �     �   � UU�UU�UU� UU� UZ� U��   �   UUU�UUX U   Z                                   � �� �     ��� ��� ��� ���                                                 ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                UZ U� �UU UZU UZU UXX U� U� UUX UX  Z            �  �� �UUU�UUUUUUUUUUXUUPUU�UU ZU �U��U�  �   �   �   �  �  �  UP UX 
U� U� U� U� U� U����������Z���� ��� ��� �UX �U� ��� �� ��� ��� ��U ��U � U� UUX  UX  UU  UX  UX  UU  UU� UU� ���������  �� 
�  �� U�Z���X �UU�UU� UU�UU�UU�UU�UU�UUZ   U   U   U  �U  �U ZU UU�UUX �P  UP ��� �P  �P  U�  P     �� U� U� U  U  U�  U�  U�  UUU UUUUU�UUUUUPUUUPUUU�UU� UX  U  �U  �X  �           �� �� UU  UU  UP U� X  �   �  ����  �  �  �� �� �� �����������  �   ��� ��������������������  �  � ������������������������� ��� ������������������  �               �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     
         U� �UZ UUU UUU UUU UUU UZU UZU  ��  ��  ��   �  ��  �� �  � ZU �ZU �UU U�U U�X UU� ZX  XP   �  �   �   �   �              U� U� �U� U� U� U� U� �U��U  UU  UP  U   U   U  U  �X  �� U�  U�  U�  U�  U  U  U   UUU�UUPUUXUU�UUU�UUUUUUUUUXUUU�UUX UUP U�  U  X     �   �   �UU�UU�UU�UU UU  UU  U  U�UUXUUU UU  UX  U�  U   �        �  �  �� �� ����  �   �   �  U�  U�  �                   U�  U   X   �     ����������� ��� ����������������������������������������������������������������������������������������������������������������  �   �   ������� ��  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             UZU UUU UU��UU� UU��UU�XUU�ZUU�U � � � U  Z  X  � ��U ��Z �UXZP  ��  �   X  �  ��              �                            �UU �UU UUX UUX UUPUUPUU�UU X  ��                �   �        U   U   �                  UUU UU� UP  UP  U         � �     �  �   �                    U                               �  ���  �                  �                                                               ����  �                        ����������� ���  ��            ������������������� �          ������  �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                UUZUUUUU�UU�UUU UUU UUU UUU UUU UU�UUX UUX UUP UU� U   U   X                                                                   UU Z  X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       UUU UU� �U�  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          	 
                        ! " # $ % & ' (                                                                                                                                                                                 ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P                                                                                                                                                                                 Q R S T U V W X Y Z [ \ ] ^ _ ` a b c d e f g h i j k l m n o p q r s t u v w x                                                                                                                                                                                 y z { | } ~  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �                                                                                                                                                                                 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �                                                                                                                                                                                 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �                                                                                                                                                                                 � � � � � � � � � � � � � � � 	
                                                                                                                                                                                 !"#$%&'()*+,-./0123456789:;<=>?@                                                                                                                                                                                ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefgh                                                                                                                                                                                ijklmnopqrstuvwxyz{|}~�����������������                                                                                                                                                                                ����������������������������������������                                                                                                                                                                                ����������������������������������������                                                                                                                                                                                �������������������������������                                                                                                                                                                                 	
 !"#$%&'()*+,-./0                                                                                                                                                                                123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWX                                                                                                                                                                                YZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�                                                                                                                                                                                ����������������������������������������                                                                                                                                                                                ����������������������������������������                                                                                                                                                                                ����������������������������������������                                                                                                                                                                                ������� 	
                                                                                                                                                                                 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGH                                                                                                                                                                                IJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnop                                                                                                                                                                                qrstuvwxyz{|}~�������������������������                                                                                                                                                                                ����������������������������������������                                                                                                                                                                                ����������������������������������������                                                                                                                                                                                ����������������������� 	
                                                                                                                                                                                 !"#$%&'()*+,-./012345678                                                                                                                                                                                9:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ~      �
u "V  �&      *   "   ����,G       @   @               �           ��ùnS@     @                          ��������    	                                                                                       �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                           ��������    	                                                                                       �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                           ��������    	                                                                                       �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                           ��������    	                                                                                       �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                           ��������    	                                                                                       �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                           ��������    	                                                                                       �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                                            �  >  >                                                                   ����������������������������������������������������������������������������������������������������������������������������������������                               �����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �����   �   �   ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �����   �   �   ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                �jx��jx�g�u��xvf%
 f%
 9l  6                      @           �   @  &   ��7�                            �     �7        `�  �   5               ��              a         ��  � j� ��         ���    ����    � v�         %      @   @                                                 @   @                                                                                                                                                                                                                                                                                                 ��         �                              �  ��.   ����ff"                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �?                       ��               �      �       p� X�                      ��������������������������������������������������������������������������������������������������������������������������������������� �     		

			


   !!""###$$%%%&&' ' ( (!(!)!)"*"*"*#+#+#,$,$-$-%-%.&.&/&/'0'0'0(1(1(2)2)2)3*3*4*4+5+5+5,6,6,7-7-8.8.8.9/9/:/:0:0;0;1<1<1=2=2=2>3>3?3?4?4@4@5A5A6B6B6B7C7C7D8D8E8E9E9F9F:G:G:G;H;H;I<I<J=J=J=K>K>L>L?M?M?M@N@N@OAOAOAPBPBQBQCRCRCRDSDSETETEUFUFUFVGVGWGWHWHXHXIYIYIZJZJZJ[K[K\K\L\L]M]M^M^N_N_N_O`O`OaPaPbPbQbQcQcRdRdRdSeSeSfTfTgUgUgUhVhViViWjWjWjXkXkXlYlYlYmZmZnZn[o[o\o\p\p]q]q]q^r^r^s_s_t_t`t`u`uavavawbwbwbxcxcydydydzeze{e{f|f|f|g}g}g~h~hhii�i�j�j�j�k�k�l�l�l�m�m�m�n�n�n�o�o�o�p�p�p�q�q�q�r�r�r�s�s�t�t�t�u�u�u�v�v�v�w�w�w�x�x�x�y�y�y�z�z�{�{�{�|�|�|�}�}�}�~�~�~����������������������������������������������������������������������������������������������������������������������������������������������������������   d   0   <      |                   �       �   ?                             u   C          uC     ~          �                       ��    ����@M~ �` >���                        