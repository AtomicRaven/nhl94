GST@�                                                            \     �                              	                  ��       �  ��            �������J���ʳ������������������        f     #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    "�j* ,  �����
�"     �j@ �    ��
  Y                                                                               ����������������������������������      ��    oo b go  4  +c  c  'c       ��       	  
    	G 7� V( 	(                 �n 1         8:8�����������������������������������������������������������������������������������������������������������������������������=?  00  45  18                        
     
                ��  �4  �  ��                  nY  	          : �����������������������������������������������������������������������������                                �>  >       Ȳ   @  #   �   �                                                                                '     �1n  	nY    H   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E > �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    A^�O@��_W��`��\|( D�H+A|f �X<��]�\W3� T0 k� �_��c�UHC"!U2d    ��    � ��A^�N@��_W��`��\|( E�H,A|f �X<��]�\W3� T0 k� �_��c�UHC"!U2d    ��    � ��A^�N@��_W��`��\|( E�D,A|f �X<��]�\W3� T0 k� �[��_�UHC"!U2d    ��    � ��A^�N@��_W��`��\|( E�D,A|f �X=��]�`W3� T0 k� �[��_�UHC"!U2d    ��    � ��A^�N@��_W��`��\|( E�D,A|f �X=��]�`W3� T0 k� �W��[�UHC"!U2d    ��    � ��A^�N@��_W��`��\|( E�D-A|f �\=��]�`W3� T0 k� �S��W�UHC"!U2d    ��    � ��A^�N@��_W��`��\|( F@-A|f �\>��]�dW3� T0 k� �S��W�UHC"!U2d    ��    � ��A^�N@��_W��`��\|( F@.A|f �\>��]�dW3� T0 k� �O��S�UHC"!U2d    ��    � ��A^�N@��_W��`��\|( F@.A|f �\>��]�dW3� T0 k� �O��S�UHC"!U2d    ��    � ��A^�N@��_W��`��\|( F@/A|f �\?��]�dW3� T0 k� �K��O�UHC"!U2d    ��    � ��A^�M@��_W��`��\|( F@0A|f �\?��]�dW3� T0 k� �K��O�UHC"!U2d    ��    � ��A^�M@��_W��`��\|( D�@0A|f �\?��]�dW3� T0 k� �G��K�UHC"!U2d    ��    � ��A^�M@��_W��`��\|( D�@0A|f �\@��]�dW3� T0 k� �G��K�UHC"!U2d    ��    � ��A^�M@��_W��`��\|( D�@1A|f �\@��]�dW3� T0 k� �C��G�UHC"!U2d    ��    � ��A^�M@��_W��`��\|( D�@1A|f �\A>�]�dW3� T0 k� �C��G�UHC"!U2d    ��    � ��A^�M@��_W��`��\|( D�@2A|f �\A>�]�dW3� T0 k� �?��C�UHC"!U2d    ��    � ��A^�M@��_W��`��\|( D�@2A|f �`B>�]�dW3� T0 k� �?��C�UHC"!U2d    ��    � ��A^�M@��_W��`��\|( D�@2A|f �`B>�]�dW3� T0 k� �;��?�UHC"!U2d    ��    � ��A^�M@��_W��`��\|( D�@3A|f �`C>�]�dW3� T0 k� �;��?�UHC"!U2d    ��    � ��A^�M@��_W��`��\|( D�D3A|f �`D>�]�dW3� T0 k� �7��;�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�D4A|f �`D>�]�dW3� T0 k� �3��7�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�D5A|f �dE>�]�dV3� T0 k� �3��7�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�D6A|f �dE>�]�dV3� T0 k� �/��3�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�H6A|f �dE>�]�dW3� T0 k� �/��3�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�H6A|f �dEN�]�dW3� T0 k� �+��/�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�H6A|f �dFN�]�dW3� T0 k� �+��/�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�H6A|f �hFN�]�dW3� T0 k� �'��+�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�L7A|f �hGN�]�dW3� T0 k� �'��+�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�L7A|f �hGN�]�dW3� T0 k� �#��'�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�L8A|f �lGN�]�dW3� T0 k� �#��'�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�L8A|f �lGN�]�dW3� T0 k� ���#�UHC"!U2d    ��    � ��A^�L@��_W��`��\|( D�L8A|g �lGN�]�hW3� T0 k� ���#�UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�L8A|g �lGN�]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�L8A|g �lG>�]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�L9A|g �pG>�]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�P9A|g �pG>�]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�P9A|g �pG>�]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�P9A|g �pG>�]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�P9A|g �pG>�]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�P9A|g �pG>�]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�P9A|g �tG>�]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�P9A|g �tG>�]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�P9A|g �tG��]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( D�T9@�|g �tG��]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( ET9@�|g �tG��]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( ET9@�|g �tG��]�hW3� T0 k� ����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( ET9@�|g �xG��]�hW3� T0 k� �����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( ET9@�|g �xG��]�hW3� T0 k� �����UHC"!U2d    ��    � ��A^�K@��_W��`��\|( EX9@�|g�xG��]�hW3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~X9@n�g�xG��]�dW3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~X9@n�h�|G��]�dW3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~X9@n�g�|H��]�dW3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~X9@n�g�|H��]�dW3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~\9@n�gހH��]�dW3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~\9B��gހH��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~\:B��gހI��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~`:B��gބI��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~`:B��gބI��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~`:B��gބJ��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L~d;B��gބJ��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�d;@n�gވJ��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�d;@n�gވJ��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�d;@n�g�J��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�h;@n�g�K��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�h<@n�g�K��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�h<@n�g�K��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�l<K��g�K��]�dX3� T0 k� ������UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�l<K��g�K��]�dX3� T0 k� �׿�ۿUHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�l<K��g�K��]�dX3� T0 k� �׿�ۿUHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�l<K��g�K>�]�dX3� T0 k� �Ӿ�׾UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�p<K��g�K>�]�dX3� T0 k� �ӽ�׽UHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�p<K��g�K>�]�dX3� T0 k� �Ͻ�ӽUHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�p<K��g�K>�]�dX3� T0 k� �ϼ�ӼUHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�p<K��g�K>�]�hX3� T0 k� �˻�ϻUHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�p<K��g�K>�]�hX3� T0 k� �˻�ϻUHC"!U2d    ��    � ��A^�K@��_W��`��\|( L�p<K��h�K>�]�hX3� T0 k� �Ǻ�˺UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�p<K��h�K>�]�hX3� T0 k� �ǹ�˹UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�p<K��h�K>�]�hX3� T0 k� �ù�ǹUHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�p<K��h�K>�]�hX3� T0 k� �ø�ǸUHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�t<K��h�KN�]�hX3� T0 k� �÷�ǷUHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�t<K΀h�KN�]�hX3� T0 k� ����÷UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�t=K΀h�KN�] hX3� T0 k� ����öUHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�t=K΀h�KN�] hX3� T0 k� ������UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�t=K΀h�KN�] hX3� T0 k� ������UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�x=K΄h�LN�] hX3� T0 k� ������UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�x=K΄h�LN�] hX3� T0 k� ������UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�x=K΄i�LN�]�lX3� T0 k� ������UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�x=K΄i�LN�]�lX3� T0 k� ������UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�x=K΄i�L>�]�lX3� T0 k� ������UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�|>K΄i�L>�]�lX3� T0 k� ������UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�|>K΄i�L>�]�lX3� T0 k� ������UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�|>K΄i�L>�]�pX3� T0 k� ������UHC"!U2d    ��    � ��A^�J@��_W��`��\|( L�|>K΄i�L>�]�pX3� T0 k� ������UHC"!U2d    ��    � ��D@@�  c�� ;�k|( E�O�@�D������C3� T0 k� �@�DUHC"!U2d   �� 
   � ��D<@�  _�� :�k|( B�K�@�D������C3� T0 k� �<�@UHC"!U2d   �� 
   � ��D8@�  [�� 8�k|( B�K�@�D�������C3� T0 k� �8�<UHC"!U2d   �    � ��D0@�  W��$7�j|( B�G�@�D�������D3� T0 k� �8�<UHC"!U2d   �    � ��AP,@�  S��$5��j|( B�G�@�D�������D3� T0 k� �4�8UHC"!U2d   ��    � ��AP(@� PO��$4�|j|( B�G�@�D�������D3� T0 k� �0�4UHC"!U2d   ��    � ��AP 	@� PK��$2�xj|( E�C�@�D�������D3� T0 k� �0�4UHC"!U2d   ��    � ��AP	@� PG��$1�pj|( E�C�@�D�������D3� T0 k� �,�0UHC"!U2d   ��    � ��AP	@� PC��$/�hi|( E�C�@�D�������D3� T0 k� �(�,UHC"!U2d   ��    � ��AP	@� P?��(.�di|( E�C�@�D�������D3� T0 k� �$�(UHC"!U2d   ��    � ��AP	@� P;��(-�\i|( E�C�@�D�������D3� T0 k� �� UHC"!U2d   ��    � ��AP	@� P7��(+�Xi|( E~?�A D������D3� T0 k� ��UHC"!U2d   ��    � ��AP
@� P3��(*�Ph|( E~?�A D������D3� T0 k� ��UHC"!U2d   ��    � ��A_�
@� P3��()�Lh|( E~?�A D ������D3� T0 k� ��UHC"!U2d   ��    � ��A_�
@� P/��('�Dh|( E~?�A D ������D3� T0 k� ��UHC"!U2d   ��    � ��A_�
@� P+��,&�@h|( E~?�A D ������D3� T0 k� ��UHC"!U2d   ��    � ��A_�
@� P'��,%�8h|( D�?�APD ������D3� T0 k� ��UHC"!U2d   ��    � ��A_�@��P#��,$�4g|( D�?�APD ������E3� T0 k� ��UHC"!U2d   ��    � ��A_�@��P��,"�0g|( D�;�APD � ����E3� T0 k� � �UHC"!U2d   ��    � ��A_�@��P��,!�(g|( D�;�APD �����E3� T0 k� � �UHC"!U2d   ��    � ��A_�@��P��, �$g|( D�;�APD �����E3� T0 k� � �UHC"!U2d   ��    � ��A_�@��P��,� g|( D�;�APD �����E3� T0 k� � �UHC"!U2d   ��    � ��A_�@��P��0�f|( D�;�A�H ����E3� T0 k� � �UHC"!U2d   ��    � ��A_�@��P��0�f|( D�;�A�D ����E3� T0 k� � �UHC"!U2d   ��    � ��A_�@��P��0�f|( D�;�A�D �	���E3� T0 k� � �UHC"!U2d   ��    � ��A_�@��P��0�f|( D�;�A�D ����E3� T0 k� �� UHC"!U2d   ��    � ��A_�@��P��0�f|( D�;�A�D ����E3� T0 k� �� UHC"!U2d   ��    � ��A_�@��P��0� f|( D�7�D0D ����E3� T0 k� �� UHC"!U2d   �    � ��A_�@��P��4��e|( D�7�D0D ����E3� T0 k� ���UHC"!U2d   ��    � ��A_�@��_���4��e|( D�7�D0D � ���E3� T0 k� ���UHC"!U2d   ��    � ��A_�@��_���8��e|( D�7�D0@ � ���E3� T0 k� �� �� UHC"!U2d    ��    � ��A_�@��_���<��e|( D�7�D0@ �����E3� T0 k� �� �� UHC"!U2d    ��    � ��A_�@��_���<��e|( D�7�D0@ �����E3� T0 k� ��!��!UHC"!U2d    .�   � ��A_�@��_��@��e|( D�7�D0< �����E3� T0 k� ��"��"UHC"!U2d    ��    � ��A_�@��_��@��d|( D�7�D0< �����F3� T0 k� ��"��"UHC"!U2d    ��    � ��A_�@��_��D��d|( D�7�D@< �����F3� T0 k� �#��#UHC"!U2d    ��    � ��A_�@��_��D��d|( D�7�D@8 �����F3� T0 k� �$��$UHC"!U2d    ��    � ��A_�@��_��H��d|( D�7�D@8 �����F3� T0 k� �$��$UHC"!U2d    ��    � ��A_�@��_��H��d|( D�3�D@4 �����F3� T0 k� �%��%UHC"!U2d    ��   � ��A_�@��_��L��d!�( D�3�D@4 �����F"�� T0 k� �&��&UHC"!U2d    ��    � ��A_�@��_��L��d!�( D�3�D@0 �����F"�� T0 k� ��&��&UHC"!U2d    ��    � ��A_�@��_ߓ�P��c!�( D�3�D@, �����F"�� T0 k� ��'��'UHC"!U2d    ��    � ��A_�@��_ߔ�P��c!�( D�3�D@, �����F"�� T0 k� ��'��'UHC"!U2d    ��    � ��A_�@��_۔�T��c!�( D�3�D@(  �����F"�� T0 k� ��(��(UHC"!U2d    ��    � ��A_�@��_۔�T��c!�( D�3�D@$! ����xF"�� T0 k� ��(��(UHC"!U2d    ��    � ��A_�@��_ה�X��c!�( D�3�D@$! ���{�tF"�� T0 k� ��)��)UHC"!U2d    ��   � ��A_�@��_Ӕ�X��c!�( D�3�DP " ���w�pF"�� T0 k� ��*��*UHC"!U2d    ��    � ��A_�@��_Ӕ�\��c!�( D�3�DP# ���s�lF"�� T0 k� ��*��*UHC"!U2d    ��    � ��A_�@��_ϔ�\��c!�( D�3�DP$ ���k�dF"�� T0 k� ��+��+UHC"!U2d    ��    � ��A_�@��_ϔ�\��b!�( D�3�DP$ ���g�`F"�� T0 k� ��+��+UHC"!U2d    ��    � ��A_�@��_˔�`��b|( D�/�DP% ���_�\F3� T0 k� ��,��,UHC"!U2d    ��    � ��A_�@��_˔�`��b|( D�/�DP&���W�XF3� T0 k� ��'��'UHC"!U2d    ��    � ��A_�@��_ǔ�`��b|( D�/�DP'���S�TF3� T0 k� ��%��%UHC"!U2d    ��    � ��A_�@��_ǔ�`��b|( D�/�DP(���K�PF3� T0 k� ��"��"UHC"!U2d    ��    � ��A_�@��_Õ�`��b|( D�/�DP)���C�HF3� T0 k� ��!��!UHC"!U2d    ��    � ��A_�@��_Õ�`��b|( D�/�DP *���?�DF3� T0 k� �� �� UHC"!U2d    ��    � ��A_�@��_Õ�`��b|( D�/�D_�+���7�@G3� T0 k� �� �� UHC"!U2d    ��    � ��A_�@��_���`��b|( D�/�Do�,���/�!<G3� T0 k� ����UHC"!U2d    ��    � ��A_�@��_���`��a|( D�/�Do�-���'�!8G3� T0 k� ����UHC"!U2d    ��    � ��A_�@��_���`��a|( D�/�Do�.���#�!4G3� T0 k� ����UHC"!U2d    ��    � ��A_�@��_���`��a|( D�/�Do�/�� ��!0G3� T0 k� �� �� UHC"!U2d    ��    � ��A_�@��_���`��a!�( D�/�Do�0�� ��!,G"s� T0 k� �� �� UHC"!U2d    ��    � ��A_�@��_���`��a!�( D�/�E_�1�� ��!(G"s� T0 k� �� �� UHC"!U2d    ��    � ��A_�@��_���`��a!�( D�, E_�2޼!R�!$G"s� T0 k� ��!��!UHC"!U2d    ��    � ��A_�@��_���`�|a!�( L^,E_�3޼!Q��! G"s� T0 k� ��!��!UHC"!U2d    ��    � ��A_�@��_���`�xa!�( L^,E_�4�"Q��!G"s� T0 k� ��"��"UHC"!U2d    ��    � ��A_�@��_���`�xa!�( L^(E_�4�"Q��!G"s� T0 k� ��"��"UHC"!U2d    ��    � ��A_�@��_���`�ta!�( L^(E_�5�#Q��!G"s� T0 k� ��#��#UHC"!U2d    ��    � ��A_�@��_���`�p`!�( L^(
E_�6�#Q��!G"s� T0 k� ��#��#UHC"!U2d    ��    � ��A_�@��_���`�p`!�( L^(C��7�#Q��!G"s� T0 k� ��#��#UHC"!U2d    ��    � ��A_�@��_���`�l`!�( L^(C�8�$Q��!G"s� T0 k� ��$��$UHC"!U2d    ��    � ��A_�@��_���`�l`!�( L^(C�9�$Q��!G"s� T0 k� ��$��$UHC"!U2d    ��    � ��A_�@��_���`�h`|( L^(C�:�$A��!G3� T0 k� ��$��$UHC"!U2d    ��    � ��A_�@��_���`�d`|( L^(C�;�%A��! G3� T0 k� ��%��%UHC"!U2d    ��    � ��A_�@��_���`�d`|( L^(C�;�%A��! G3� T0 k� ��%��%UHC"!U2d    ��    � ��A_�@��_���`�``|( L^(C�<�&A�� �G3� T0 k� ��&��&UHC"!U2d    ��    � ��A_�@��_���`�``|( L^(C�=�&A�� �G3� T0 k� ��&��&UHC"!U2d    ��    � ��A_�@��_���`�\`|( L^(C�>�&��� �G3� T0 k� ��&��&UHC"!U2d    ��    � ��A_�@��_���`�\`|( Ln(C�>�'��� �G3� T0 k� ��'��'UHC"!U2d    ��    � ��A_�@��_���`�X`|( Ln(C�?�'��� �G3� T0 k� ��'��'UHC"!U2d    ��    � ��A_�@��_���`�X`|( Ln( C�|@�'�� �G3� T0 k� ��'��'UHC"!U2d    ��    � ��A_�@��_���`�T`|( Ln("C�tA�(�w� �G3� T0 k� ��(��(UHC"!U2d    ��   � ��A_�@��_���`�T_|( Ln($C�lA�(�o� �G3� T0 k� ��(��(UHC"!U2d    ��    � ��A_�@��_���`�P_|( Ln(%C�hB�(�g� �G3� T0 k� ��(��(UHC"!U2d    ��    � ��A_�@��_���`�P_|( Ln('C�`C�(�_� �G3� T0 k� ��(��(UHC"!U2d    ��    � ��A_�@��_���`�L_|( Ln((C�XD�)�W� �G3� T0 k� ��(��(UHC"!U2d    ��    � ��A_�@��_���`�L_|( Ln(*E�PD�)�O� �H3� T0 k� ��(��(UHC"!U2d    ��    � ��A_�@��_���`�H_|( Ln(+E�LE�)�G� �H3� T0 k� ��(��(UHC"!U2d    ��    � ��A_�@��_���`�H_|( Ln(-E�DF�*�?� �H3� T0 k� ��)��)UHC"!U2d    ��    � ��A_�@��_���`�D_|( Ln$.E�<G�*�7� �H3� T0 k� ��)��)UHC"!U2d    ��    � ��A_�@��_���`�D_|( Ln$0E�4H�*�/� �H3� T0 k� ��)��)UHC"!U2d    ��    � ��A_�@��_���`�D_|( Ln$1E�0H�*�'� �H3� T0 k� ��*��*UHC"!U2d    ��    � ��A_�@��_���`�@_|( Ln$3E�(I�+�� �H3� T0 k� ��*��*UHC"!U2d    ��    � ��A_�@��_���`�@_|( Ln$4D? J�+�� �H3� T0 k� ��*��*UHC"!U2d    ��    � ��A_�@��_���`�<_|( Ln$5D?K�+�� �H3� T0 k� ��*��*UHC"!U2d    ��    � ��A_�@��_���`�<_|( Ln$7D?L�,�� �H3� T0 k� ��+��+UHC"!U2d    ��    � ��A_�@��_���`�<_|( Ln$8D?M�,�� �H3� T0 k� ��+��+UHC"!U2d    ��    � ��A_�@��_���`�8_|( Ln$9D?M�,��� �H3� T0 k� ��+��+UHC"!U2d    ��    � ��A_�@��_���`�8_|( Ln$;I� N�,����H3� T0 k� ��+��+UHC"!U2d    ��    � ��A_�@��_���`�4^|( Ln$<I��O�-����H3� T0 k� ��,��,UHC"!U2d    ��    � ��A_�@��_���`�4^|( Ln$=I��O�-����H3� T0 k� ��,��,UHC"!U2d    ��    � ��A_�@��_���`�4^|( Ln$>I��P�-�� �H3� T0 k� ��,��,UHC"!U2d    ��    � ��A_�@��_���`�0^|( Ln$?I��P�-�� �H3� T0 k� ��,��,UHC"!U2d    ��    � ��A_�@��_���`�0^|( Ln$AI��Q�-���H3� T0 k� ��-��-UHC"!U2d    ��    � ��A_�@��_���`�0^|( Ln$BI��Q�.���H3� T0 k� ��-��-UHC"!U2d    ��    � ��A_�@��_���`�,^|( Ln$CI��Q�.���H3� T0 k� ��-��-UHC"!U2d    ��    � ��A_�@��_���`�,^|( Ln$DI��Rސ. ��H3� T0 k� ��-��-UHC"!U2d    ��    � ��A_�@��_���`�,^|( Ln$EI��Rސ. ��H3� T0 k� ��.��.UHC"!U2d    ��    � ��A_�@��_���`�(^|( Ln$FL>�Rތ/ ��H3� T0 k� ��.��.UHC"!U2d    ��    � ��A_�@��_��`�(^|( Ln$GL>�Rތ/ ��H3� T0 k� ��.��.UHC"!U2d    ��    � ��A_�@��_��`�(^|( Ln$HL>�Sތ/ ��H3� T0 k� ��.��.UHC"!U2d    ��    � ��A_�@��_��`�$^|( Ln$IL>�Sތ/ ���H3� T0 k� ��.��.UHC"!U2d    ��    � ��A_�@��_��`�$^|( Ln$JL>�S ��/ ���H3� T0 k� ��3��3UHC"!U2d    ��    � ��A_�@��_��`�$^|( Ln$KL>�S ��0 ���H3� T0 k� ��6��6UHC"!U2d    ��    � ��A_�@��_{��`� ^|( Ln$LL>�T ��0 ���H3� T0 k� �|8��8UHC"!U2d    ��    � ��A_�@��_{��`� ^|( Ln$ML>�T ��0����H3� T0 k� �|:��:UHC"!U2d    ��    � ��A_�@��_{��`� ^|( Ln$NL>�T ��0����H3� T0 k� �|;��;UHC"!U2d    ��    � ��A_�@��_{��`� ^|( Ln$OL>�T ��0�|��H3� T0 k� �|=��=UHC"!U2d    ��    � ��A_�@��_{��`�^|( Ln$PL>�T ��1�t��H3� T0 k� �|>��>UHC"!U2d    ��    � ��A_�@��_{��`�^|( L^$QL>�U ��1�p�|H3� T0 k� �|?��?UHC"!U2d    ��    � ��A_�@��_w��`�^|( L^$RL>�U ��1�l	�xH3� T0 k� �x?�|?UHC"!U2d    ��    � ��A_�@��_w��`�^|( L^$SL>�U ��1�h	�tH3� T0 k� �x?�|?UHC"!U2d    ��    � ��A_�@��_w��`�^|( L^$TLN�U ��1�`
�lH3� T0 k� �x?�|?UHC"!U2d    ��    � ��A_�@��_w��`�^|( L^$ULN�U ��1�\
�hH3� T0 k� �x@�|@UHC"!U2d    ��    � ��A_�@��_w��`�]|( L^$ULN�V ��2�X
�dH3� T0 k� �x@�|@UHC"!U2d    ��    � ��A_�@��_w��`�]|( D�$VLN�V ��2�T�\H3� T0 k� �x@�|@UHC"!U2d    ��    � ��A_�@��_s��`�]|( D�$WLN�V ��2�L�XH3� T0 k� �x@�|@UHC"!U2d    ��    � ��A_�@��_s��`
�]|( D�$XLN�V ��2�H PH3� T0 k� �t@�x@UHC"!U2d    ��    � ��A_�@��_s��`
�]|( D�$YLN�V ��2�D LH3� T0 k� �t@�x@UHC"!U2d    ��    � ��A_�@��_s��`
�]|( D�$ZLN�W ��2�@ DI3� T0 k� �tA�xAUHC"!U2d    ��    � ��A_�@��_s��`
�]|( D�$[LN�W ��3�8 @I3� T0 k� �tA�xAUHC"!U2d    ��    � ��A_�@��_s��`
�]|( D� \LN�W ��3�4 8I3� T0 k� �tA�xAUHC"!U2d    ��    � ��A_�@��_s��`
�]|( D� ^LN�W ��3�0 0I3� T0 k� �tA�xAUHC"!U2d    ��    � ��A_�@��_s��`
�]|( D� _LN�W ��3�, ,I3� T0 k� �tA�xAUHC"!U2d    ��    � ��A_�@��_o��`
�]|( D� `LN�W ��3�( $I3� T0 k� �tA�xAUHC"!U2d    ��    � ��A_�@��_o��`
�]|( D� aLN�X �|3�$ I3� T0 k� �pA�tAUHC"!U2d    ��    � ��A_�@��_o��`
�]|( F cLN�X �|3�  I3� T0 k� �pB�tBUHC"!U2d    ��    � ��A_�@��_o��`
�]|( F$dLN|X �|4  I3� T0 k� �pB�tBUHC"!U2d    ��    � ��A_�@��_o��`
�]|( F$eLN|X �|4 I3� T0 k� �pB�tBUHC"!U2d    ��    � ��A_�@��_o��`
�]|( F$gLNxX �|4  I3� T0 k� �pB�tBUHC"!U2d    ��    � ��A_�@��_o��`
�]|( F$hLNxX �|4 �I3� T0 k� �pB�tBUHC"!U2d    ��    � ��A_�@��_o��`
�]|( F$iLNtY �|4 �I3� T0 k� �pB�tBUHC"!U2d    ��    � ��A_�@��_k��`
�]|( F$kLNtY �|4 �I3� T0 k� �pB�tBUHC"!U2d    ��    � ��A_�@��_k��`
�]|( F(lLNpY �|4  �I3� T0 k� �pC�tCUHC"!U2d    ��    � ��A_�@��_k��`
�]|( F(mLNpY �|4��I3� T0 k� �lC�pCUHC"!U2d    ��    � ��A_�@��_k��`
�]|( F(oLNlY �x5��I3� T0 k� �lC�pCUHC"!U2d    ��    � ��A_�@��_k��`	�]|( E�,pLNlY �x5���I3� T0 k� �lC�pCUHC"!U2d    ��    � ��A_�@��_k��`	�]|( E�,rLNhY �x5���I3� T0 k� �lC�pCUHC"!U2d    ��    � ��A_�@��_k��`	�]|( E�0tLNdZ �x5���I3� T0 k� �lC�pCUHC"!U2d    ��    � ��A_�@��_k��`	� ]|( E�4vLNdZ �x5���I3� T0 k� �lC�pCUHC"!U2d    ��    � ��A_�@��_k��`	� ]|( E�4wLN`Z �x5���I3� T0 k� �lD�pDUHC"!U2d    ��    � ��A_�@��_g��`	� ]|( E�8xLN`Z �x5���I3� T0 k� �lD�pDUHC"!U2d    ��   � ��A_�@��_g��`	� ]|( E�<zLN\Z �x5���I3� T0 k� �lD�pDUHC"!U2d    ��    � ��A_�@��_g��`	� ]|( E�@{LN\Z �x6���I3� T0 k� �lD�pDUHC"!U2d    ��    � ��A_�@��_g��`	� ]|( E�@|LNX[ �x6���I3� T0 k� �hD�lDUHC"!U2d    ��    � ��A_�@��_g��`	��]|( E�D}LNX[ �t6���tI3� T0 k� �hD�lDUHC"!U2d    ��    � ��A_�@��_g��`	��]|( E�HLNT[ �t6���lI3� T0 k� �hD�lDUHC"!U2d    ��    � ��A_�@��_g��`	��]|( E�L�LNT[ �t6���dI3� T0 k� �hD�lDUHC"!U2d    ��    � ��A_� @��_g��`	��]|( E�P�LNT[ �t6���\I3� T0 k� �hD�lDUHC"!U2d    ��    � ��A_� @��_g��`	��]|( E�TLNP[ �t6��OTI3� T0 k� �hD�lDUHC"!U2d    ��    � ��A_� @��_g��`	��]|( E�XLNP[ �t6��OLI3� T0 k� �hE�lEUHC"!U2d    ��    � ��A_�!@��_g��`	��]|( E�\LNL[ �t6��ODI3� T0 k� �hE�lEUHC"!U2d    ��    � ��A_�!@��_c��`	��]|( E�`~L>L[ �t6��O8I3� T0 k� �hE�lEUHC"!U2d    ��    � ��A_�!@��_c��`	��]|( E�d~L>L\ �t7��O0I3� T0 k� �hE�lEUHC"!U2d    ��    � ��A_�!@��_c��`	��]|( E�h}L>H\ �t7��O(J3� T0 k� �hE�lEUHC"!U2d    ��    � ��A_�"@��_c��`	��]|( E�l}L>H\ �t7��O J3� T0 k� �hE�lEUHC"!U2d    ��    � ��A_�"@��_c��`	��]|( E�p|L>D\ �t7��OJ3� T0 k� �hE�lEUHC"!U2d    ��    � ��A_�"@��_c��`	��]|( E�t|L>D\ �t7��OJ3� T0 k� �dE�hEUHC"!U2d    ��    � ��A_�#@��_c��`	��]|( E�x{L>D\ �p7��OK3� T0 k� �dE�hEUHC"!U2d    ��    � ��A_�#@��_c��`	��]|( E�|zL>D\ �p7����K3� T0 k� �dE�hEUHC"!U2d    ��    � ��A_�$@��_c��`	��]|( E��zL>@\ �p7����K3� T0 k� �dE�hEUHC"!U2d    ��   � ��A_�$@��_c��`	��]|( E��yL>@\ �p7����K3� T0 k� �dF�hFUHC"!U2d    ��    � ��A_�$@��_c��`	��]|( KވxL>@\ �p7����L3� T0 k� �dF�hFUHC"!U2d    ��    � ��A_�%@��_c��`	��]|( KތwL>@\�p7����L3� T0 k� �dB�hBUHC"!U2d    ��   � ��A_�%@��_c��`	��]|( KސwL>@\�p8��	~�L3� T0 k� �d?�h?UHC"!U2d    ��    � ��A_�&@��_c��`��]|( KޔvL>@\�p8��	~�L3� T0 k� �d=�h=UHC"!U2d    ��    � ��A_|&@��__��`��]|( KޘuL>@\�p8��	~�L3� T0 k� �d;�h;UHC"!U2d    ��    � ��A_|&@��__��`��\|( KޜtA�@\�p8��	~�L3� T0 k� �d:�h:UHC"!U2d    ��    � ��A_x'@��__��`��\|( KޠtA�@\�p8��	~�L3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_t'@��__��`��\|( KޤsA�@\�p8��	��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_t(@��__��`��\|( KިrA�@\�p8��	��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_p(@��__��`��\|( KެrA�@\�p8��	��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_l)@��__��`��\|( KެqA�@\�p8��	��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_l)@��__��`��\|( KްpA�@\�p8�� 	��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_h*@��__��`��\|( K޴pA�@\�p8��!��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_d*@��__��`��\|( K޸oA�@\�p8��!��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_d*@��__��`��\|( K�oA�@\�l8��!��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_`+@��__��`��\|( K�nA�@\�l8��"��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_\+@��__��`��\|( K��mA�@\�l9Ϙ#��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_\,@��__��`��\|( K��mBN@\�l9ϔ#��L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_X,@��__��`��\|( K��lBN@\�l9ϐ$�|L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_T-@��__��`��\|( K��lBN@\�l9ό%�xL3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_P-@��__��`��\|( K��kBN@\�l9ό&�pL3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_P.@��__��`��\|( K��kBN@\�l9ψ&�lL3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_L.@��__��`��\|( K��j@@\�l9ψ&�hL3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_H/@��_[��`��\|( K��j@@\�l9τ'�dL3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_D/@��_[��`��\|( K��i@@\�l9π(`L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_D0@��_[��`��\|( K��i@@\�l9π)\L3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_@1@��_[��`��\|( K��h@@\�l9�|*XL3� T0 k� �d8�h8UHC"!U2d    ��    � ��A_<1@��_[��`��\|( K��hB�D\�l9�x+TL3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_82@��_[��`��\|( K��gB�D\�l9�t,PL3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_42@��_[��`��\|( K��gB�D\�l9�t,LL3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_43@��_[��`��\|( K��fB�H\�l9�t,LL3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_03@��_[��`��\|( K��fB�H\�l9�p-LL3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_,4@��_[��`��\|( K��eB�H\�l9�l.LL3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_(4@��_[��`��\|( K��eB�H\�l:�h/LL3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_$5@��_[��`��\|( K��dB�H\�l:�d0LL3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_ 5@��_[��`��\|( K��dB�H\�l:�`1LL3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_ 6@��_[��`��\|( K��cB�H\�l:�`1LL3� T0 k� �d9�h9UHC"!U2d    ��    � ��A_6@��_[��`��\|( K��cB�H\�l:�`2LL3� T0 k� �`9�d9UHC"!U2d    ��    � ��A_7@��_[��`��\|( K��cB�H\�l:�\3LL3� T0 k� �`9�d9UHC"!U2d    ��    � ��A_7@��_[��`��\|( K��bB�H\�l:�X4LL3� T0 k� �`9�d9UHC"!U2d    ��    � ��A_8@��_[��`��\|( K��bB�H\�l:�T5LL3� T0 k� �`9�d9UHC"!U2d    ��    � ��A_8@��_[��`��\|( K� aB�H\�h:�P6LL3� T0 k� �`9�d9UHC"!U2d    ��    � ��A_9@��_[��`��\|( K� aB�H\�h:�L7LL3� T0 k� �`9�d9UHC"!U2d    ��    � ��A_9@��_[��`��\|( K�aB�H\�h:�H8LL3� T0 k� �`9�d9UHC"!U2d    ��    � ��A_:@��_[��`��\|( K�`B�H\�h:�D9LL3� T0 k� �`9�d9UHC"!U2d    ��    � ��A_ :@��_[��`��\|( K�`B�H\�h:�@;LL3� T0 k� �`9�d9UHC"!U2d    ��    � ��A^�:@��_[��`��\|( K�`B�H\�h:�<<LL3� T0 k� �`9�d9UHC"!U2d    ��    � ��A^�;@��_[��`��\|( K�_B�H\�h:�8=LL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�;@��_[��`��\|( K�_B�H\�h:�4>LL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�<@��_[��`��\|( K�_B�H\�h:�4>LL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�<@��_[��`��\|( K�^B�H\�h:�0?LL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�=@��_[��`��\|( K�^B�H\�h:�,@LL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�=@��_W��`��\|( K�^B�H\�h:�(ALL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�=@��_W��`��\|( K�]B�H\�h:� CLL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�=@��_W��`��\|( K�]B�H\�h;�DLL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�=@��_W��`��\|( K�]B�H\�h;�ELL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�=@��_W��`��\|( K�\B�H\�h;�GLL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�>@��_W��`��\|( K�\B�H\�h;�HLL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�>@��_W��`��\|( K� \B�H\�h;�ILL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�?@��_W��`��\|( K� [B�H\�h;�JLL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�?@��_W��`��\|( K� [B�H\�h;� LLL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�?@��_W��`��\|( CO$[B�H\�h;��MLL3� T0 k� �`:�d:UHC"!U2d    ��    � ��A^�@@��_W��`��\|( CO$ZB�H\ �h;��NLL3� T0 k� �\>�`>UHC"!U2d    ��    � ��A^�@@��_W��`��\|( CO$ZB�H\ �h;��OLL3� T0 k� �\A�`AUHC"!U2d    ��    � ��A^�@@��_W��`��\|( CO(YB�H\ �h;��PLL3� T0 k� �\C�`CUHC"!U2d    ��    � ��A^�A@��_W��`��\|( CO(YB�H\ �h;��Q�LL3� T0 k� �\E�`EUHC"!U2d    ��    � ��A^�A@��_W��`��\|( CO,XB�H\ �h;��S�LL3� T0 k� �\F�`FUHC"!U2d    ��    � ��A^�A@��_W��`��\|( CO,XB�H\ �h;��T�LL3� T0 k� �\G�`GUHC"!U2d    ��    � ��A^�A@��_W��`��\|( CO,WB�H\ �h;��T�LL3� T0 k� �\H�`HUHC"!U2d    ��    � ��A^�B@��_W��`��\|( CO0VB�H\ �h;	��U�LL3� T0 k� �\I�`IUHC"!U2d    ��    � ��A^�B@��_W��`��\|( CO0VB�H\ �h;	��V�LL3� T0 k� �\I�`IUHC"!U2d    ��    � ��A^�B@��_W��`��\|( CO0UB�H\ �h;	��W�LL3� T0 k� �\I�`IUHC"!U2d    ��    � ��A^�C@��_W��`��\|( E�4TB�H\ �h;	��XNLL3� T0 k� �\I�`IUHC"!U2d    ��    � ��A^�C@��_W��`��\|( E�4SB�H\ �h;	��XNLL3� T0 k� �\J�`JUHC"!U2d    ��    � ��A^�C@��_W��`��\|( E�4RB�H\ �h;	��YNLL3� T0 k� �\J�`JUHC"!U2d    ��    � ��A^�D@��_W��`��\|( E�4QB�H\ �h;	��ZNLL3� T0 k� �\J�`JUHC"!U2d    ��    � ��A^�D@��_W��`��\|( E�8PB�H\ �h;	��ZNLL3� T0 k� �\J�`JUHC"!U2d    ��    � ��A^�D@��_W��`��\|( E�8OB�H\ �h;	��[>LL3� T0 k� �\J�`JUHC"!U2d    ��    � ��A^�D@��_W��`��\|( E�8NB�H\ �h;	��[>LL3� T0 k� �\J�`JUHC"!U2d    ��    � ��A^�E@��_W��`��\|( E�<MB�H\ �h;	��\>LL3� T0 k� �\J�`JUHC"!U2d    ��    � ��A^�E@��_W��`��\!�( E�<LB�L] �h;	��\>LL"s� T0 k� �\J�`JUHC"!U2d    �    � ��A^�E@��_W��`��\!�( E�<KB�L] �h;	��\>HL"s� T0 k� >XI�\IUHC"!U2d    ��    � ��A^�E@��_W��`��\!�( E�<JB�P] �h;	��]>HL"s� T0 k� >TH�XHUHC"!U2d   ��    � ��A^�F@��_W��`��\!�( E�<HB�P] �h;	��].HM"s� T0 k� >TG�XGUHC"!U2d   ��    � ��A^�F@��_W��`��\!�( E�<GB�T] �h;	��].DM"s� T0 k� >PG�TGUHC"!U2d   ��    � ��A^�F@��_W��`��\!�( E�<FB�T] �h;	��].DM"s� T0 k� >PF�TFUHC"!U2d   ��    � ��A^�F@��_W��`��\!�( E�<EB�T] �d;	��].DM"s� T0 k� �LE�PEUHC"!U2d   ��    � ��A^�G@��_W��`��\!�( E�<CB�T^ �d;	��].@M"s� T0 k� �LD�PDUHC"!U2d   ��    � ��A^�G@��_W��`��\!�( E�<BB�T^ �d;	��].@M"s� T0 k� �HC�LCUHC"!U2d   ��    � ��A^�G@��_W��`��\!�( E�<AB�T^ �d;	��]@N"s� T0 k� �HC�LCUHC"!U2d   ��    � ��A^�G@��_W��`��\!�( E�<@B�X^ �d;	��]@N"s� T0 k� �DB�HBUHC"!U2d   ��    � ��A^�H@��_W��`��\|( E�8?E�X^ �d;	��]@N3� T0 k� �@A�DAUHC"!U2d   ��    � ��A^�H@��_W��`��\|( E�8>E�X^ �d;	��]@O3� T0 k� �@@�D@UHC"!U2d  	 ��    � ��A^�H@��_W��`��\|( E�8<E�X^ �d;	��]@O3� T0 k� �<?�@?UHC"!U2d  	 ��    � ��A^�I@��_W��`��\|( E�4;E�X^ �d;�]�@O3� T0 k� �<?�@?UHC"!U2d  
 ��    � ��A^�I@��_W��`��\|( E�4:E�X^ �d;�]�@O3� T0 k� �8>�<>UHC"!U2d   ��    � ��A^�I@��_W��`��\|( E�09E�\^ �d;�]�DO3� T0 k� N8=�<=UHC"!U2d   ��    � ��A^�I@��_W��`��\|( E�08E�\^ �d;�]�DO3� T0 k� N4<�8<UHC"!U2d   ��    � ��A^�I@��_W��`��\|( E�,7E�\^ �d;�]�DO3� T0 k� N0;�4;UHC"!U2d   ��    � ��A^�J@��_W��`��\|( E�,6E�\^ �d;�]�DO3� T0 k� N0;�4;UHC"!U2d   ��    � ��A^�J@��_W��`��\|( E�(5E�\^ �d;�]�DO3� T0 k� N,:�0:UHC"!U2d   ��    � ��A^�J@��_W��`��\|( E�$4K�\^ �`;.�]�DO3� T0 k� .,9�09UHC"!U2d   ��    � ��A^�J@��_W��`��\!�( D?$4K�`^ �`;.�]�DO"�� T0 k� .(8�,8UHC"!U2d   ��    � ��A^�J@��_W��`��\!�( D? 3K�`^ �`;.�]�DO"�� T0 k� .(7�,7UHC"!U2d   ��    � ��A^�J@��_W��`��\!�( D?2K�`_ �`;.�]�HO"�� T0 k� .$7�(7UHC"!U2d   ��    � ��A^�K@��_W��`��\!�( D?2K�d_ �`;.�]�HO"�� T0 k� . 6�$6UHC"!U2d   ��    � ��A^�K@��_W��`��\!�( D?1K�d_ �`;.�]�HO"�� T0 k� > 5�$5UHC"!U2d   ��    � ��A^�K@��_W��`��\!�( D?1K�d_ �`;.�]�HP"�� T0 k� >4� 4UHC"!U2d   ��    � ��A^�K@��_W��`��\!�( E�0K�d_ �`;.�]�HP"�� T0 k� >3� 3UHC"!U2d   ��    � ��A^�K@��_W��`��\!�( E�0K�h` �`;.�]�HP"�� T0 k� >3�3UHC"!U2d   ��    � ��A^�K@��_W��`��\!�( E�/K�h` �`;�]�HP"�� T0 k� >2�2UHC"!U2d   ��    � ��A^�K@��_W��`��\!�( E�/K�h` �`;�]�HP"�� T0 k� �1�1UHC"!U2d   ��    � ��A^�K@��_W��`��\!�( E� /K�l` �`;�]�HQ"�� T0 k� �0�0UHC"!U2d   ��    � ��A^�K@��_W��`��\|( E��.K�l` �`;�]�HQ3� T0 k� �/�/UHC"!U2d   ��    � ��A^�K@��_W��`��\|( E��.K�l` �`;�]�HQ3� T0 k� �/�/UHC"!U2d   ��    � ��A^�K@��_W��`��\|( E��.K�l` �`;�]�HQ3� T0 k� �.�.UHC"!U2d   ��    � ��A^�L@��_W��`��\|( E��.K�pa �`;�]�HQ3� T0 k� �-�-UHC"!U2d   ��    � ��A^�L@��_W��`��\|( E��.K�pa �`;�]�HR3� T0 k� �,�,UHC"!U2d   ��    � ��A^�L@��_W��`��\|( E��-K�pa�`;�]�HR3� T0 k� �+�+UHC"!U2d   ��    � ��A^�L@��_W��`��\|( E��-K�pa�`:�]�LR3� T0 k� �+�+UHC"!U2d   ��    � ��A^�L@��_W��`��\|( L^�-K�pa�`:�]�LR3� T0 k� � *�*UHC"!U2d   ��    � ��A^�L@��_W��`��\|( L^�-K�pa�\:�]�LR3� T0 k� ��)� )UHC"!U2d   ��    � ��A^�L@��_W��`��\|( L^�-K�pb�\:�]�LS3� T0 k� ��(� (UHC"!U2d   ��    � ��A^�L@��_W��`��\|( L^�-K�pb�\:�]�LS3� T0 k� ��'��'UHC"!U2d   ��    � ��A^�L@��_W��`��\|( L^�-K�pb�\:�]�LS3� T0 k� -�'��'UHC"!U2d   ��    � ��A^�L@��_W��`��\|( L^�-K�pb�\:�]�LS3� T0 k� -�&��&UHC"!U2d   ��    � ��A^�L@��_W��`��\|( L^�,K�pb�\:^�]�LS3� T0 k� -�%��%UHC"!U2d   ��    � ��A^�L@��_W��`��\|( L^�,K�tb�\:^�]�LT3� T0 k� -�$��$UHC"!U2d   ��    � ��A^�L@��_W��`��\|( L^�,K�tb�\:^�]�PT3� T0 k� -�#��#UHC"!U2d   ��    � ��A^�L@��_W��`��\|( L^�,K�tb�\:^�]�PT3� T0 k� ��#��#UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�,K�tc�\:^�]�PT3� T0 k� ��"��"UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�,K�tc�\:��]�PT3� T0 k� ��!��!UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�,K�tc�\:��]�PT3� T0 k� �� �� UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�,K�tc�\:��]�PU3� T0 k� ����UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�+K�xc�\:��]�PU3� T0 k� ����UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�+K�xc�\:��]�PU3� T0 k� ����UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�+K�xc�\:��]�PU3� T0 k� -���UHC"!U2d  
 ��    � ��A^�M@��_W��`��\|( Ln�+K�xc�\:��]�PU3� T0 k� -���UHC"!U2d  
 ��    � ��A^�M@��_W��`��\|( Ln�+K�xd�\:��]�PU3� T0 k� -���UHC"!U2d  	 ��    � ��A^�M@��_W��`��\|( Ln�+K�xd�\:��]�TV3� T0 k� -���UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�+K�xd�\:��]�TV3� T0 k� -���UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�+K�xd�\:��]�TV3� T0 k� ����UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�+K�xd�\:��]�TV3� T0 k� ����UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�*K�xd�\:��]�TV3� T0 k� ����UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�*K�xd�\:��]�TV3� T0 k� ����UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�*K�xd�\:��]�TV3� T0 k� ����UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�*K�xd�\:��]�TV3� T0 k� ����UHC"!U2d   ��    � ��A^�M@��_W��`��\|( Ln�*K�xe�\:��]�TW3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Ln�*K�xe�\:��]�TW3� T0 k� -���UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Ln�*K�xe�\:��]�TW3� T0 k� -���UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Ln�*K�xe�\:��]�TW3� T0 k� -���UHC"!U2d    ��    � ��A^�N@��_W��`��\|( Ln�*K�xe�\:��]�TW3� T0 k� -���UHC"!U2d    ,�    � ��A^�N@��_W��`��\|( Ln�*K�xe�\:��]�XW3� T0 k� -���UHC"!U2d    ��    � ��A^�N@��_W��`��\|( Ln�*K�|e�\:��]�XW3� T0 k� ����UHC"!U2d    ��    � ��A^�N@��_W��`��\|( Ln�)K�|e�X:��]�XW3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Ln�)K�|e�X:��]�XW3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Ln�)K�|e�X:��]�XW3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Ln|)K�|f�X:��]�XW3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Ln|)K�|f�X:��]�XW3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Ln|)K�|f�X:��]�XW3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Lnx)B�|f�X:��]�XW3� T0 k� -�
��
UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Lnx)B�|f�X:��]�XW3� T0 k� -�	��	UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Lnt)B�|f�X:��]�XW3� T0 k� -���UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Lnt)B�|f�X:��]�XW3� T0 k� -���UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Lnp)B�|f�X:��]�XX3� T0 k� -���UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Lnp)B�|f�X:��]�\X3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Lnl)B�|f�X:��]�\X3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Lnl)B�|f�X:��]�\X3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Lnh(@n|f�X:��]�\X3� T0 k� ����UHC"!U2d   ��    � ��A^�N@��_W��`��\|( Lnh(@n|f�X:��]�\X3� T0 k� ����UHC"!U2d   ��    � ��A^�O@��_W��`��\|( Lnh(@n|f�X:��]�\X3� T0 k� ����UHC"!U2d   ��    � ��A^�O@��_W��`��\|( L^d(@n|f�X:��]�\X3� T0 k� ����UHC"!U2d   ��    � ��A^�O@��_W��`��\|( L^d(@n|f�X:��]�\X3� T0 k� -� �� UHC"!U2d   ��    � ��A^�O@��_W��`��\|( L^`(@n|f�X:��]�\X3� T0 k� -� �� UHC"!U2d   ��    � ��A^�O@��_W��`��\|( L^`(@n|f�X:��]�\X3� T0 k� -�����UHC"!U2d   ��    � ��A^�O@��_W��`��\|( L^`(@n|f�X:��]�\X3� T0 k� -�����UHC"!U2d   ��    � ��A^�O@��_W��`��\|( L^\(@�|f�X:��]�\X3� T0 k� -�����UHC"!U2d   ��    � ��A^�O@��_W��`��\|( D�\(@�|f�X:��]�\X3� T0 k� ������UHC"!U2d   ��    � ��A^�O@��_W��`��\|( D�\(@�|f�X:��]�\X3� T0 k� �����UHC"!U2d   ��    � ��A^�O@��_W��`��\|( D�X(@�|f �X:��]�\X3� T0 k� �����UHC"!U2d   ��    � ��A^�O@��_W��`��\|( D�X(@�|f �X:��]�\X3� T0 k� �{���UHC"!U2d   ��    � ��A^�O@��_W��`��\|( D�X)@�|f �X:��]�\X3� T0 k� �{���UHC"!U2d   ��    � ��A^�O@��_W��`��\|( D�T)@�|f �X:��]�\X3� T0 k� �w��{�UHC"!U2d   ��    � ��A^�O@��_W��`��\|( D�T)@�|f �X:��]�\X3� T0 k� �w��{�UHC"!U2d    ��    � ��A^�O@��_W��`��\|( D�T)@�|f �X:��]�\X3� T0 k� -s��w�UHC"!U2d    ��    � ��A^�O@��_W��`��\|( D�P*@�|f �X:��]�\X3� T0 k� -s��w�UHC"!U2d    ��    � ��A^�O@��_W��`��\|( D�P*@�|f �X:��]�\X3� T0 k� -o��s�UHC"!U2d    .�    � ��A^�O@��_W��`��\|( D�P*@�|f �X:��]�\X3� T0 k� -k��o�UHC"!U2d    ��    � ��A^�O@��_W��`��\|( D�L*A|f �X:��]�\X3� T0 k� -k��o�UHC"!U2d    ��    � ��A^�O@��_W��`��\|( D�L*A|f �X;��]�\X3� T0 k� �g��k�UHC"!U2d    ��    � ��A^�O@��_W��`��\|( D�L+A|f �X;��]�\X3� T0 k� �g��k�UHC"!U2d    ��    � ��A^�O@��_W��`��\|( D�H+A|f �X;��]�\X3� T0 k� �c��g�UHC"!U2d    ��    � ��A^�O@��_W��`��\|( D�H+A|f �X;��]�\W3� T0 k� �c��g�UHC"!U2d    ��    � ��                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��#8 ]�2�2� h �� Jڧ          ����     J���0    ���              ��          �     ���   	@	
          ����           ����m    �������m                   
     ��         �      ���   8�          ��/�           ��[    ��/���[                      	   �         @     ���   (
	          �          ��.      ���.                        ��$          ��     ���   H$
          \�P     	   .����     \�P����           
            �$          �     ���   H
!
           ��  ��     B�
h�      ���
h�                            ���5              C  ���      0             >g� � �
	   V����     >I���s(    ��         # R Z��         � �    ��`   8
           i�� � �
	   j��Zq     i{���O�    7 �            :	 Z��         $��    ��`   0
%            L��  � �	   ~���-     L������    �            B Z��         P�  	  ��h   0
           ]"�  � �
   ���U�     ]"���U�                      P	 Z��         	 p�    ��`   8          X�  * *	      ���ǻ     X���[}      8             $  Z��         
  ���     ��@   P
	
            ��
	      � �4�       �4�                          	  �p����             C  ��@    P                   ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��j'  ��        ��*'    ����*��    �b�C "               x                j  �   �   �                         ��    ��        ��+      ��  �+           "                                                 �                         �����������
���������� ����*�+ 
         	       
   J   ��� ��D       � @r@ �� `r� �D s� �d s� V� s� �� n� � �m@ �  n@ V� s� G$ k� H� s� �� s� � s� >  s@ � r� �  r�  s  �d u� � �r@ �  s@ 
� V� 
�� V� 
�\ W  
�\ W� 
� W� 
�\ W� �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� � }`���� � 
�| V  
� V� 
�� V� 
�\ W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������� �� Y  ������  
�fD
��L���"����D" � j  "  B   J jF�"    "�j * , ����
��"     �j @�    �
� �  �  
�  ;��  ��     ���  �   ��    ��     ���       L��  ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  ��      �� �T ���        � �  ���        �        ��        �        ��        � 	  G�    E���� u        ��                         T�) , ��� ��                                     �                ����              E�� ���%��   ����                8 Geoff Sanderson     0:01                                                                        7  6     �f � �e � � �c�K � c�C � c�C �kV2 � k^2 � k_B � 	k`B � 
ka7 � kb< �kj] � kre � ksU �ktU � kv] � kw` �c~? �c�G � c�@ �c�? �c�J �c�A �c�L � c�T � c�E � c�= �J�< � J�< �C � � C � � C � � !C" � �"J� � �#"� � � $"� � �%"� � �&*� � �'"�6 � ("�H �)�6 � 
�E � 
�E � 
�3 � 
�4 � 
�1 � 
�1X  "H �P 1"O �X  "H � �3!� x8 4"I �H 5"P �P 6"O �X  "H �X  "H �X  "H �X :"G �X  "K �8 <"D �P ="C �X >"G �X  "K �                                                                                                                                                                                                                         �� P @       �     @ 
        :     Y P E g  ���� \               	�������������������������������������� ���������	�
��������                                                                                          ��    �^~�
� ��������������������������������������������������������   �4, F  H � X� r� ��@(	��@9��@�	 A�g�������&�                                                                                                                                                                                                                                                                                                 @�����                                                                                                                                                                                                                                           
 ! &    	��  H�J      ��  	                           �������������������������������������������������������                                                                                                                                    �        9              �    �9    H        
 	  
	 
 	 	 ������������������������������������������� �� ������� ������� ���������������� �� ��� �������� ��� �������� �������������������� ���������� �������������������������������� � ����� ��� ��� ��������������� ������ ���� ���� ������                          O    .     �  D�J    	  �                             ������������������������������������������������������                                                                          	                                                      
      �      �      �        n        n  �         	  
 	 
 	 	 ������������ �� ��� ��������������� ���������������������� �������������������� �����������  � ������� ������� ������������������������������ ������������������ ������ ����������� �������������������������������� ����������������� �������      	  	   ~       	                                                                                                                                                                                                                                                                                                     �             


            �   }�         ��������������������  N�������������  V����������������  }���������  Rt  N�����������������������������                                                                 R�               ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" = E 8                	                 � xݟ� �\                                                                                                                                                                                                                                                                                     �1n  	nY                      k            e                                                                                                                                                                                                                                                                                                                                                                                                                                   2 �  2�  J�   d  <�  F_e�  �������8�X��8����B��������̞�����������b7          .  ��  � x          	�   & AG� �  q   
           �f�                                                                                                                                                                                                                                                                                                                                      C B   �         "             !��                                                                                                                                                                                                                            Y   �� �� Ѱ��      �� Z      ������������������������������������������� �� ������� ������� ���������������� �� ��� �������� ��� �������� �������������������� ���������� �������������������������������� � ����� ��� ��� ��������������� ������ ���� ���� ������������������ �� ��� ��������������� ���������������������� �������������������� �����������  � ������� ������� ������������������������������ ������������������ ������ ����������� �������������������������������� ����������������� �������   �� �     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    4      F   #  ��                       I     �  �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$    `d  �@���6 ��  �@���6 �$ ^$ �r@  �@  �r@   1 
�T ��   1 
   ���   ���� ��   ���� �$ ^$   �   �           r  ��     H � ��� �� � ��� �$ c �  ��c  �      �  ��    �����������J g���  �     f ^�         �� 4              ��#��������J���J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �   3       �  �3 3�=������<��̼��� �3 33==ƙ�<ə�ƙ�3ƙ��ƙ���i� 3= ��3=�l�ә��<��l<��l<��l<���<    �   3=  �30 ��� ���=��������                        +   3     0  �<  3� 3� =� =� 0� 0������������������3�33033�0�3�0��;f��;��̽�������3��3��<���<�f���̳=�=�������3303<�<00�<30�3����������������=��=��3�3�=�3�0  �=  �3  �3� ��0 ̳0 �0 �0  0� =� =� 3�  3�  �<  0  33�0�3�0�3�0�3303�303�303�303303��<���0<��0<033<033003300330033030�30�<00�<0330333033303330333033�0��<���0�03303303=03=03��0 ̳0 ��0 �3� �3� �=  0  3�     �                           <�03=��3=�� 3��  �=  �        033003300330�330��303= ��33    330333033303330333<��333ݰ    0=�0<3���;�3 �=  3�             �                           wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "! ""! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "! ""! " "" """ "!   " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                        "! ""! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                              "  .���"    �     �                                                                                                                                                                                     �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   �   ��  � � ��      �    �   �   �"  ""  !� �� ��  �               �   ������  ��                      �   �                      �������  ���    ��   �   ��� ������ �   �      �       �                        �   ��  ���  � �    �                                                                                                                                       	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                        �          �   � � �  ��� ��  �                       �   �                      �������  ���    �       �  �  �  �                   �     �                                                                                                                                                                                   �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �   �   "   "   "  !�    ��                              �                        ���� ��� ����                � ��                    ���� �                                                                                                                                                                                        �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                ��� ���� ��  ���� �                                                                                                                                                                                                                �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                          �  �  �  �� ݚ� }�Ȫ��˙������˼� ��  ��  ��  ��  ��  I� H� �E X�T X�S T�D �[ ˻  ˸  ��  
� �,"��"" "  �" �  ""� �� ˻ �˻ ��ݪ��کɨ��ˀ�̽ ��� ��  ̽  ̻  ̻  ˉ  ��  �D  DC  C3  #;  ;�� �� ��  �� "�  "  �"/ / ����� ��  �      �   �          �  �  "     "  "  "   "�  �  �   �   
                            �          �   �          �                    ��  ���� ��    �����                         �     �                                       �   ���                            �   �                                                                                                  "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��                       "  "  "                                                                                                                                                                               � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �                         ���                                                                                                                                                                                                                 " �"  �      �    "" ""  "!� !������������ ����  ��  "  ""  "!  "���                     
         �  � "��""- �"- "   � "� ""� ""$ "$  C  3  �  �  �   �   +w{� �װ vw� �w� ��� ɪ������˹��̻����̰݊� �ɨ �˅@̻�@�D�@4U�@4U� 4U� 4U� 3UXP�EX��U����  ��                    �  ��� ݼ� �    �    �   �                     �  �  �   �   �   �                   �   �               �  ��� ݼ� w{� �װ vw�                    �   ���                            �   �                                                                                                                         
   �   �  ��  �� ������-�� "��  �  
�  �C 
UU US �UD TE0 �� 
�� ʐ �  ̻  "�  "   " �� ����   �  �˰ ̻� �ݰ �w� ��� ����������˹�̹���ڙ��ٻ��ݰ̻� ˘  ��  3D  TD� 340 340 3D0 30 
��  ��  "/  "/  �� ���� �    ��                  "      �           �  �   �   ��  �             ��  ��  �                            �   �    �   �       �   �   �                .                         � ��                  �  �˰ ��� �wp ���                                                                                                                                                                        �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��                  �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqf � �e � � �c�K � c�C � c�C �kV2 � k^2 � k_B � 	k`B � 
ka7 � kb< �kj] � kre � ksU �ktU � kv] � kw` �c~? �c�G � c�@ �c�? �c�J �c�A �c�L � c�T � c�E � c�= �J�< � J�< �C � � C � � C � � !C" � �"J� � �#"� � � $"� � �%"� � �&*� � �'"�6 � ("�H �)�6 � 
�E � 
�E � 
�3 � 
�4 � 
�1 � 
�1X  "H �P 1"O �X  "H � �3!� x8 4"I �H 5"P �P 6"O �X  "H �X  "H �X  "H �X :"G �X  "K �8 <"D �P ="C �X >"G �X  "K �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.����������������������������������������� ��=�K�X�X�_��B�G�Q�K� � � � � � � � � � �2�0�.�����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������2�0�.� ��"�������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������/�.�7� �� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 