GST@�                                                            \     �                                               �   �                        ���2���� 
 ʱ������ĸ����������        i      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    "�j��,  " ��
  Y                                                                               ����������������������������������       ��    =b 0Qb 4 114  4c  c  c        	 
      	   
       ��G �� � ( �(                 Enn )1         88�����������������������������������������������������������������������������������������������������������������������������oo    og     +      '            ��                     	  7  V  	                  �            :8 �����������������������������������������������������������������������������                                ��  �       *�   @  #   �   �                                                                                '      E)n1n  �    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    I��XnϿD��7n�FHT|0 ���A_|bA* ��_8<3��T0 k� �W��[�%�0d  U8D"!8 ��?    � <��I��Xn��D��8n�FLU|0 ���A_xbA* ��_8<3��T0 k� NS��W�%�0d  U8D"!8 ��?    � <��I��Xn��D��9n�E�TW|0 ���A_tbA* ��_8<3��T0 k� NO��S�%�0d  U8D"!8 ��?    � <��L�Xn��D��:n�E�XX|0 ���A_pbA* ��_4<3��T0 k� NK��O�%�0d  U8D"!8 ��?    � <��L�Xn��D��<n�E�\Y|0 ���A_lbA* ��_4<3��T0 k� NC��G�%�0d  U8D"!7 ��?    � <��L�Xn��D��=n�E�`[|0 ���A_lbA* ��_0<3��T0 k� N?��C�%�0d  U8D"!7 ��?    � <��L�Xn��F�?n�D�h\|0 ���A_hbA+ ��_0<3��T0 k� �;��?�%�0d  U8D"!7 ��?   � <��L�X~��F�@n�Dl]|0 ���A_dbA+ ��_0<3��T0 k� �7��;�%�0d  U8D"!7 ��?    � <��L�X~��F�An�Dp^|0 ���A_`bA + ��_,<3��T0 k� �/��3�%�0d  U8D"!6 ��?    � <��L�X~��F�Cn�Cx`|0 ���A_\bA�+ ��_,<3��T0 k� �+��/�%�0d  U8D"!6 ��?    � <��L�X~��F�En�Cx`|0 ���A_\bA�+ ��_,<3��T0 k� �'��+�%�0d  U8D"!5 ��?    � <��L�X~��F�Fn�C|a|0 ���A_XbA�+ ��_(<3��T0 k� .��#�%�0d  U8D"!5 ��?    � <��L�X~��F�Hn�C�c|0 ���A_TbA�+ ��_(<3��T0 k� .���%�0d  U8D"!5 ��?    � <��L.�X~��F�In�B�d|0 ���A_PbA�+ ��_(<3��T0 k� .���%�0d  U8D"!4 ��?    � <��L.�W~��E��Kn�B��f|0 ���A_LbA�+ ��_$<3��T0 k� .���%�0d  U8D"!4 ��?    � <��L.�W~��E��Mn�B��g|0 ���A_LbA�+ ��_$=3��T0 k� .���%�0d  U8D"!3 ��?    � <��L.�W~��E��Nn�B��i|0 ���A_HbA�+ ��_$=3��T0 k� ����%�0d  U8D"!3 ��?    � <��L.�W~��E��Pn�A��j|0 ���A_DbA�+ ��_$=3��T0 k� ����%�0d  U8D"!2 ��?    � <��L.�VN��E��Rn�A��k|0 ���A_DbA�+ ��_ =3��T0 k� �����%�0d  U8D"!1 ��?    � <��L.�VN��E��Sn�A��l|0 ���A_@bA�+ ��_ =3��T0 k� ������%�0d  U8D"!1 ��?   � <��L.�VN�E��Un�A��m|0 ���A_<bA�+ ��_ =3��T0 k� ������%�0d  U8D"!0 ��?    � <��L.�VN{�E��Vn�@��n|0 ���A_<bA�+ ��_=3��T0 k� =�����%�0d  U8D"!/ ��?    � <��L.�VN{�E��Xn�@��o|0 ���A_8bA�+ ��_=3��T0 k� =�����%�0d  U8D"!/ ��?    � <��L.�UNw�E��Zn�@��p|0 ���A_4bA�+ ��_=3��T0 k� =�����%�0d  U8D"!. ��?    � <��L.�UNs�B��[n�@��q|0 ���A_4bA�+ ��_=3��T0 k� =�����%�0d  U8D"!- ��?    � <��L.�UNo�B��]n�@~�r|0 ���A_0bA�+ ��_=3��T0 k� =�����%�0d  U8D"!, ��?    � <��L.�UNo�B��^n�?~�s|0 ���A_,bA�+ ��_=3��T0 k� ������%�0d  U8D"!, ��?    � <��L.�UNk�B��`n�?~�s|0 ���A_,bA�+ ��_=3��T0 k� ������%�0d  U8D"!+ ��?    � <��L.�TNg�B��bn�?~�t|0 ���A_(bA�+ ��_=3��T0 k� ������%�0d  U8D"!* ��?    � <��L.�TNc�E��c^�?~�t|0 ���A_(bA�+ ��_=3��T0 k� ������%�0d  U8D"!) ��?    � <��L.�T^c�E��e^�?~�u|0 ���A_$bA�+ ��_=3��T0 k� ����ÿ%�0d  U8D"!( ��?    � <��L.�T^_�E��f^�>~�u|0 ���A_$bA�+ ��_=3��T0 k� -�����%�0d  U8D"!' ��?    � <��L.�T^[�E��h^�>~�v|0 ���A_ bA�+ ��_=3��T0 k� -�����%�0d  U8D"!& ��?    � <��L.�T^W�E��j^�>~�v|0 ���A_bA�+ ��_=3��T0 k� -�����%�0d  U8D"!% ��?    � <��L.�S^TL��k^�>~�v|0 ���A_bA�+ ��_=3��T0 k� -�����%�0d  U8D"!$ ��?    � <��L.�S^PL��m��>n�v|0 ���A_bA�+ ��_=3��T0 k� -�����%�0d  U8D"!# ��?    � <��L.�S^LL��n��>n�v|0 ���A_bA�+ ��_=3��T0 k� ������%�0d  U8D"!" ��?    � <��L.�S^LL��p��=n�v|0 ���A_bA�+ ��_=3��T0 k� ������%�0d  U8D"!! ��?    � <��L.�S^H
L��q��=n�w|0 ���A_bA�+ ��_=3��T0 k� ������%�0d  U8D"!  ��?    � <��L.�S^HL��s��=n�w|0 ���A_bA�+ ��_=3��T0 k� ������%�0d  U8D"! ��?    � <��L.�R>DL��u��=n�v|0 ���A_bA�+ ��_<3��T0 k� ������%�0d  U8D"! ��?    � <��L.�R>@L��v��=n�v|0 ���A_bA�+ ��_<3��T0 k� M�����%�0d  U8D"! ��?    � <��L.�R>@L��x��=n�v|0 ���A_bA�+ ��_<3��T0 k� M�����%�0d  U8D"! ��?    � <��L.�R><L��y��=n�v|0 ���A_bA�+ ��_<3��T0 k� M����%�0d  U8D"! ��?    � <��L.�R><L� {��<>�v|0 ���A_bA�+ ��_<3��T0 k� Mw��{�%�0d  U8D"! ��?   � <��L.�R>8L� |��<>�v|0 ���A_bA�+ ��_<3��T0 k� Ms��w�%�0d  U8D"! ��?    � <��L.�R>4L�~��<>�v|0 ���A_bA�+ ��_<3��T0 k� �o��s�%�0d  U8D"! ��?    � <��L.�Q>4L���<>�u|0 ���A_bA�+ ��_<3��T0 k� �k��o�%�0d  U8D"! ��?    � <��L.�Q>0L����<>�u|0 ���A_ bA�+ ��_<3��T0 k� �c��g�%�0d  U8D"! ��?   � <��L.�Q>0 L����<>�u|0 ���A_ bA�+ ��_<3��T0 k� �_��c�%�0d  U8D"! ��?    � <��L.�Q.,"L����<? t|0 ���A^�bA�+ ��_<3��T0 k� �[��_�%�0d  U8D"! ��?    � <��L.�Q.,%L����<? t|0 ���A^�bA�+ ��_<3��T0 k� -W��[�%�0d  U8D"! ��?    � <��L.�Q.,'L���;? t|0 ���A^�bA�, ��_<3��T0 k� -O��S�%�0d  U8D"! ��?    � <��L.�Q.()L���;? s|0 ���A^�bA�, ��_<3��T0 k� -K��O�%�0d  U8D"! ��?    � <��L�Q.(+L���;?s|0 ���A^�bA�, ��_<3��T0 k� -G��K�%�0d  U8D"!
 ��?    � <��L�P�$-L�~��;?s|0 ���A^�bA�, ��_<3��T0 k� -?��C�%�0d  U8D"! ��?    � <��L�P�$/L� ~��;?r|0 ���A^�bA�, ��_<3��T0 k� �;��?�%�0d  U8D"! ��?    � <��L�P�$1L�$~��;?r|0 ���A^�bA�, ��_<3��T0 k� �7��;�%�0d  U8D"! ��?    � <��L�P� 2L�$}��;?r|0 ���A^�bA�, ��_<3��T0 k� �3��7�%�0d  U8D"! ��?    � <��L�P� 4L�(}^�;?q|0 ���A^�bA�, ��_<3��T0 k� �+��/�%�0d  U8D"! ��?    � <��L�P� 6E�,|^�;?q|0 ���A^�bA�, ��_<3��T0 k� �'��+�%�0d  U8D"!  ��?    � <��L�P�8E�0|^�:?q|0 ���A^�bA�, ��_<3��T0 k� =#��'�%�0d  U8D"!  ,�?    � <��L�P�:E�0|^�:?q|0 ���A^�bA�, ��_<3��T0 k� =��#�%�0d  U8D"!  ��?    � <��L�P�<E�4{^�:?q|0 ���A^�bA�, ��_<3��T0 k� =���%�0d  U8D"! ��?    � <��L�P�=E�8{^�:Oq|0 ���A^�bA�, ��_<3��T0 k� =���%�0d  U8D"! ��?    � <��L�P�?E�<z^�:Oq|0 ���A^�bA�, ��_<3��T0 k� =���%�0d  U8D"! ��?    � <��L�P�AE�@z^�:Op|0 ���A^�bA�, ��_<3��T0 k� ����%�0d  U8D"! ��?    � <��L�P�BE�Dy^�:Op|0 ���A^�bA�, ��_<3��T0 k� ����%�0d  U8D"! ��?    � <��L�P�DE�Hy^�:Op|0 ���A^�bA�, ��_<3��T0 k� �����%�0d  U8D"! ��?    � <��L�P�EE�Px^�:Op|0 ���A^�bA�, ��_<3��T0 k� ������%�0d  U8D"! ��?    � <��L�P�GE�Tx^�:Oo|0 ���A^�bA�, ��_<3��T0 k� �����%�0d  U8D"! ��?    � <��L�P�IE�Xw^�:Oo|0 ���A^�bA�, ��_<3��T0 k� ,���%�0d  U8D"! ��?    � <��L�P�JE�\v^�9Oo|0 ���A^�bA�, ��_<3��T0 k� ,���%�0d  U8D"! ��?    � <��L�P�LE�`un�9Oo|0 ���A^�bA�, ��_<3��T0 k� ,���%�0d  U8D"! ��?   � <��L�P�ME�hun�9On|0 ���A^�bA�, ��_<3��T0 k� ,߁��%�0d  U8D"! ��?    � <��L�P�OE�ltn�9On|0 ���A^�bA�, ��_<3��T0 k� ,ۀ�߀%�0d  U8D"!	 ��?    � <��L�P�PE�psn�9On|0 ���A^�bA�, ��_<3��T0 k� ����%�0d  U8D"!	 ��?    � <��L�P�QE�xrn�9On|0 ���A^�bA�, ��_<3��T0 k� ��}��}%�0d  U8D"!
 *�?    � <��L.�P�SE�|qn�9On|0 ���A^�bA�, ��_<3��T0 k� ��~��~%�0d  U8D"!
 ��?    � <��L.�P�TE��pn�9Om|0 ���A^�bA�, ��_<3��T0 k� ��~��~%�0d  U8D"!	 ��?    � <��L.�P�UE��on�9Om|0 ���A^�bA�, ��_<3��T0 k� ��~��~%�0d  U8D"!	 ��?    � <��L.�P�WE��nn�9Om|0 ���A^�bA�, ��_<3��T0 k� ܿ��%�0d  U8D"!	 ��?    � <��L.�P�XE��mn�9Om|0 ���A^�bA�, ��_<3��T0 k� ܷ��%�0d  U8D"! ��?    � <��L.�P�YE��kn�9Om|0 ���A^�bA�, ��_<3��T0 k� ܳ��%�0d  U8D"! ��?    � <��L.�P�[E��jn�8Ol|0 ���A^�bA�, ��_<3��T0 k� ܯ����%�0d  U8D"! ��?    � <��L.�P�\E��jn�8Ol|0 ���A^�bA�, ��_<3��T0 k� ܫ����%�0d  U8D"! ��?    � <��L.�P�]E��jn�8Ol|0 ���A^�aA�, ��_<"���T0 k� ������%�0d  U8D"! ��?    � <��L.�P� ^E��in�8Ol|0 ���A^�aA�, ��_<"���T0 k� ������%�0d  U8D"! ��?    � <��L.�P� `E��hn�8Ol|0 ���A^�`A�, ��_<"���T0 k� ������%�0d  U8D"! ��?    � <��L.�P� bEΠgn�8Ok|0 ���A^�`A�, ��_<"���T0 k� ������%�0d  U8D"! ��?    � <��L.�P� cEΠfn�8Ok|0 ���A^�_A�, ��_<"���T0 k� ܋����%�0d  U8D"! ��?    � <��L.�P��dEΠen�8Ok|0 ���A^�_A�, ��_<"���T0 k� ܇����%�0d  U8D"! ��?    � <��L.�P��eEΤdn�8Ok|0 ���A^�_A�, ��_<"���T0 k� ܃����%�0d  U8D"! ��?    � <��L.�P��fEΤcn�8Ok|0 ���A^�^A�, ��_<"���T0 k� �����%�0d  U8D"! ��?    � <��L.�P��gEΤbn�8Oj|0 ���A^�^A�, ��_<"���T0 k� �w��{�%�0d  U8D"! ��?    � <��L.�P��hEΤbn�8Oj|0 ���A^�]A�, ��_<"���T0 k� �s��w�%�0d  U8D"! ��?   � <��L.�P��jEΤan�8Oj|0 ���A^�]A�, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��L.�P��kEΤ`n�8Oj|0 ���A^�]A�, ��_<3��T0 k� �k��o�%�0d  U8D"!  ,�?    � <��L.�P��lEΤ`n�8Oj|0 ���A^�\A�, ��_<3��T0 k� �c��g�%�0d  U8D"!  ��?    � <��L.�P��mEΤ_n�8Oj|0 ���A^�\A�, ��_<3��T0 k� �_��c�%�0d  U8D"!  ��?    � <��L.�P��nEΤ_n�7O j|0 ���A^�\A�, ��_<3��T0 k� [��_�%�0d  U8D"!  ��?    � <��L.�P��oEΤ_n�7O i|0 ���A^�\A|, ��_<3��T0 k� W��[�%�0d  U8D"! ��?    � <��L.�P��oEΤ_n�7O i|0 ���A^�[A|, ��_<3��T0 k� O��S�%�0d  U8D"! ��?    � <��L.�P��pEΤ_n�7O i|0 ���A^�[A|, ��_<3��T0 k� K��O�%�0d  U8D"! ��?    � <��L.�O��qEΤ^n�7? i|0 ���A^�[A|, ��_<3��T0 k� G��K�%�0d  U8D"! ��?    � <��L.�O��rEΤ^n�7? i!�0 ���A^�ZA|, ��_<3��T0 k� C��G�%�0d  U8D"! ��?    � <��L.�O��sEΤ^n�7? i!�0 ���A^�ZA|, ��_<3��T0 k� ?��C�%�0d  U8D"! ��?    � <��L.�O��tEΤ^n�7? i!�0 ���A^�ZA|, ��_<"s��T0 k� 7��;�%�0d  U8D"! ��?    � <��L.�O��uEΤ^n�7? h!�0 ���A_ YAx, ��_<"s��T0 k� 3��7�%�0d  U8D"! ��?    � <��L.�O��vEΤ^n�7? h!�0 ���A_ YAx, ��_<"s��T0 k� /��3�%�0d  U8D"! ��?    � <��L.�N��wA�^n�7?$h!�0 ���A_ YAx, ��_<"s��T0 k� �+��/�%�0d  U8D"! ��?    � <��L.�N��wA�^n�7?$h!�0 ���A_YAx, ��_<"s��T0 k� �#��'�%�0d  U8D"! ��?    � <��L.�N��xA�^n�7? h!�0 ���A_XAx, ��_<"s��T0 k� ���#�%�0d  U8D"! ��?    � <��L.�N��yA�^^�7? g!�0 ���A_XAx, ��_<"s��T0 k� ����%�0d  U8D"! ��?    � <��L.�N��zA�^^�7? g!�0 ���A_XAx, ��_<"s��T0 k� ����%�0d  U8D"! ��?    � <��L.�N��{A�^^�7o g!�0 ���A_XAx, ��_<"s��T0 k� ����%�0d  U8D"! ��?    � <��L.�N��{A�^^�7o g|0 ���A_WAt, ��_<"s��T0 k� ����%�0d  U8D"! ��?    � <��L.�M��zA�^^�7o g|0 ���A_WAt, ��_<"s��T0 k� ����%�0d  U8D"! ��?    � <��L�M��zA�^^�7o g|0 ���A_VAt, ��_<3��T0 k� ����%�0d  U8D"! ��?    � <��L�M��zA�^��7og|0 ���A_VAt, ��_<3��T0 k� �����%�0d  U8D"! ��?    � <��L�M��zA�^��7_g|0 ���A_VAt, ��_<3��T0 k� ������%�0d  U8D"! ��?    � <��L�M��zA�^��7_f|0 ���A_UAt, ��_<3��T0 k� �����%�0d  U8D"! ��?    � <��L�M��zA�^��7_f|0 ���A_UAt, ��_<3��T0 k� ����%�0d  U8D"!  ��?    � <��L�M��zA�^��7_f|0 ���A_UAt, ��_<3��T0 k� ����%�0d  U8D"!  ��?    � <��L�M-�zA�^��6_f|0 ���A_TAt, ��_<3��T0 k� ����%�0d  U8D"!  ��?    � <��A^�M-�zA�^��6�f|0 ���A_TAp, ��_<3��T0 k� ߎ��%�0d  U8D"!  /�?    � <��A^�L-�zA�^��6�e|0 ���A_SAp, ��_<3��T0 k� ۏ�ߏ%�0d  U8D"!  ��?    � <��A^�L-�zA�^��6�e!�0 ���A_SAp, ��_<3��T0 k� ׏�ۏ%�0d  U8D"!  ��?    � <��A^�L-�yA�^��6�e!�0 ���A_SAp, ��_<3��T0 k� ӏ�׏%�0d  U8D"!  ��?    � <��A^�L�yA�^��6�e!�0 ���A_SAp, ��_<3��T0 k� ː�ϐ%�0d  U8D"!  ��?    � <��A��L yA�^��6�e!�0 ���A_RAp, ��_<3��T0 k� ǐ�ː%�0d  U8D"!  ��?    � <��A��LyA�^��6�d!�0 ���A_RAp, ��_<3��T0 k� Ð�ǐ%�0d  U8D"!  ��?    � <��A��LxA�^��6� d!�0 ���A_RAp, ��_<3��T0 k� ���Ñ%�0d  U8D"!  ��?    � <��A��LxA�^��6��d!�0 ���A_QAp, ��_<3��T0 k� �����%�0d  U8D"!  ��?    � <��A��LxA�^��6��d!�0 ���A_QAp, ��_<3��T0 k� �����%�0d  U8D"!  ��?    � <��A��L�xA�^��6��d!�0 ���A_QAp, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��A��L�wA�^��6��d!�0 ���A_PAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��A��L�wA�^��6��c!�0 ���A_PAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��A��L�wA�^��6��c|0 ���A_PAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��A��L�vA�^��6��c|0 ���A_PAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��A��L� vA�^��6��c|0 ���A_ OAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��BN�L�$uA�^��6��c|0 ���A_ OAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��BN�L�(uA�^��6��d|0 ���A_ OAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��BN�L�,tA�^��6��d|0 ���A_ OAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��BN�L�0tA�^��6��d|0 ���A_ NAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��BN�L�4sA�^��6��d|0 ���A_$NAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��DބL�8rA�^��6��d|0 ���A_$NAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��DބL�@rA�^��6��d|0 ���A_$NAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��DބM�DqA�^��6��d|0 ���A_$MAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��DބM�HpA�^��6��c|0 ���A_$MAl, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��DވM�LoA�^��6��c|0 ���A_$MAh, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��DވM�PoA�^��6��c|0 ���A_(MAh, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��DވM�XnA�^��6��c|0 ���A_(LAh, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��DވM�\mA�^��6>�c|0 ���A_(LAh, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��D�M�`lA�^��6>�c|0 ���A_(LAh, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��D�M�dkA�^��6>�b|0 ���A_(LAh, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��D�M�ljA�^��6>�b|0 ���A_(LAh, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��D�M~ljA�^��6>�b|0 ���A_(KAh, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��D�M~pjA�^��6>�b|0 ���A_,KAh, ��_<3��T0 k� ������%�0d  U8D"!  ��?    � <��BN�M~pjA�]��6>�a|0 ���A_,KAh, ��_<3��T0 k� �����%�0d  U8D"!  ��?    � <��BN�M~tjA�]��6^�a|0 ���A_,KAh, ��_<3��T0 k� �����%�0d  U8D"!  ��?    � <��BN�M~tjA�]��6^�a|0 ���A_,KAh, ��_<3��T0 k� �{���%�0d  U8D"!  ��?    � <��BN�M^tjA�]��6^�a|0 ���A_,JAh, ��_<3��T0 k� �{���%�0d  U8D"!  ��?    � <��BN�M^tjA�]��6^�`|0 ���A_,JAh, ��_<3��T0 k� �{���%�0d  U8D"!  ��?    � <��L^�L^tjA�]��6^�`|0 ���A_,JAh, ��_<3��T0 k� �{���%�0d  U8D"!  ��?    � <��L^�L^tjA�\^�6��`|0 ���A_,JAh, ��_<3��T0 k� �w��{�%�0d  U8D"!  ��?    � <��L^�L^tjA�\^�6��`|0 ���A_0JAh, ��_<3��T0 k� �w��{�%�0d  U8D"!  ��?    � <��L^�K^tjA�\^�6��`|0 ���A_0IAh, ��_<3��T0 k� �w��{�%�0d  U8D"!  ��?    � <��L^�K^tjA�\^�6��_|0 ���A_0IAd, ��_<3��T0 k� �w��{�%�0d  U8D"!  ��?    � <��L^�K^tjA�[^�6��_|0 ���A_0IAd, ��_<3��T0 k� �s��w�%�0d  U8D"!  ��?    � <��L^�K^tjA�[^�6�_|0 ���A_0IAd, ��_<3��T0 k� �s��w�%�0d  U8D"!  ��?    � <��L^�J^tjA�[^�5�_|0 ���A_0IAd, ��_<3��T0 k� �s��w�%�0d  U8D"!  ��?    � <��L^�J^xjA�[^�5�_|0 ���A_0IAd, ��_<3��T0 k� �s��w�%�0d  U8D"!  ��?    � <��L^�JnxjA�[^�5�_|0 ���A_0HAd, ��_<3��T0 k� �s��w�%�0d  U8D"!  ��?    � <��L^�JnxjA�Z^�5�^|0 ���A_4HAd, ��_<3��T0 k� �s��w�%�0d  U8D"!  ��?    � <��L^�InxjL��Z^�5�^|0 ���A_4HAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�In|jL��Z^�5�^|0 ���A_4HAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�In|jL��Z^�5�^|0 ���A_4HAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�In|iL��Z^�5�^|0 ���A_4HAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�In|iL��Zn�5�^|0 ���A_4HAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Hn|iL��Zn�5�^|0 ���A_4GAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Hn|iL��Zn�5�^|0 ���A_4GAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Hn�iL��Zn�5�^|0 ���A_4GAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Hn�iL��Zn�5.�]|0 ���A_4GAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Gn�iL��Yn�5.�]|0 ���A_8GAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Gn�iM�Yn�5.�]|0 ���A_8GAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Gn�iM�Yn�5.�]|0 ���A_8GAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Gn�iM�Yn�5.�]|0 ���A_8GAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Gn�iM�Yn�5.�]|0 ���A_8FAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Gn�iM�Yn�5.�]|0 ���A_8FAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln�Fn�iM�Yn�5.�]|0 ���A_8FAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?   � <��Ln|Fn�iM�Yn�5.�]|0 ���A_8FAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|Fn�iM�Yn�5.�]|0 ���A_8FAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|Fn�iM�Yn�5.�\|0 ���A_8FAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|Fn�iL��Xn�5.�\|0 ���A_8FAd, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|En�iL��Xn�5.�\|0 ���A_<FA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|En�iL��Xn�5.�\|0 ���A_<FA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|En�iL��Xn�5.�\|0 ���A_<EA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|En�iL��Xn�5.�\|0 ���A_<EA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|En�iL��Xn�5.�\|0 ���A_<EA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|En�iL��Xn�5.�\|0 ���A_<EA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|Dn�iL��Xn�5.�\|0 ���A_<EA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|Dn�iL��Wn�5.�\|0 ���A_<EA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|Dn�iL��Wn�5.�\|0 ���A_<EA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|Dn�iL��Wn�5.�\|0 ���A_<EA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|Dn�iL��Wn�5.�\|0 ���A_<EA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Ln|Dn�iA�Wn�5.�[|0 ���A_<EA`, ��_<3��T0 k� �o��s�%�0d  U8D"!  ��?    � <��Hdp`��G��<I!�|0 �{�I,cE�+��Q��T0 k� �7��7%�0d  U8D"! ��*    � - �Hdp`��@���@J!�|0 �{�I$0cE�+��R��T0 k� �8��8%�0d  U8D"! ��*    � - �Hdp`��@���DK��|0 �{�I$0cE�+��S��T0 k� �9��9%�0d  U8D"! ��*    � - �Hdp`��@���HL��|0 �{�I$0cA�+��	�S��T0 k� �9��9%�0d  U8D"! ��*    � - �Hdt`��@���HM��|0 �{�I$4cA�,���T��T0 k� �:��:%�0d  U8D"! �*    � - �Hdt`��@���LO��|0B{�I$4cA�,���U��T0 k� ��;��;%�0d  U8D"! ��*    � - �Hdt`���O2��PP��|0B{�I4cA�,���V��T0 k� ��<��<%�0d  U8D"! ��*    � . �Hdt`���O2��PQ��|0B{�I4cA�-���V��T0 k� ��<��<%�0d  U8D"! ��*    � . �Hdx`���O2��TS���|0B{�I4cER -Ҽ�X��T0 k� ��>��>%�0d  U8D"! ��*    � / �Hdx`���O2��TT���|0�{�I4cER .Ҽ�X��T0 k� ��>��>%�0d  U8D"!  ��*    � 0 �Hdt_���O2��TU���|0�{�D�4dER .Ҽ�Y��T0 k� ��?��?%�0d  U8D"!  ��*    � 1 Hdt_���O2��XV���|0�{�D�4dEQ�.Ҽ�Z��T0 k� ��@��@%�0d  U8D"!  ��*    � 2 Hdt_���O2��XW���|0�{�D�4dEQ�/Ҽ�Z��T0 k� ��@��@%�0d  U8D"!  .�*    � 2 Hdt_���O2��XX���|0�{�D�4dEQ�/���[��T0 k� ��G��G%�0d  U8D"!  ��*   � 3 Hdt^���O2��XY���|0�{�D�4eEA�/����\��T0 k� ��M��M%�0d  U8D"!  ��*    � 4 A�t^���O2��XZ���|0�{�D�8eEA�0����\��T0 k� ��Q��Q%�0d  U8D"!  ��*    � 4 A�t^���O2��T\���|0�{�D�8fEA�0����^��T0 k� ��V��V%�0d  U8D"!  ��*    � 5 A�t^���O2��T\���|0�w�D�<fEA�0����^��T0 k� ��X��X%�0d  U8D"!  ��*    � 6 A�t]���O2��T]���|0�w�D�<gC��0����_��T0 k� ��Z��Z%�0d  U8D"!  ��*    � 7 A�p]���O2��P^���|0�w�D�<gC��0����_��T0 k� ��[��[%�0d  U8D"!  ��*    � 7 ATp]���O2��P_���|0�s�D�@hC��0����`��T0 k� ��]��]%�0d  U8D"!  ��*    � 8 ATp]���O2��La���|0�o�D�DiC��0����a��T0 k� �b�b%�0d  U8D"!  ��*    � 9 ATp]���O2��Lb���|0�o�D�DjC��0����b��T0 k� �f�f%�0d  U8D"!  ��*    � : ATp]��O2�Hc���|0�k�D�DjC��0����b��T0 k� �i�i%�0d  U8D"!  ��*    � : C�l]��O2�Dc���|0�k�D�DjC��0����c��T0 k� �k�k%�0d  U8D"!  ��*    � ; C�l]��O2�Dd���|0�g�D�DjC��0����d� T0 k� �m�m%�0d  U8D"!  ��*    � < C�l]��O2�<f���|0�c�D�@jC��0����d� T0 k� � p�$p%�0d  U8D"!  ��*    � < C�h]��O2�8g���|0�_�D�DkC��/����e�T0 k� � q�$q%�0d  U8D"!  ��*    � < C�h]��E� 4g��|0�[�E�DkC��/��� f�T0 k� �$r�(r%�0d  U8D"!  ��*    � < e�d\�#�E� 4h��|0�W�E�@kC��/��� f�T0 k� �$r�(r%�0d  U8D"!  ��*    � < e�d\�/�E�,j��|0�O�E�@kC��.��� g�T0 k� �v� v%�0d  U8D"!  ��*    � < �e�`\�3�E�$j��|0�K�E�DkC��-��� h�T0 k� �x�x%�0d  U8D"!  ��*   � < �e�`\�7�E�
 k��|0�G�B�DkC��-�� �h�T0 k� �z�z%�0d  U8D"!  ��*    � < �e�\\�?�E�
l��|0�C�B�DkC��-�� �i�T0 k� �{�{%�0d  U8D"!  ��*    � < �e�\[�C�E�	l��|0�?�B�DkEA�,�� �i�T0 k� � |�|%�0d  U8D"!  ��*    � < �e�\[�G�E�m�߹|0�;�B�HkEA�+�� �j�T0 k� ��}� }%�0d  U8D"!  ��*    � < �e�X[�S�E�n�ۻ|0�/�B�HkEA�*�� �l�T0 k� ��}��}%�0d  U8D"!  ��*    � < �e�X[W�E�o�׼|0�+�B�HkEA�*����l�T0 k� ��}��}%�0d  U8D"!  ��*    � < �e�XZ_�E��p�Ӽ|0�#�B�HkEA�)����m�T0 k� ��}��}%�0d  U8D"!  ��*    � < �e�TZc�E��p�Ͻ|0��B�HkEA�(����n�T0 k� ��}��}%�0d  U8D"!  ��*    � < �e�TZk�E��q�Ǿ|0��B�DkEA�(���� o�T0 k� ��}��}%�0d  U8D"!  ��*    � < �e�TZo�E��r�ÿ|0��B�DkEA|'���� p�T0 k� ��~��~%�0d  U8D"!  ��*    � < �e�PZw�E���r��|0��B�DjEAx&���� q�T0 k� ��z��z%�0d  U8D"!  ��*    � < �e�PY�E���s��|0��B�DjE1t%���� r�T0 k� ��x��x%�0d  U8D"!  ��*    � < �e�PY��E� ��t��|0���B�DjE1h$�����s�T0 k� ��w��w%�0d  U8D"!  ��*    � < �e�LY���E����u��|0���B�DjE1d#�����t�T0 k� ��v��v%�0d  U8D"!  ��*    � < �e�LY���E����u��|0��B�@jE1`"�����u�T0 k� ��v��v%�0d  U8D"!  ��*    � < �e�LY���E���v��|0�B�@iE1\!�����v�T0 k� ��v��v%�0d  U8D"!  ��*    � < �e�LX���E���v��|0�B�@iE1T ���c�w�T0 k� ��v��v%�0d  U8D"!  ��*    � < �e�HX���E���w��|0۱B�@iE1P���c�x�T0 k� �w��w%�0d  U8D"!  ��:    � < �e�HX���E���x��|0ӲB�@iE1L���c�x�T0 k� �x��x%�0d  U8D"!  ��:    � < �e�HX���E���y��|0ǳB�<iE1D���c�z�T0 k� �z��z%�0d  U8D"!  ��:    � < �e�DW���E���y{�|0��B�<iCA@���c�{�T0 k� �z��z%�0d  U8D"!  ��:    � < �e�DW���E���zw�|0��B�<iCA<���c�{�T0 k� �{��{%�0d  U8D"!  ��:    � < �e�DWs��E���zo�|0��B�<hCA8���c�|�T0 k� �|��|%�0d  U8D"!  ��:    � < �e�DWs��E���|{g�|0��B�<hCA4���c�}�T0 k� �}��}%�0d  U8D"!  ��:    � < �e�@Ws��E���t{c�|0��B�<hCA,���c�~�T0 k� �}��}%�0d  U8D"!  ��:    � < �e�@Ws�E���d|S�|0��B�<hE1$��c�~�T0 k� �}��}%�0d  U8D"!  ��:    � < �e�@Vs��D3��\}K�|0��B�8hE1 ��s�~�T0 k� �|~��~%�0d  U8D"!  ��:    � < �e�<Vs��D2���T}C�|0�B�8hE1��s�~�T0 k� �|��%�0d  U8D"!  ��:    � < �e�<Vt�D2���L~?�|0w�B�8hE1��s�~�T0 k� �x�|%�0d  U8D"!  ��:    � < �e�<Vt�D2���D~7�|0s�B�8gE1��s�~�T0 k� �p�t%�0d  U8D"!  ��:    � < �e�<Vt�D2��</�|0	�k�B�8gE1
��s�~�T0 k� �l�p%�0d  U8D"!  ��:    � < �e�<Vt�D2��4'�|0	�c�B�8gE1	��s�~�T0 k� �h�l%�0d  U8D"!  ��:    � < �e�8Ut�D2��(��|0	�W�B�8gE!��s�~�T0 k� �\�`%�0d  U8D"!  ��:    � < �A�8Ud'�D2�� ��|0	�S�@8gE!��s�~�T0 k� �X�\%�0d  U8D"!  ��:    � < �A�8Ud+�D2���|0	�K�@8gE! ��s�~�T0 k� �P�T%�0d  U8D"!  ��:    � < �A�4Ud/�D2����|0	�G�@8gE! ��s�~� T0 k� �L�P%�0d  U8D"!  ��:    � < �A�4Ud3�D2����|0	�C�@8gE ������~� T0 k� �@�D%�0d  U8D"!  ��:    � < �A�4Ud;�DB�� ��|0	�;�@8fE ������~� T0 k� �4�8%�0d  U8D"!  ��:    � < �D40VdC�DB�� �~��|0	�3�B�4fE �����t~� T0 k� �$�(%�0d  U8D"!  ��:    � < �D4,VdG�DB���~���|0	�/�B�4fE �����p~� T0 k� �� %�0d  U8D"!  ��:    � < �D4,VdK�DB���~���|0	�+�B�4fE �����h~� T0 k� ��%�0d  U8D"!  ��:    � < �D4(VdK�ER���}���|0	�'�B�4fE �����`~� T0 k� ��%�0d  U8D"!  ��:    � < �D4$VdO�ER���}��|0	�#�B�4fE �����X~� T0 k� ��%�0d  U8D"!  ��:    � < �D4$VdS�ER���}��|0	��@d4fE�����P~� T0 k� � �%�0d  U8D"!  ��:    � < �D4 VTW�ER���}��|0	��@d4fE�����L~��T0 k� ����%�0d  U8D"!  ��:    � < �DDWT[�ER���|���|0	��@d4fE�����<~"C�T0 k� ����%�0d  U8D"!  ��:    � < �DDWT[�ER���|���|0	��@d4fE�����4~"C�T0 k� ��~��~%�0d  U8D"!  ��:    � < �DDWT_�ER���|���|0	��@�4fE�����,~"C�T0 k� ��~��~%�0d  U8D"!  ��:    � < �DDW�[�C����|��|0	��@�0fE�����$~"C�T0 k� ��~��~%�0d  U8D"!  ��:    � < �DDX�W�C�����|�w�|0	��@�0fE�����~"C�T0 k� ��~��~%�0d  U8D"!  ��:    � < �DDX�S�C�����{�o�|0	��@�0eE�����~"C�T0 k� ��~��~%�0d  U8D"!  ��:    � < DDY�O�C�����{�g�|0	���@�0eE�����"C�T0 k� �~��~%�0d  U8D"!  ��:    � < }DD Y�C�C����t{�W�|0���A0eE���{���"C�T0 k� �~��~%�0d  U8D"!  ��:    � < zES�Z�?�C����l{�O�|0���A0eE���w���"C�T0 k� �~��~%�0d  U8D"!  ��:    � < wES�Z�;�C����dz�C�|0��A0eE����w����T0 k� �~��~%�0d  U8D"!  ��:    � < tES�[�7�C����\z�;�|0��A0eE����s����T0 k� ���%�0d  U8D"!  ��:    � < rES�[�/�C���Tz�3�|0��A0eE����o����T0 k� �~��~%�0d  U8D"!  ��:    � < pES�[�+�C���Lz�+�|0��C�0eE����k����T0 k� �}��}%�0d  U8D"!  ��:    � < nES�\�#�C���Dz�#�|0�߸C�0eE����g����T0 k� �}��}%�0d  U8D"!  ��:    � < lES�\��C���4y��|0�ӸC�,eE����c����T0 k� �}��}%�0d  U8D"!  ��:    � < jES�]��C���,y �|0�ϸC�,eE����_�Ҹ�T0 k� �}��}%�0d  U8D"!  ��:    � < hES�]��C���$y��|0�˸C�(eE���[�Ұ�T0 k� �}��}%�0d  U8D"!  ��:    � < eC��^��C���y��|0�øC�(eE���[�Ҩ�T0 k� �}��}%�0d  U8D"!  ��:    � < cC��^���C���y��|0�C�$eE���W�Ҡ�T0 k� �x}�|}%�0d  U8D"!  ��:    � < aC��^���C���y��|0�C�$eEq��S�Ҙ"S�T0 k� �p}�t}%�0d  U8D"!  ��:    � < _C�_��C����xo��|0�C� dEq��K�҈"S�T0 k� �`}�d}%�0d  U8D"!  ��:    � < ]C�_��C���xo��|0�C�dEq��G��"S�T0 k� �\x�`x%�0d  U8D"!  ��:    � < [C�`�ۊC���xo��|0�C�dEq��C��x"S�T0 k� �Tt�Xt%�0d  U8D"!  ��:    � < YC�`ӉD���xo��|0 ��C�dD���?��t"S�T0 k� �Pq�Tq%�0d  U8D"!  ��:    � < WC�`ωD���xo��|0 ��C�dD���;��l"S�T0 k� �Ho�Lo%�0d  U8D"!  ��:    � < UC�a��D{�o�xo��|0 ��C�dD���3��\"S�T0 k� �<l�@l%�0d  U8D"!  ��:    � < SC�a��Dw�o�xo��|0 �C�dD���/��T~"S�T0 k� �4k�8k%�0d  U8D"!  ��:   � < PC�|b��Do�o�xo��|0 w�C�dD�#�+��L~"S�T0 k� �,j�0j%�0d  U8D"!  ��:    � < NC�tb��Dk�o�x��|0 o�C� dD�#�'��D~�T0 k� �$i�(i%�0d  U8D"!  ��:    � < LC�lb��Dk�o�y��|0 g�C��dD�'�#��<~�T0 k� �k�k%�0d  U8D"!  ��:    � < JC�`c��Dc�o�y��|0 [�C��dD�+���,}�T0 k� �k�k%�0d  U8D"!  ��:    � < GC�Xc��D[��y��|0 S�D�dD�/���$}�T0 k� ��l��l%�0d  U8D"!  ��:    � < DC�Pc{�DW��z��|0K�D�dD�/��� }�T0 k� ��m��m%�0d  U8D"!  ��:    � < BC�Hds�DS��z��|0C�D�dD�3���}�T0 k� ��m��m%�0d  U8D"!  ��:    � < @C�@dk�DK��{�|0;�D�dD�3���|�T0 k� ��m��m%�0d  U8D"!  ��:    � < >C�8dc�DG��{{�|03�D�dD�7����|�T0 k� ��m��m%�0d  U8D"!  ��:    � < <C�(eO�DG��|s�|0#�D�dD�;������{�T0 k� ��l��l%�0d  U8D"!  ��:    � < :D eG�DC��}o�|0�D�dD�;������{�T0 k� ��k��k%�0d  U8D"!  ��:    � < 8De?�D?��}�k�|0�D�dD�?������z�T0 k� �k��k%�0d  U8D"!  ��:    � < 6Df7�D7��}�c�|0�D�dD�?������z�T0 k� �k��k%�0d  U8D"!  ��:    � < 4Df/�D3�?|~�_�|0��D�dD�?������y�T0 k� �j��j%�0d  U8D"!  ��:    � < 2Df'�D+�?x~�[�|0��D�dD�C������y�T0 k� �j��j%�0d  U8D"!  ��:    � < 0D�f��C�'�?t�W�|0��D�cD�C������x�T0 k� �i��i%�0d  U8D"!  ��:    � < .D�g��C��?p�S�|0��D�cD�G������x�T0 k� �i��i%�0d  U8D"!  ��:    � < ,D�g��C��?l�K�|0�߸D�cD�G������w�T0 k� �h��h%�0d  U8D"!  ��:    � < *D�g��C��?h��G�|0�׸D�cD�K������w�T0 k� �h��h%�0d  U8D"!  ��:    � < (D�g��C��?`�;�|0�ǸD�cD�K������v�T0 k� �tf�xf%�0d  U8D"!  ��:    � < &D�h��C��?\�4|0߿�DxcD�O������u�T0 k� �lf�pf%�0d  U8D"!  ��:    � < $D�h��C��?X�0|0߷�DpcD�O�q����u�T0 k� �de�he%�0d  U8D"!  ��:    � < "D�h�ہC���?T(|0߫�DhcD�S�q��ѐt�T0 k� �Xd�\d%�0d  U8D"!  ��:    � <  D�h�ρC���?P~$|0ߣ�D`cD�S�q��шs�T0 k� �Pb�Tb%�0d  U8D"!  ��:    � < D�i�ǂC���?L~|0ߛ�C�XcEqS�q��рs�T0 k� �Ha�La%�0d  U8D"!  ��:    � < D�i⿂C���?H~|0ߓ�C�LcEqW�q���xr�T0 k� �@a�Da%�0d  U8D"!  ��:    � < D�i�C���?@}
|0߃�C�<cEq[����lq�T0 k� �4_�8_%�0d  U8D"!  ��:    � < D�i�C�� ?<}
|0�{�C�4cEq[����dp�T0 k� �,_�0_%�0d  U8D"!  ��:    � < D�j�C�� ?8}
�|0�s�C�,cEq[����\o�T0 k� �$^�(^%�0d  U8D"!  ��:    � < D�j�C�� ?4}
�|0�k�C�$cEq_����To�T0 k� �]� ]%�0d  U8D"!  ��:    � < C�xj�C� ?4|
�|0�c�C�cEq_����Pn�T0 k� �\�\%�0d  U8D"!  ��:    � < C�pj�C� ?0|
�|0�_�C�cEa_�����Hm�T0 k� �\�\%�0d  U8D"!  ��:    � < C�`k�s�C�?(|
�|0	�O�C� cEac�����8l�T0 k� � Z�Z%�0d  U8D"!  ��:    � < C�Xk�k�C�?$|
�|0	�K�C��cEac�����0k�T0 k� ��Y��Y%�0d  U8D"!  ��:    � < 
C�Pk�c�C�?${ �|0	�C�C��cEac�����,j�T0 k� ��Y��Y%�0d  U8D"!  ��:    � < C�Hk[�D�? { �|0	�?�C��cEac�����$i�T0 k� ��X��X%�0d  U8D"!  ��:    � < C�@kS�D|?{ �|0	�7�C��cEac�
A���i3�T0 k� ��W��W%�0d  U8D"!  ��:    � < C�<kG�Dt?{ �|0	�3�C��cEa_�
A���h3�T0 k� ��V��V%�0d  U8D"!  ��:    � < C�4l?�Dl?{ �|0	�+�C��cEa_�
A���g3�T0 k� ��V��V%�0d  U8D"!  ��:    � <  C�$l/�DX?z �|0	�#�C�cEa[�
A��� e3�T0 k� ��T��T%�0d  U8D"!  ��:    � <��C�l'�DP?z �|0	��C�cEaW�!����e3�T0 k� ��S��S%�0d  U8D"!  ��:    � <��C�l�DH?z �|0��C�cEaW�!����d3�T0 k� �S��S%�0d  U8D"!  ��:    � <��C�l�D@?z �!�0��C�cEaS�!����c3�T0 k� �S��S%�0d  U8D"!  ��:    � <��C�m�D4�z �!�0��C�cEQO�!����b3�T0 k� �S��S%�0d  U8D"!  ��:    � <��C��m�D,� y � !�0��D�cEQO�!����a3�T0 k� �R��R%�0d  U8D"!  ��:    � <��EQ�m��D$� y �!!�0���D�cEQK�1����`3�T0 k� �Q��Q%�0d  U8D"!  ��:    � <��EQ�m�D��y �!!�0���DxcEQG�1��P�`3�T0 k� �V��V%�0d  U8D"!  ��:    � <��EQ�m�D�x �"!�0��DdcEQC�1��P�^3�T0 k� �Y��Y%�0d  U8D"!  ��:    � <��EQ�nۇD �w �#!�0��D\cEQ?�1��P�]3�T0 k� �[��[%�0d  U8D"!  ��:    � <��EQ�nӈD��w |#!�0��DTcEQ;�A��P�]3�T0 k� �]��]%�0d  U8D"!  ��:    � <��EQ�nˈE���v |$!�0�۴DLcEQ7�A��P�\3�T0 k� ��^��^%�0d  U8D"!  ��:    � <��EQ�n��E���v x$!�0�״D@cEQ3�A��`�[3�T0 k� �t]�x]%�0d  U8D"!  ��:    � <��EQ�n��E����u t$|0�ӳD8cC�/�A��`�Z3�T0 k� �d[�h[%�0d  U8D"!  ��:    � <��EQ�n��E����t t$|0�˲D0cC�+�A��`�Z3�T0 k� �XZ�\Z%�0d  U8D"!  ��:    � <��EA�n��E����t p%|0�ǲD(cC�'�Q��`�Y3�T0 k� �LY�PY%�0d  U8D"!  ��:    � <��EA�oᗉE���r l%|0���DbC� Q��P�X3�T0 k� �<X�@X%�0d  U8D"!  ��:    � <��EA�oᏉE���q l%|0���DbC�Q��P|W3�T0 k� �8W�<W%�0d  U8D"!  ��:    � <��EA�oᇉE���q h%|0���DbC�Q��PtV3�T0 k� �0W�4W%�0d  U8D"!  ��:    � <��Eрo�{�E��~�p h%|0���D�bC�Q��PlV3�T0 k� �(V�,V%�0d  U8D"!  ��:    � <��E�xo�s�D0�~�o h%|0��D�bC�Q��PhU3�T0 k� �$U�(U%�0d  U8D"!  ��:    � <��E�po�k�D0�~�n d%|0��D�bC� Q��P`U3�T0 k� �U� U%�0d  U8D"!  ��:    � <��E�ho�c�D0�~�m d%|0��D�bC��a��P\T3�T0 k� �T�T%�0d  U8D"!  ��:    � <��E�`o�[�D0x~�l d%!�0��D�bC��a��PTS3�T0 k� �T�T%�0d  U8D"!  ��:    � <��E�\o�S�D0p~�l d%!�0��D�bC��a��PPS3�T0 k� �S�S%�0d  U8D"!  ��:    � <��E�To�K�D0h~�k d%!�0��C��bC��	a��PHR3�T0 k� �R�R%�0d  U8D"!  ��:    � <��C�Lo�?�D0`	~�j d%!�0��C�bC��
a��PDR3�T0 k� � R�R%�0d  U8D"!  ��:    � <��C�Dp�7�D0T	~�i d%!�0��C�bC��Q��P<Q3�T0 k� ��Q��Q%�0d  U8D"!  ��:    � <��C�<p�/�D0L	~�i
d%!�0��C�bC��Q��P8P3�T0 k� ��Q��Q%�0d  U8D"!  ��:    � <��C�4p�'�D0D	��h
d%!�0��C�bC��Q��P4P3�T0 k� ��P��P%�0d  U8D"!  ��:    � <��C�,p��D0<
��g
`%!�0��C�bC��Q��P,O3�T0 k� ��P��P%�0d  U8D"!  ��:    � <��EA$o��D00
��f
`%!�0���C�bC��Q��P(O3�T0 k� ��O��O%�0d  U8D"!  ��:    � <��EAo��D@(
��f
`%!�0��C�bC��Q��P$N3�
T0 k� ��N��N%�0d  U8D"!  ��:    � <��EAo��D@ 
��e
\%!�0��C�|bC�A��PN3�
T0 k� ��N��N%�0d  U8D"!  ��:    � <��EAo���D@��d
\%|0�{�C�tbC�A��PM3�	T0 k� ��M��M%�0d  U8D"!  ��:    � <��EAo��D@��d
\%|0�{�C�hbD �A��PM3�	T0 k� ��M��M%�0d  U8D"!  ��:    � <��E@�o��D@��c
X%|0�w�C�`bD �A��PL3�T0 k� ��L��L%�0d  U8D"!  ��:    � <��C��o��DO���b
X%|0�w�C�XbD �A��PL3�T0 k� ��L��L%�0d  U8D"!  ��:    � <��C��n�ۋDO���b
T%|0�w�C�PbD �A��PK3�T0 k� ��K��K%�0d  U8D"!  ��:    � <��C��n ӌDO���a
P%|0�w�C�DbD �A��P K3�T0 k� /�J��J%�0d  U8D"! �:    � <��C��n ǌDO���`
.P%|0�w�C�<bEP�A����J3�T0 k� /�I��I%�0d  U8D"! ��?    � <��C��m ��DO���`
.L%|0�w�C�4bEP� �����J3�T0 k� /�G��G%�0d  U8D"! ��?    � <��C��m ��DO���_
.D%|0�w�C� bEPp �����I3�T0 k� /�E��E%�0d  U8D"! ��?    � <��C��l ��D_���^
.D%|0�w�C�bEPh �����I3�T0 k� /�C��C%�0d  U8D"!	 ��?    � <��C��l ��D_���^
.@%|0�w�C�bEP` �����H3�T0 k� ��B��B%�0d  U8D"! ��?    � <��C��l ��D_���]
.<%|0�w�C�bEPX �����H3�T0 k� ��@��@%�0d  U8D"! ��?    � <��C��k ��D_���\
.8%|0�w�C��bEPP �����G3�T0 k� ��?��?%�0d  U8D"! ��?    � <��C��k ��D_���\
.4%|0�{�D �bEPL �����G3�T0 k� ��>��>%�0d  U8D"! ��?    � <��C��j {�D_���[
.0%|0�{�D �bEPD �����G3�T0 k� ��<��<%�0d  U8D"! ��?    � <��C��js�D_���[
.,%|0�{�D �bEP< �����F3�T0 k� ?�;��;%�0d  U8D"! ��?    � <��C��ik�D_���Z
$%|0�{�D �bE@4A����F3�T0 k� ?|9��9%�0d  U8D"! ��?    � <��C��ic�D_t��Z
 %|0�{�D �bE@,A����E3�T0 k� ?x8�|8%�0d  U8D"! �?    � <��C�|h[�E�l��Y
%|0��AP�bE@$A����E3�T0 k� ?t7�x7%�0d  U8D"! �?    � <��E�thO�E�d��Y
%|0��AP�bE@A����E3�T0 k� ?p5�t5%�0d  U8D"! ��?    � <��E�lgPG�E�\��X
%|0��AP�bE@A���D3�T0 k� �h4�l4%�0d  U8D"! ��?   � <��E�dgP?�E�T��X�%|0��AP�bE@ ����D3�T0 k� �d2�h2%�0d  U8D"! ��?    � <��E�\fP7�E�H��W�%|0��AP�bE@ ����D3�T0 k� �`1�d1%�0d  U8D"! ��?    � <��E�TfP/�E�@��W�%|0 ��AP�bE@  ����C3�T0 k� �X0�\0%�0d  U8D"! ��?    � <��E�PeP'�E�8��V�%|0 ���AP�bEO�  ����C3�T0 k� �T.�X.%�0d  U8D"! ��?    � <��E�HeP�E�0��V�%|0 ���AP�bA�  ����C3�T0 k� /P-�T-%�0d  U8D"! ��?    � <��E�@e@�E�$��U�%|0 ���AP�bA�! ����B3�T0 k� /L+�P+%�0d  U8D"!  ��?    � <��E�8d@�E���U�&|0 ���AP|bA�! ����B3�T0 k� /D*�H*%�0d  U8D"!" ��?    � <��C�0d@�E���U�&|0 ���APtbA�" ����B3�T0 k� /@)�D)%�0d  U8D"!# ��?    � <��C�(cO��E���T� &|0 ���APlbA�" ����A3�T0 k� /<'�@'%�0d  U8D"!$ ��?    � <��C� cO�E���T� &|0 ���APdbA�# ����A3�T0 k� �8&�<&%�0d  U8D"!% ��?    � <��C�bO�E����S� '|0 ���AP`bA�# ����A3�T0 k� �0$�4$%�0d  U8D"!& ��?    � <��C�bO�E����S� '|0 ���APXbA�# ����@3�T0 k� �,#�0#%�0d  U8D"!' ��?    � <��C�bO׏E����S��'|0 ���APPbA�$ ����@3�T0 k� �("�,"%�0d  U8D"!( ��?    � <��C�aOϐE����R��(|0 ���APHbA�$ ����@3�T0 k� �  �$ %�0d  U8D"!) ��?    � <��C��aOǐE����R��(|0 ���APDbA�% ����?3�T0 k� O� %�0d  U8D"!* ��?    � <��C��aO��E����Q��)|0 ���AP<bA�% ����?3�T0 k� O�%�0d  U8D"!* ��?    � <��C��`?��E����Q��)|0 ���AP4bA�% ���_�?3�T0 k� O�%�0d  U8D"!+ ��?    � <��C��`?��D����Q��*|0 ���AP0bA�& ���_�?3�T0 k� O�%�0d  U8D"!, ��?    � <��C��_?��D����P��*|0 ���AP(bA�& ���_�>3�T0 k� O�%�0d  U8D"!- ��?    � <��C��_?��D����P�+|0 ���AP bA�' ���_�>3�T0 k� ��%�0d  U8D"!. ��?    � <��C��_?��D����P�+|0 ���APbA�' ���_|>3�T0 k� ��� %�0d  U8D"!. ��?    � <��C��^?��D����O�,|0 ���APbA�' ���_x>3�T0 k� ����%�0d  U8D"!/ ��?    � <��C��^?��E����O -|0 ���APbA�( ���_x=3�T0 k� ����%�0d  U8D"!0 ��?    � <��C��^?�E����O -|0 ���APbA�( ���_t=3�T0 k� ����%�0d  U8D"!1 ��?    � <��C��]?w�E����N .|0 ���APbA�( ���_t=3�T0 k� .���%�0d  U8D"!1 ��?    � <��C��]?s�E�x ��N/|0 ���A_�bA|) ���_p=3�T0 k� .���%�0d  U8D"!2 ��?    � <��C��]Ok�E�p!��N0|0 ���A_�bAx) ���_l<3�T0 k� .���%�0d  U8D"!2 ��?    � <��C��\Oc�E�h"^�M1|0 ���A_�bAt) ���_l<3�T0 k� .���%�0d  U8D"!3 ��?    � <��C��\O[�E�\"^�M1|0 ���A_�bAp* ���_h<3�T0 k� .���%�0d  U8D"!3 ��?    � <��C��\OW�E�T#^�M2|0 ���A_�bAl* ���_h<3�T0 k� ��
��
%�0d  U8D"!4 ��?    � <��D�\OO�FL$^�L3|0 ���A_�bAh* ���_d;3�T0 k� ��	��	%�0d  U8D"!4 ��?    � <��Dx[OG�FD%^�L4|0 ���A_�bAh* ���_d;3� T0 k� ����%�0d  U8D"!5 ��?    � <��Dp[OC�F<&^�L5|0 ���A_�bAd* ���_`;3� T0 k� ����%�0d  U8D"!5 ��?    � <��Dh[O;�F4'^�K6|0 ���A_�bA`* ���_\;3� T0 k� ����%�0d  U8D"!6 ��?    � <��DdZO7�F4'^�K7|0 ���A_�bAX* ���_\<3� T0 k� >���%�0d  U8D"!6 ��?    � <��D\ZO/�D�0'^�K9|0 ���A_�bAT* ���_X<3� T0 k� >���%�0d  U8D"!6 ��?    � <��DTZO'�D�((^�K:|0 ���A_�bAP* ���_X<3� T0 k� >� �� %�0d  U8D"!7 ��?    � <��DLZO#�D�$(^�J<|0 ���A_�bAL* ���_T<3� T0 k� >�����%�0d  U8D"!7 ��?    � <��DDY_�D� )^�J=|0 ���A_�bAH* ���_T<3� T0 k� >�����%�0d  U8D"!7 ��?    � <��D<Y_�D�*^�J?|0 ���A_�bAH* ���_P<3� T0 k� ������%�0d  U8D"!8 ��?    � <��D4Y_�D�*^�J @|0 ���A_�bAD* ���_P<3� T0 k� ������%�0d  U8D"!8 ��?    � <��D,Y_�D�+n�I. B|0 ���A_�bA@* ���_L<3� T0 k� ������%�0d  U8D"!8 ��?   � <��D$X_�D�,n�I.$D|0 ���A_�bA<* ���_L<3��T0 k� ������%�0d  U8D"!8 ��?    � <��DX_�D�-n�I.$E|0 ���A_�bA8* ���_L<3��T0 k� ������%�0d  U8D"!8 ��?    � <��DX^��D� -n�I.(G|0 ���A_�bA4* ���_H<3��T0 k� .�����%�0d  U8D"!8 ��?    � <��DX^��D��.n�H.,H|0 ���A_�bA0* ���_H<3��T0 k� .�����%�0d  U8D"!8 ��?    � <��I�W^�D��/n�H0J|0 ���A_�bA,* ���_D<3��T0 k� .{���%�0d  U8D"!9 ��?    � <��I� W^�D��0n�H4K|0 ���A_�bA(* ���_D<3��T0 k� .w��{�%�0d  U8D"!9 ��?    � <��I��W^�D��1n�H4M|0 ���A_�bA(* ���_@<3��T0 k� .s��w�%�0d  U8D"!9 ��?    � <��I��Wn�D��2n�G8N|0 ���A_�bA$* ���_@<3��T0 k� �o��s�%�0d  U8D"!9 ��?    � <��I��WnߺD��3n�G<P|0 ���A_�bA * ���_@<3��T0 k� �g��k�%�0d  U8D"!9 ��?    � <��I��Wn׻D��4n�G@Q|0 ���A_�bA* ��_<<3��T0 k� �c��g�%�0d  U8D"!8 ��?    � <��I��XnӽD��6n�FDS|0 ���A_�bA* ��_<<3��T0 k� �_��c�%�0d  U8D"!8 ��?    � <��                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��N� ]�'�'� H �� D9_  � �	    ���0�     D]���<i    ���R              L Z���         +@�  	  ���   0
% 	           i[g   � �	    ����2     id�����    �q�            q Z��         �P�    ���   0
 
          W�.        ���     W�.���                    p	 Z��         ��     ���  8	           5��   � �	    ���n     5������    ����   
            o  Z��          � �    ���   8          [�l   � �
	   .����     \
8���     ���i            D Z��         �@�    ���   P
	
          ��  ��	      B�2�     ���2�                             ���               �  ���    P             ���l   `       V��O�    ���q��O�     K              � 6         0     ��@   (          E
�         j����     E!�����    ��               r 6         �     ��@   8�           ,{+       ~���     ,{+����      ��           �� @         	`     ��@   	@


          ��m   U      � �$�    �� �$�     ,                    X         	 Ґ     ��@ @ H	$
          <�W    
	  ���p     <�W��p                          �         
 �     ��J   H!	         ��< ��
     � ���    ��< ���                             ���I              [  ��@      0                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         ���A  ��        ���I�    ��Q���I�    
                     x                j  �   �
   �                         ��    ��        ���      ��  ��           "                                                �                         ����������������� ��� �������    	 
            
  % 
  4� S��I       � �`� �  a� �d b  ۄ b  �� b  � b  #� `e� $d f����. ����< ����J ����X ����J ����X � 
�< V� 
�� V� 
�\ W  
�� V� 
�\ W  
�< W� 
� W� 
�\ W� �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �� �R� � }`���� � 
�| W ���� � 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������� <�� Y  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    "�j�� , " �
� �  �  
�  K    ��     �    �    5��  ��     ���       <    ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �?!!      ��CT ���        �T ���        �        ��        �        ��        �  
  ��     ���`-��        ��                         T�) ,  ���                                    �                 ����           
 K  
���%��   <����               85 Petr Klima on i     0:01                                                                        3  1      � �k~ � �k� � �J� �J� �J� � J� � �J� �B�) �	B�* �
B�" � B�1 �B�  �K �K �C � � K �C � �C � �C � � C" � �C# � �C. � C6' � C7 � C8 � C9 � C: �c� � � c�  �kj � kr � "� � � !"� � �""� � �#*� � �$"� � � %"� �&� � �'
� � � (*Kt � )*>|7  *l �+**| �,*l � -*Fd �.*2t/*:d/ 0*Gd?  *Ad?  *Bd/  *Et4*:d 5*Pt-6)�dE 7*&|U **|X **|3:)�dK ;*&|[ **|< )�d? )�d2  *Kd                                                                                                                                                                                                                         �� R @      �    @ 
        >     a P E c  ��        
           	 �������������������������������������� ���������	�
��������                                                                                          ��    �7H�� ��������������������������������������������������������   �4, :  * X� �	@��A	�����	���	                                                                                                                                                                                                                                                                                                                               �                                                                                                                                                                                                                                               ^    )    ��  D�J    	  P  	                           ������������������������������������������������������                                                                     	                                                                  �      �      �        �          �     �    	  
 	 
 	 	 � ��������������������������������� ����������� ����� ����������������� ������������ ������� � ������������������������ � ������������������������������������������������� ������������������������ �� �����  ���������������� �� ���������                          	       %  	  3    �	�  H�J      �a                             ������������������������������������������������������                                                                                                                                  
       � �     �      �        �    ��              
 	  
	 
 	 	 ������������� �� ����  ��������� �� ����������� �������� ��������������� ��� ����� ������� ��  �������������������������� ���������������������������������������������������������������������  ���������������� �������������  �� �����              �                                                                                                                                                                                                                                                                                           
                  �             


            �   }�                       O           N�                              R�              'u      ������������������������������������    ����������������    ��������  's  's����������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" A C 6               	                  � �x� �\                                                                                                                                                                                                                                                                                      E)n1n  �             W       m      m      l            a                                                                                                                                                                                                                                                                                                                                                                                                                       
 R  >�  J�  (�  (�  EZmw ����.��v���H������ �N =���������������                ���G :����        	 �   & AG� �   A                 �                                                                                                                                                                                                                                                                                                                                      p B C   =                       !��                                                                                                                                                                                                                            Y��   �� �� ��      �� B 	     � ��������������������������������� ����������� ����� ����������������� ������������ ������� � ������������������������ � ������������������������������������������������� ������������������������ �� �����  ���������������� �� ���������������������� �� ����  ��������� �� ����������� �������� ��������������� ��� ����� ������� ��  �������������������������� ���������������������������������������������������������������������  ���������������� �������������  �� �����               ���������������������������������������������������f��ff�fff�ff���������l�ff�ffffl��ff˼fllf������l��̼�ʗ���˹�ffjz�fkyl�l��fƨ�����������������������̼��̉������������������������������f���f�fff�ff�ffl�ff�flfl�l��xl�wwl���l̻�����˺��fl����l�xx��w��̻���l�f�f�ƻ�fl�����ffl�ffffffff���f���̚���ffflffflfffffffffflfffff������������������������l���l������f����������������������������l��lf��f�fff�f��l˪���ww��w�����flflffffffff�̼̙��fww��w��fx�̻�llffff�ffff���fl���f�l�l�˶����fffl��fflfll����ff��ff��lfl�lf��l���l�����������l�������l�������ʼ�j˚��̩��ʨ��ɘ���xxxȈ��ɉ�x���̇�̺������www��ww��xw���x��xk�����������wx��������������x����l�ƈ��Ƈ���w��Ɨ��̩z�̩yf̪�f�������������������������������̙i���ɖ�yɌ��ˌȉ̚ə̩���ə��Ɉ����x�̹x�̹�����������ƺ�������������������ˈ������˙������̫��̺�������˪�������������̸��̗�����̇��̇�����������������������̈���xx����x���w���ɉ��̨���k���̛̻�������������l��Ʀl�Ɗl�l���̻�lk��̺�f̩�l��f�ɫ�ˉ�lɊ�˙���ʚ���˙�˫̼���ɬ�̚��̼�����̼���̬������̼�����˻������������f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff���m�    ;      @     ��                       B     �   ���������J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �f ��        p���� ��   p���� �$     \   �4  \ >�������J J  \ \   �4  \   i  ��   �    >  H��� ��  H��� �$ ^$      H    | 
l� �� | 
l� �$ ^$ � ��� �� � ���  � � � �  �� �  �      �  ��   �������2����   g���  �     f ^�         ��  <            ��O>���2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "" "  """               "  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               ""   "! " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """               "  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        ۻ� ۽� ��� H�DH�D�DP�E X�T H�P H�@ Ȥ� ̻� ˘ �� "*� �/�""/""/���                       ��  ۼ� ݻ� w�� b}ذgvz�w������ɨ�ͨ���ڋ��٭���ۻݻ� �   �          �   �   .   ."  ""  ""  ,   �   
            "  "  ""  "�   �           �   ��  �      �                                     �  �  �  ��  �  �  �  ��  �             �   �   �             � � "            � "�",�"+� ",                       "  .���"    �     �                         � �������������  �                                �   �    ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         ۻ� ۽� ��� H�DH�D�DP�E X�T H�P H�@ Ȥ� ̻� ˘ �� "*� �/�""/""/���                       ��  ۼ� ݻ� w�� b}ذgvz�w������ɨ�ͨ���ڋ��٭���ۻݻ� �   �          �   �   .   ."  ""  ""  ,   �   
            "  "  ""  "�   �           �   ��  �      �                                     �  �  �  ��  �  �  �  ��  �             �   �   �             � � "            � "�",�"+� ",                       "  .���"    �     �                       �   ��  ���  � �    �                                                                                                                                        
� �� ���̹����̹������������̳��#3 �"T .� "U 
�U 
�U ET EC DL ��� ��  �� �� "  ""/"/�����  �           �z�����̙�����ؚ��ک��Ћ�� ˻  ��@ ��@4D����U T4UPCDEPC4U@0�D@0��� ��  ��  ""  """ "" �"������� �                         �   �   �� �� .� .� ��"       �   �                            �� ۼ�����wp���vvp�ww�             �                  �  �  �                              �  �� ��  �    � ���                                                                                                                                                                                             ۻ� ۽� ��� H�DH�D�DP�E X�T H�P H�@ Ȥ� ̻� ˘ �� "*� �/�""/""/���                       ��  ۼ� ݻ� w�� b}ذgvz�w������ɨ�ͨ���ڋ��٭���ۻݻ� �   �          �   �   .   ."  ""  ""  ,   �   
            "  "  ""  "�   �           �   ��  �      �                                     �  �  �  ��  �  �  �  ��  �             �   �   �             � � "            � "�",�"+� ",                       "  .���"    �     �                                                                                                                                                                                         �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��  ��  �   ��  �                                                                                                                                                                                                                       �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                    �  ��� ��� }�� wݪ �� 	�� �� �ͼ ��� ��� ̘� �ͻ +���"�8"8  8� �� �U��EU��3 ̻�"̰""�" ��" �"                             �   ��� �˹��˚���ڍ�̽���ͽ��ͽ���ݼ��л�� ��D �UT EUT UU0 C3  2"  ""  -�  ��  ��  �   � ��"/ �" � ���    �        �   ��  ��  ��  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��� ���� ��             �  �˰ ��� �wp ���                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  �   �   �                           �   �   �   �      �  �                         �  ���       ����������                                ��  ��  ��� �"�!/"�  �                                                                                                                                                                                                �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �        �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����            �  �  ��  �   �   �        �  �  �   �   ��  �                            �   ���                            �   �    ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                             �  ɪ� ɪ� ̚� �ȍ ͷ  "�  "� .( 3># �4�
�T��T�"�UN"�UN(�Dɜ� ʨ����, � /�������� � ��                                ��  ��  ��  g}  �א vz� gz� ̊� �ɩ 8̜ D<� T� @��  �� ɀ ��  ��  "   .          �  ��� �������  ��                           "  "  "  "                                              ��                  �                        ���� ��� ����                            �   ���       ���� �                                                                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                    ""  ."  �"    �   ��  �   �                  �  �  �  �                                       �  �   ��                     �    � �  ��                  ���                                      ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                                     �� ̻ ��˛��  �� �˚̻���ۚ����I���䘼�^���^�٘�:�^�� ^�� D�( �) �) �) ��) ˹� ț�+��,��,����  �𫝝 ��� �ɍ ��ݨ��ډ�݊�� ��D@ �D�  J�� ݩ� ��� �ۻ �ک �ڹ�ɻ��̸���������� ����������            �   ��  ��  ��  ��  ��                                          �� ��� ��� ��  �                         �   �                    �          �         �   �  �  �   �               �   �                               � ����ݼ� ����                                                                                                                                                                             �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                             DD A@A@DD@ DD                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=LL����������D����3333DDDD    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����������A������ x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx""""�������I�I������ w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww""""�������I��D���I�������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(�D�M�D���M������3333DDDD �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""�����AMAD������ M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M""""������������������ � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �k~ � �k� � �J� �J� �J� � J� � �J� �B�) �	B�* �
B�" � B�1 �B�  �K �K � K � K �C � �C � �C � � C" � �C# � �C. � C6' � C7 � C8 � C9 � C: �c� � � c�  �kj � kr � "� � � !"� � �""� � �#*� � �$"� � � %"� �&� � �'
� � � (*Kt � )*>|7  *l �+**| �,*l � -*Fd �.*2t/*:d/ 0*Gd?  *Ad?  *Bd/  *Et4*:d 5*Pt-6)�dE 7*&|U **|X **|3:)�dK ;*&|[ **|< )�d? )�d2  *Kd3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�����������������������������������������#��-�X�G�O�M��<�O�S�V�Y�U�T� � � � � � � �/�.�7����������������������������������������#� ��9�K�Z�X��5�R�O�S�G� � � � � � � � � � �/�.�7�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������/�.�7� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            