GST@�                                                            \     �                                               �   �                        ���2���
�	 ʰ������̸��h�������        i      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     "�j  " ���
��
�"    B�jl �   B ��
  C�                                                                              ����������������������������������      ��    oo= 0 go4  1  +      '      ��                 	� 7� V� 	�                 � 
         8:�����������������������������������������������������������������������������������������������������������������������������=o  0  4g  1                      �                         �  �  �  �                  ͛  	          8 �����������������������������������������������������������������������������                                ��  �       �   @  #   �   �                                                                                '    �
  	��    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E & �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    D�@�۶E�� C��m�'|(D1c��@P���`6Z3��CT0 k� ������%2't �H%1p   ��8    � #��Eq@�׷E��C��
=�&|(D1[��8P���`5Z3��BT0 k� ������%2't �H%1p   ��8    � "��EqD�ϸE��C��=�$|(D1S��0P���`4Z3��@T0 k� �����%2't �H%1p   ��8    � !��EqD�ǹEмC��=�#|(D1K��(P���`4Z3���?T0 k� �{���%2't �H%1p   ��8    �  ��EqH���EаC�l=� |(E�;��P���`2Z3���;T0 k� �s��w�%2't �H%1p   ��8    � ��EaL���EШC�d =�|(E�3��P���`1Z3���:T0 k� �o��s�%2't �H%1p   ��8    � ��EaL���EРC�_�=�|(E�'��P���`0Z3���8T0 k� �k��o�%2't �H%1p   ��8    � ��EaL���EИC�W�=�|(E���P���`/Z3���7T0 k� �g��k�%2't �H%1p   ��8    � ��EaP���C��C�O�M�|(E����P���`.Z3���5T0 k� �_��c�%2't �H%1p   ��8    � ��EaP	���C��C�G�M�|(E����P{��`-Z3���3T0 k� �[��_�%2't �H%1p   ��8    � ��D1P
���C��C�?�M�|(E�� �Pw��`,Z3���1T0 k� �W��[�%2't �H%1p   ��8    � ��D1P���C�pC�+�M�|(E��� �Po��`*Z3���.T0 k� �K��O�%2't �H%1p   ��8    � ��D1T�{�C�lC�#�M�|(E��� �@g��`)Z3���,T0 k� �G��K�%2't �H%1p   ��8    � ��D1T�s�C�d	C��M�|(E��� �@c��`(Z3���*T0 k� �?��C�%2't �H%1p   ��8    � ��D1T�o�C�\C��M�|(E��� �@[��`&Z3���)T0 k� �;��?�%2't �H%1p   ��8    � ��D1T�g�C�TC��M�|(E��� �@W��`%Z3���'T0 k� �3��7�%2't �H%1p   ��8    � ��D1P�_�C�LC��M�|(E��� �@O��`$Z3���%T0 k� �/��3�%2't �H%1p   ��8    � ��D1P�W�C�@C���M�|(E��� ��K��`#Z3���#T0 k� �'��+�%2't �H%1p   ��8    � ��D1P�S�C�8C���]�
|(E�� ��C��`!Z3���!T0 k� �#��'�%2't �H%1p   ��8    � ��D1P�C�C�(C���]�|(E�� ��7��`Z3�q�T0 k� ����%2't �H%1p   ��8    � ��DAL�?�C�#�C���]�|(E��x�/��`Z3�q�T0 k� ����%2't �H%1p   ��8    � ��DAL�7�C��C���]�|(E��p�+��`Z3�q�T0 k� ����%2't �H%1p   ��8    � ��DAL�/�C��C�����|(E��d�#��`Z3�q�T0 k� �����%2't �H%1p   ��8    � ��DAH�'�C��C����� |(E���\���`Z3�q�T0 k� ������%2't �H%1p   ��8    � ��DAH�#�C��E������|(F ��T���`Z3�q�T0 k� ������%2't �H%1p   ��8    � ��DAH��C���EϿ����|(F �H��c`Z3�q�T0 k� ������%2't �H%1p   ��8    � 
��DAD��C���Eϳ����|(F s�4���c`Z3�q�T0 k� ������%2't �H%1p   ��8    � 	��DA@��C���Eϫ����|(F o�,���c\Z3�q�T0 k� ������%2't �H%1p   ��8    � 	��DA@���D��Eϧ����|(F g� ���c\Z3�q�T0 k� ������%2't �H%1p   ��8    � ��DA<���D��Eϟ����|,F c����c\Z3�q�	T0 k� ������%2't �H%1p   ��8    � ��DQ8 ���D��Eϛ����|,F [�����c\Z3�q�T0 k� ������%2't �H%1p   ��8    � ��DQ8!���D��Eϓ���|,F W�����c\Z3�q�T0 k� ������%2't �H%1p   ��8    � ��DQ4#���D��Eϋ���|,F S������c\
Z3�q�T0 k� ������%2't �H%1p   ��8    � ��DQ0$���E߫�Eχ���|, F O������c\Z3�q�T0 k� ������%2't �H%1p   ��8    � ��DQ,'���Eߛ�E�w���|, F G���߳�c\Z3�q��T0 k� ������%2't �H%1p   ��8    � ��DQ((���Eߓ�E�s���|, E�C���_��c\Z3�q��T0 k� ������%2't �H%1p   ��8    � ��DQ$*��Eߋ�E�k���|, E�?���_��c\Z3�q��T0 k� �����%2't �H%1p   ��8    � ��DQ +��E��E�c���|, E�;���_��c\Z3�q��T0 k� �w��{�%2't �H%1p   ��8    � ��DQ,��E�w�E�_���|, E�;��_��c\ Z3�q��T0 k� �o��s�%2't �H%1p   ��8    � ��DQ.��E�o�E�W���|, E�7��_��c_�Z3�q��T0 k� �g��k�%2't �H%1p   ��8    � ��Da/П�E�g�E�O���|, E�3��_��c_�Z3�q��T0 k� �c��g�%2't �H%1p   ��8    � ��Da1Л�E�[�E�G���!�/�E�3���_�c_�Z3�q��T0 k� �[��_�%2't �H%1p   $�8    � ��Da2Г�E�S�E�C����!�/�E�/���Ow�c_�Z3�q��T0 k� �[��_�%2't �H%1p   ��8    � ��Da6Ѓ�E�C�E�3����!�/�E�+��|Og�c[�Z3����T0 k� �K��O�%2't �H%1p   ��8    � ��Ea 7�{�E�7�E�+����!�/�E�( �tO_�c[�Z3����T0 k� �?��C�%2't �H%1p   ��8    � ��E`�9�s�E�/�E�'����!�/�Ep(OhOW�c[�Z3����T0 k� �7��;�%2't �H%1p   ��8    �  ��E`�:�k�E�#�E�����!�/�Ep$O`O�c[�Z3����T0 k� �'��+�%2't �H%1p   ��8    �  ��E`�<�c�E��E�����!�/�Ep$OXG�c[�Z3����T0 k� ����%2't �H%1p   ��8    �  ��E`�?�S�E��E�����!�/�Ep OD3�cW�Z3����T0 k� ����%2't �H%1p   ��8    �  ��E`�@�K�E���E�����!�/�Ep 
O8+�cW�Z3����T0 k� ������%2't �H%1p   ��8    ����E`�BPG�E���E������|/�Ep O0 #�cS�Z3����T0 k� ������%2't �H%1p   ��8    ����|E`�CP?�E���E�����|/�EpO( �cS�Z3����T0 k� ������%2't �H%1p   ��8    ����zE`�EP7�E���E�����|/�EpO!�cS�Z3����T0 k� ������%2't �H%1p   ��8    ����wEP�FP/�E���D.߳���|/�Ep	!�cO�Z3����T0 k� ������%2't �H%1p   ��8    ����uEP�IP�E���D.Ǵ��|/�Ep	"��cO�Z3����T0 k� ������%2't �H%1p   ��8    ����rEP�K��E���D.����|/�E`	~�".��cK�Z3����T0 k� ������%2't �H%1p   ��8    ����oEP�L��E���D.�����|/�E`	~�".��cK�Z3����T0 k� ������%2't �H%1p   ��8    ����lEP�M��E���D.�����|/�E`	~�".��cK�Z3����T0 k� ������%2't �H%1p   ��8    ����jEP�O���D���D.�����|/�E`	��#.��cG�Z3����T0 k� ������%2't �H%1p   ��8    ����hEP�P���D���D.�����|/�E`	��#.��cG�Z3����T0 k� ������%2't �H%1p   ��8    ����fEP�R���D���D.����!�/�E`!	��#.��cG�Z3����T0 k� ������%2't �H%1p   ��8    ����dEP�S���D���D.{���!�/�E`#	��#.��cC�Z3����T0 k� ������%2't �H%1p   ��8    ����bC�T���D���D.o���!�/�D0%	��#.��cC�Z3����T0 k� ������%2't �H%1p   ��8    ����`C��W�� D�s�D.[���!�/�D0 )	~�#.��c?�Z3����T0 k� �s��w�%2't �H%1p   $�8    ����]C��X�� I�k�D.O���!�/�D0 +	~�#.��S?�Z3�q��T0 k� .s��w�%2't �H%1p   ��8    ����[C��Y�I�c�D.O���!�/�D?�-	~�#>��S?�Z3�q��T0 k� .g��k�%2't �H%1p   ��8    ����YC��Z��I�[�D.K���!�/�D?�/	~�#>��S;�Z3�q��T0 k� .[��_�%2't �H%1p   ��8    ����VC��\��I�W�D.G���!�/�Eo�1	~�$>��S;�Z3�q��T0 k� .S��W�%2't �H%1p   ��8    ����TC��]��I�O�D.C�N�!�/�Eo�3Δ$>w�S7�Z3�q��T0 k� .K��O�%2't �H%1p   ��8    ����RC�t_��I�C�D.;�N�!�/�Eo�7Έ$>g�S3�Z3�q��T0 k� �;��?�%2't �H%1p   ��8    ����PC�l`��I�;�D.7�N�|/�Eo�9΀%>_�S/�Z3�q��T0 k� �3��7�%2't �H%1p   ��8    ����NC�ha��I�7�D.3�N�|/�Eo�;�x%>W�S/�Z3�q��T0 k� �+��/�%2't �H%1p   ��8    ����LC�`b�|I�/�D./���|/�Eo�=�p&>O�S+�Z3�q��T0 k� �#��'�%2't �H%1p   ��8    ����JC�\d�tI�+�D.+���|/�Eo�?�h&>O��'�Z3�a��T0 k� ����%2't �H%1p   ��8    ����HC�Pf�`I��D.#��#�|/�Eo�C�X'>?���Z3�a��T0 k� ����%2't �H%1p   ��8 	   ����GC�HgXI��E���#�|/�Eo�E�P'N?���Z3�a��T0 k� ����%2't �H%1p   ��8 	   ����FC�DhP	I��E���#�|/�Eo�G�H(N7���Z3�a��T0 k� ����%2't �H%1p   ��8 	   ����EC�<iH	I��E���#�|/�E_�I�@(N/���Z3�a��T0 k� ������%2't �H%1p   ��8 	   ����DC�8j@
I��E���#�|/�E_�K�8)N'���Z3�a��T0 k� ������%2't �H%1p   ��8 	   ����CC�(l0I���E���'�|/�E_�O�(*N���Z3�a��T0 k� ������%2't �H%1p   ��8 	   ����BC�$m(I���E���'�|/�E_�Q� *N���Z3�a��T0 k� ������%2't �H%1p   ��8 	   ����AD n I���E���'�|/�E_�R�*N����Z3�a��T0 k� ������%2't �H%1p   ��8 	   ����@D oI���E��'�|/�E_�T�+N����Z3�a��T0 k� ������%2't �H%1p   ��8 	   ����?D qI���D}��#�|/�E_�X��,M�����Z3�a��T0 k� ������%2't �H%1p   ��8 	   ����>D q Em��D}��#�|/�C�Z��,�����Z3�Q�T0 k� ������%2't �H%1p   ��8 	   ����=D�r�Em��D}��#�|/�C�[��,�����Z3�Q�T0 k� ������%2't �H%1p   ��8 	   ����<D�s�Em��D}��^#�|/�C�]��,�����Z3�Q�T0 k� ������%2't �H%1p   ��8 
   ����;D�t�Em��D}��^�|/�C�_��,�����Z3�Q�T0 k� ������%2't �H%1p   �? 
   ����:D�u�Em��O}��^�|/�C�`��-��R��Z3�Q�T0 k� ������%2't �H%1p   ��8 
   ����9D�w��Em��O}��^�|/�C�c�-&���R˿Z3�Q�T0 k� ������%2't �H%1p   ��8 
   ����8D�x��Em��O}����|/�C�|e�-&���RǿZ3�QߍT0 k� ������%2't �H%1p   ��8 
   ����8D�x�E]��O}����|/�C�xg�-&���R��Z3�QۋT0 k� ������%2't �H%1p   ��8 
   ����8D�y�E]��O}����|/�C�ph�-&���R��Z3�Q׊T0 k� ������%2't �H%1p   ��8 
   ����8D�z�E]��O}����|/�C�lj�-&���B��Z3�QӈT0 k� ������%2't �H%1p   ��8 
   ����8D�{�E]��O}����|/�C�dkm�,&���B��Z3�QφT0 k� ������%2't �H%1p   ��8 
   ����8D�|�E]��O}����|/�C�Xnmt,&���B��Z3�AǃT0 k� �s��w�%2't �H%1p   ��8    ����8D�}>�E]� O}����|/�C�Pomh,&���B��Z3�AÁT0 k� �k��o�%2't �H%1p   ��8    ����8D�~>�E]�O}����|/�C�Lqm`,&���B��Z3�A�T0 k� �g��k�%2't �H%1p   ��8    ����8D�>|E]xO}�����|/�C�DrmT,&���B��Z3�A��T0 k� �c��g�%2't �H%1p   ��8    ����8D�>pC�pO}�����|/�C�<tmL+&�{�B��Z3�A��T0 k� �[��_�%2't �H%1p   ��8    ����8C>hC�hO}�����|/�C�4umD+&�s�B�Z3����T0 k� �S��W�%2't �H%1p   ��8    ����8C>`C�`O}����|/�C�0vm8+&�o�B{�Z3����T0 k� �O��S�%2't �H%1p   ��8    ����8C�|>XC�XO}����|/�C�(xm0*&�g��s�Z3����T0 k� �G��K�%2't �H%1p   ��8    ����8C�t>PC�LO}����|/�C� y]$*&�c��k�Z3����T0 k� �@ �D %2't �H%1p   ��8    ����8C�d>@E]<O}����|/�C�|])&�S��_�Z3����T0 k� �4�8%2't �H%1p   ��8    ����8E_`>8E]4	O}��Mߛ|/�D}])&�O��W�Z3�я�T0 k� �0�4%2't �H%1p   ��8    ����8E_X~>0E],	O}��Mכ|/�D~] (&�G��O�Z3�ы�T0 k� �(�,%2't �H%1p   ��8    ����8E_P~N(E] 
O}��Mӛ|/�D�\�(&�C��K�Z3�у�T0 k� �$�(%2't �H%1p   ��8    ����8E_H~NE]O}��Mϛ|/�D��\�(&�;��C�Z3��{�T0 k� �� %2't �H%1p   ��8    ����8E_@~NE]O}��M˛|/�D��\�'&�7��;�Z3��w�T0 k� ��%2't �H%1p   ��8   ����8E_8}NE]O}��MǛ|/�E^�\�'&�/��3�Z3��o�T0 k� ��%2't �H%1p   ��8    ����8E_,}��E\�Em�����|/�E^�\�&&�'��#�Z3��c�T0 k� ��%2't �H%1p   ��8    ����8E_$}��I��Em�����|/�E^�\�&&����Z3��[�T0 k� � 	�	%2't �H%1p   ��8    ����8E_|��I��Em�����|/�E^�\�&&����Z3��S�T0 k� ��	��	%2't �H%1p   ��8    ����8EO|��I��Em�����|/�E^�~L�&&� ��Z3��O�T0 k� ��
��
%2't �H%1p   ��8    ����8EO|��I��Em�����|/�E^�~L�%&���Z3��G�T0 k� ����%2't �H%1p   ��8   ����8EN�{��I��Em�M��|, E^�~L�%&����Z3��7�T0 k� ����%2't �H%1p   ��8    ����8EN�{��I��Em{�M��|,E^�}L�%&����Z3��/�T0 k� ����%2't �H%1p   ��8    ����8EN�{�I��Emw�M��|,EN�}Lx%&����Z3��'�T0 k� ����%2't �H%1p   ��8    ����8EN�z��I��Ems�M��|,EN�}Lp%&���ߵZ3���T0 k� ����%2't �H%1p   ��8    ����8EN�z��
I��Eml M��|,EN�|Ld%���׵Z3���T0 k� ����%2't �H%1p   ��8    ����8EN�y��
I��Em`=w�|,ENt|�P%���ǴZ3���T0 k� ��
��
%2't �H%1p   ��8    ����8C��y��
I��EmX=s�|,ENl{�H%��ῴZ3����T0 k� ��	��	%2't �H%1p   ��8    ����8C��y��
I��EmP=o�|,ENd{�<%��ᷴZ3���T0 k� ��	��	%2't �H%1p   ��8    ����8C��x��
I��EmH=g�|,EN\z�4%���Z3���T0 k� ��
��
%2't �H%1p   ��8    ����8C��x��
I��Em@=c�|,ENTz�,%��	�Z3���T0 k� ����%2't �H%1p   ��8    ����8EN�w��	I�tEm4=W�|,C�@yL&��
�Z3��ӐT0 k� ����%2't �H%1p   ��8    ����8EN�v��	I�pEm,=S�|,C�8xL&̼�Z3��ːT0 k� ����%2't �H%1p   �8    ����8EN�v��	I�lEm$	=O�|,C�0xL&ܸA��Z3��ÑT0 k� ��
��
%2't �H%1p  ��?    ����8EN�u��I�hEm
=K�|,C�(wK�&ܰA�Z3��T0 k� �t�x%2't �H%1p  ��?    ����8EN�t�xI�`E]M?�|,C�vK�'ܨAo�Z3��T0 k� �`�d%2't �H%1p  $�?    ����8EN|t�tI�\E]M;�|,C�uK�'ܠAg�Z3��T0 k� ,d�h%2't �H%1p  ��?    ����8ENts�pI�XE\�M7�|,	C�tK�(�A_�Z3��T0 k� ,h�l%2't �H%1p  ��?    ����8ENls�lI�XE\�M/��,C� tK�(��W�Z3� ��T0 k� ,l�p%2't �H%1p  ��?    ����8EN`r�dI�TI��M'��,C��rK�)��G�Z3� {�T0 k� ,p�t%2't �H%1p  ��?    ����8ENXq�`I�PI��M#��,C��r;�)��?�Z3� s�T0 k� ,t�x%2't �H%1p  ��?    ����8E>Pp�\I�LI��M��,C��q;�*��7�Z3� k�T0 k� �x�|%2't �H%1p  ��?    ����8E>Lp�XI�LI��M��(C��p;�+��/�Z3� c�T0 k� �|��%2't �H%1p  ��?    ����8E>Do�TI�HI��M��(C��p;�+��'�Z3� [�T0 k� ����%2't �H%1p  ��?    ����8E><n�P I�DI��M��(C��o;�,���Z3� S�T0 k� ����%2't �H%1p   ��?    ����8E>0mmK�EL<I��M��(EM�m;x.�|��Z3� ?�T0 k� ����%2't �H%1p   ��?    ����8E>(lmG�EL8I��]��(EM�m;p/�x��Z3� 7�T0 k� <���%2't �H%1p   /�?    ����8E>$kmC�EL4I��\���(EM�l;h/�t��Z3�/�T0 k� <���%2't �H%1p   ��?    ����8E>jm?�EL0I��\���$EM�k;h0�p���Z3�'�T0 k� <���%2't �H%1p   ��?    ����8CNim;�EL,I��\���$EM�j;l1�l��Z3��T0 k� <���%2't �H%1p   ��?    ����8CNhm7�E<(I��\���$EM�i;l3�h��Z3��T0 k� <� �� %2't �H%1p   ��?    ����8CNem/�E< I��<���$EM|h+p5�`�۸Z3��T0 k� �� �� %2't �H%1p   ��?    ����8CN dm+�E<I��<���$EMtg+t6�\�ӹZ3���T0 k� �� �� %2't �H%1p   ��?    ����8CM�cm'�E<I��<���$EMlf+x7�X�˹Z3��T0 k� �� �� %2't �H%1p   ��?    ����8CM�bm�E<I��<���$C�de+x8�X�úZ3��T0 k� ������%2't �H%1p   ��?    ����8CM�`m�E<I��<��� C�\d+|:�T���Z3��T0 k� ������%2't �H%1p   ��?    ����8CM�^]�E<I��<��� C�Lb+�<�T���Z3�ϚT0 k� ������%2't �H%1p   ��?    ����8CM�]]�E<I��,��� C�Da+�>�P���Z3��ǚT0 k� ������%2't �H%1p   ��?    ����8CM�[]�E<I��,��� C�<`+�?�L���Z3�ￛT0 k� ������%2't �H%1p   ��?    ����8C]�Z]�E,I��,��� C�4_+�@�H���Z3�﷛T0 k� ������%2't �H%1p   ��?    ����8C]�Y\��E,I��,��� C�,^+�B�H���Z3�ﯛT0 k� ������%2't �H%1p   ��?    ����8C]�V\��E+�I��,��� C�]�E�@��Z3�O��T0 k� ������%2't �H%1p   ��    ����8C]�U	���E+�Eܐ,��� C�\�F�<�w�Z3�O��T0 k� ������%2't �H%1p   ��    ����8I]�S	���E+�E܌,��� E�[�G�8�s�Z3�O��T0 k� ������%2't �H%1p   ��    ����8I]�R	���E+�E܌,��� E�Z�I�8�k�Z3�O��T0 k� ������%2't �H%1p   ��    ����8I]�P	���E+�E܈����E��X��K�8�[�Z3�Os�T0 k� ������%2't �H%1p   �    ����8I]�N	���fK�E����| E��W��M�4�S�Z3�Ok�T0 k� ������%2't �H%1p   ��    ����8E=�M	���fK�E����|  EL�V��N�4�K�Z3�Oc�T0 k� ������%2't �H%1p   ��    ����8E=�J	���fK�E�|���|#�EL�S��P�4�?�Z3��O�T0 k� ������%2't �H%1p   ��    ����8E=�I	���fK�E�x̛�|#�EL�R��R�0�7�Z3��G�T0 k� ������%2't �H%1p   ��    ����8E=�G	���fK�D�x̗�|#�EL�Q��S�0�/�Z3��?�T0 k� ������%2't �H%1p   ��    ����8E=�F	���fK�D�t̓��#�I|�P��T�0�'�Z3��7�T0 k� ������%2't �H%1p   ��    ����8E=�C	���fK�D�p̋��#�I|�O��V�0��Z3��'�T0 k� ������%2't �H%1p   ��    ����8E=�A	���f[�D�l̇��'�I|�N��W�0��Z3���T0 k� ������%2't �H%1p   ��    ����8E=�@	���f[�D�l���'�I|�M��Y�0��Z3���T0 k� ������%2't �H%1p   ��    ����8E-�>\��f[�D�l�{��'�I|�L��Z�0��Z3���T0 k� ������%2't �H%1p   ��    ����8E-x;\��f[�D�h�s��'�EL�J�\�0���Z3����T0 k� ������%2't �H%1p   ��    ����8E-x9\��f[�BLd�o��'�EL�J�]�0���Z3���T0 k� ������%2't �H%1p   ��    ����8E-t7\��f[�BLd �g��'�EL�I�^�0���Z3���T0 k� ������%2't �H%1p   ��    ����8E-p6��fk�BLd �c��'�EL�H� _�0���Z3���T0 k� ������%2't �H%1p   ��    ����8E-l2��fk�BL` �c��#�E<tF�0a�0���Z3��өT0 k� ������%2't �H%1p   ��    ����8E-l1��fk�F`!�c�|�E<lD�8b�0���Z3��˪T0 k� ������%2't �H%1p   ��    ����8E-h/��fk�F`!�c�|�E<hC�@c�0���Z3��êT0 k� ������%2't �H%1p   ��    ����8E-h- ���fk�F`"�_�|�E<`B�Hd�0���Z3����T0 k� ������%2't �H%1p   ��    ����8E-d) ���fk�F`"�_�|�E<T?�Xf�0���Z3����T0 k� ������%2't �H%1p   ��    ����9Ed( ���fk�E�`#�[�|�E<P>�dg�0
ߧ�Z3�	~��T0 k� ������%2't �H%1p   ��    ����:Ed& ���f[�E�`#�[�|�E<H=�lh�0
ߟ�Z3�	~��T0 k� ������%2't �H%1p   ��    ����;E`$ l��f[�E�`#�W�|�E<D;�ti0
ߗ�Z3�	~��T0 k� ������%2't �H%1p   �    ����<E`# l��f[�E�d$�W�|�E<<9�|j,
ߓ�Z3�	~��T0 k� ������%2't �H%1p   ��    ����=E`! l��f[�E�d$�W�|�E,88̈k,ߋ�Z3�	~��T0 k� ������%2't �H%1p   ��    ����>Ed l��f[�E�h%LS�|�E,05̘m$�{�Z3�	~w�T0 k� ������%2't �H%1p   ��    ����?Ed l��f[�E�h%LS�|�E,(3ܠn�$�s�Z3�	�s�T0 k� ������%2't �H%1p   ��    ����@Ed ��fK�E�l%LP |�E,$1ܨn� �o�b��	�k�T0 k� ������%2't �H%1p   ��    ����AEd ��fK�E�l%LP|�E, 0ܴo� �g�b��	�g�T0 k� ����%2't �H%1p   ��    ����BEd ��fK�E�p%LP|�B�.ܼp��_�b��	�_�T0 k� ����%2't �H%1p   ��    ����CEh ��fK�CLp%LP|�B�,��q��W�b��	�[�T0 k� ����%2't �H%1p   ��    ����DE�h ��fK�CLt%LP|�B�+��r��O�b��NW�T0 k� ����%2't �H%1p   ��    ����EE�l ,��fK�CLx%LL|�B�'��s��C�b��NK�T0 k� �#��'�%2't �H%1p   ��    ����FE�p ,��fK�CLx%LL|�E,'��t�O;�b��NC�T0 k� �+��/�%2't �H%1p   ��    ����HE�p ,��@�CLx$LL|�E,&��u�O3�b��N?�T0 k� �/��3�%2't �H%1p   ��    ����JD�t ,��@�CL|$LL|�E,$�v�O#�b��>3�T0 k� �7��;�%2't �H%1p   ��    ����LD�x ,��@�CL�#LL|�E,#�w�O�Z3�>+�T0 k� �;��?�%2't �H%1p   ��    ����ND�| ,��@�CL�#LL|�E,"�x�O�Z3�>'�T0 k� �C��G�%2't �H%1p   ��    ����PD�|
 <��B��CL�"LH	|�E,!� y�O�Z3�>�T0 k� �K��O�%2't �H%1p   ��    ����RE�� <��B��CL�!LH
|�B�$�4z�N��Z3�>�T0 k� �S��W�%2't �H%1p   ��    ����TE�� <��B��C\� LH
|�B�,�<{�N��Z3�>�T0 k� �[��_�%2't �H%1p   ��    ����VE�� <��B��C\�LH|�B�0�D{� >��Z3�>�T0 k� �_��c�%2't �H%1p   ��    ����XE�� <��B��C\�LH|�B�0�P|� >��Z3�>�T0 k� �c��g�%2't �H%1p   �    ����ZE�� =�B��C\��H|#�O�8�`}��>��Z3�=��T0 k� �k��o�%2't �H%1p   ��    ����\E�� =�B��C\��H|#�O�@�l~��>��Z3�=��T0 k� �o��s�%2't �H%1p   ��    ����^E�� =�B��C\��H
|#�O�D�t��>��bs�=��T0 k� ������%2't �H%1p   �    ����iE}�M�B��C\��L
|#�O�H�|��>��bs�-��T0 k� ������%2't �H%1p   ��    ����tE}�M�B��C\��L
|#�O�L�����>��bs�-��T0 k� ������%2't �H%1p   ��    ����~E}�M�B��C\��L	|'�O�T�����>��bs�-��T0 k� ������%2't �H%1p  ��    �����E}�M#�B��Cl��L	|'�O�\����>��bs�-��T0 k� ������%2't �H%1p  ��    �����D��M#�B��Cl��L	|'�O�\�� >��bs�-��T0 k� ������%2't �H%1p  ��    �����D��]'�B��Cl��L|'�O�`�� >��bs�-��T0 k� ����%2't �H%1p  ��    �����D��]+�B��Cl��L|'�O�d�� .��bs�-��T0 k� ����%2't �H%1p  ��    �����D��]/�B�� Cl��L|'�O�h�~� .��bs�-��T0 k� �/��3�%2't �H%1p  ��    �����D��]3�B�� Cl��P|'�O�l�~� .��bs�-��T0 k� �?��C�%2't �H%1p  ��    �����D��]7�B�� Cl��P|'�O�p�~� .��Z3�-��T0 k� �S��W�%2't �H%1p  ��    �����D��m;�B� I\��P|'�O�t�~� .��Z3�-��T0 k� �g��k�%2't �H%1p  ��    �����D��m;�B� I\�
�P|'�O�t�}� .��Z3�-��T0 k� �w��{�%2't �H%1p  ��    �����F�m?�B�!I\�	�P|'�O�x�}�.� Z3���T0 k� ������%2't �H%1p  ��    �����F�mC�B�!I\��P|'�O�|�}�.|Z3���T0 k� ������%2't �H%1p  ��   �����F�mG�B�!I\��P|'�O���}�.xZ3���T0 k� ������%2't �H%1p  ��    �����F�mG�B�!I\��P|'�O���|�.tZ3���T0 k� ������%2't �H%1p  ��    �����F�mK�B� !Il��P|'�O��� |�tZ3���T0 k� ������%2't �H%1p  ��    �����E��mO�B�(!Il��T|'�O���(|�pZ3���T0 k� ������%2't �H%1p  ��    ��� E��mS�B�,"Il��T|'�O���4{�lZ3���T0 k� �����%2't �H%1p  ��    ��� 	E��mS�B�4"Il��T|'�O���<{�h
Z3����T0 k� ����%2't �H%1p  ��    ��� E��mW�B�8"Il��T|'�O���Hz�hZ3����T0 k� �#��'�%2't �H%1p  ��    ��� E��m[�B�@"I\� �T|'�O���Pz��dZ3����T0 k� �7��;�%2't �H%1p  ��    ��� B��m[�B�D"I\���T|'�E,��Xy��`Z3����T0 k� �G��K�%2't �H%1p   ��    ��� "B��m_�B�L"I\���T|'�E,��dy��`Z3����T0 k� �[��_�%2't �H%1p   ��    ��� (B��mc�B�T#I\���T|'�E,��lx��\Z3����T0 k� �o��s�%2't �H%1p   ��    ��� .B��mc�B�\#I\���T|'�E,��tw��\Z3����T0 k� ������%2't �H%1p   /�    ��� 4B��mg�B�`#Il���T|'�E,�ހw��\Z3����T0 k� ������%2't �H%1p   ��   ��� :B��mk�B�h#Il���X|'�E�ވv��XZ3����T0 k� ������%2't �H%1p   ��    ��� @B��mk�B�p#Il���X|'�E�ސv��XZ3����T0 k� ������%2't �H%1p   ��    ��� FB� mo�B�x#Il���X|'�E�ޜu��XZ3����T0 k� ������%2't �H%1p   ��    ��� LB�mo�B܀$Il���X|'�E�ޤt��TZ3����T0 k� ������%2't �H%1p   ��    ��� QB��s�B��$I\���X|'�E�ެt��TZ3����T0 k� ������%2't �H%1p   ��    ��� VB��w�B��$I\���X|'�B��޸s��TZ3����T0 k� ����%2't �H%1p   ��    ��� [B��{�B��$I\���X|'�B����r��TZ3����T0 k� ����%2't �H%1p   ��    ��� `B��{�B��$I\���X|'�B����q�.T Z3����T0 k� �'��+�%2't �H%1p   ��    ��� eB���B��%I\���X|'�B����p�.T!Z3����T0 k� �;��?�%2't �H%1p   ��    ��� jB�$���B��%E,���\|'�B����p�.P#Z3����T0 k� �O��S�%2't �H%1p   ��    ��� oB�(���B��%E,���\|'�B����o�.P%Z3����T0 k� �_��c�%2't �H%1p   ��    ��� tB�0���B��%E,���\|'�B����n�.T&Z3����T0 k� �s��w�%2't �H%1p   ��    ��� yB�4���B��&E,���\|'�B����m�T(Z3����T0 k� ������%2't �H%1p   ��    ��� ~B�<���B��&E,���\|'�B��� l�T)Z3����T0 k� ������%2't �H%1p   ��   ��� �B�@���B��&E���`|'�B��k�T*Z3����T0 k� ������%2't �H%1p   ��    ��� �B�H���B��&E���`|'�B��k�T,Z3����T0 k� ������%2't �H%1p   ��    ��� �B�P���B��&E���`|'�B��j�X-Z3����T0 k� ������%2't �H%1p   ��    ��� �B�T���B��'E���`|'�B��$i��X/Z3����T0 k� ������%2't �H%1p   ��   ��� �B�\���B��'E���`|'�B�$�,h��X0Z3����T0 k� ������%2't �H%1p   ��    ��� �B�d���B��'E���`|'�B�,�8g��\1Z3����T0 k� ����%2't �H%1p   ��    ��� �B�l���B�'E���d|'�B�4�@f��\3Z3���T0 k� ����%2't �H%1p   ��    ��� �B�p���B�(E���d|'�B�<�He��`4Z3���T0 k� �'��+�%2't �H%1p   ��    ��� �B�x���B�(E���d|'�B�D�Pd��`5Z3���T0 k� �;��?�%2't �H%1p   ��    ��� �B΀���B�$(E���d|+�B�L�Xc��d7Z3��#�T0 k� �K��O�%2't �H%1p   ��    ��� �BΈ���B�,(E���d|+�B�T�db��d8Z3��, T0 k� �_��c�%2't �H%1p   ��    ��� �Bΐ��B�4(E����d|+�B�`�la��h9Z3��8T0 k� �o��s�%2't �H%1p   ��    ��� �BΘ��B�@)E����h|+�B�h�t`�l:Z3��DT0 k� �����%2't �H%1p   �    ��� �E����B�H)E����h|+�@pO|_�l;Z3� �PT0 k� ������%2't �H%1p   �    ��� �E����B�T)E����h|+�@xO�^�p=Z3� �XT0 k� ������%2't �H%1p   ��    ��� �E����B�\)E����h|+�@�O�]�t>Z3� �dT0 k� ������%2't �H%1p   ��    ��� �E����B�d)E����h|+�@�O�\�x?Z3� �pT0 k� ������%2't �H%1p   ��    ��� �E����B�p*E����h|+�@�O�[�|@Z3���xT0 k� ������%2't �H%1p   ��    ��� �E����B�x*E����h|+�@�O�Z��AZ3����T0 k� ������%2't �H%1p   ��    ��� �E���B̈́*E����l|+�@�O�Y��BZ3����T0 k� ������%2't �H%1p   ��    ��� �E���B͌*E����l|+�@�O�X��CZ3���T0 k� ����%2't �H%1p   ��    ��� �E����B͔*E����l|+�@�O�W��DZ3���T0 k� ���#�%2't �H%1p   ��    ��� �E����B͠*E����l|+�@�O�V���EZ3���T0 k� �/��3�%2't �H%1p   ��    ��� �B����Bͨ+B���l|+�@�O�U���FZ3���T0 k� �C��G�%2't �H%1p   ��    ��� �B��#�Bݰ+B���l|+�@�O�U���GZ3���	T0 k� �S��W�%2't �H%1p   ��    ��� �B��+�Bݼ+B���l|+�@�O�T���HZ3���	T0 k� �c��g�%2't �H%1p   ��    ��� �B�  �3�B��+B���p|+�@�O�S���IZ3���
T0 k� �w��{�%2't �H%1p   ��    ��� �B�/��;�B��+B���p|+�@�O�R���JZ3���
T0 k� ������%2't �H%1p   ��    ��� �B�;��C�B��+B���p|+�@�O�Q���JZ3���T0 k� ������%2't �H%1p   ��    ��� �B�G��K�B��+B�'��p|+�@�O�P���KZ3���T0 k� ������%2't �H%1p   ��    ��� �B�O��S�B��,B�+��p|+�@�O�P���LZ3���T0 k� ������%2't �H%1p   ��    ��� �B�[��[�B��,B�3��p|+�@�@ O���LZ3���T0 k� ������%2't �H%1p   ��    ��� �B�g��c�B��,B�7��p|+�@�@N�N�MZ3���T0 k� ������%2't �H%1p   ��    ��� �B�s��k�B�,B�?��p|+�@ �M�N�MZ3���T0 k� ������%2't �H%1p   ��    ��� �B�{��s�B�,B�G��t|+�@�M�N�NZ3���T0 k� �����%2't �H%1p   ��    ��� �B���{�B�,B�O��t|+�@�L�N�NZ3���T0 k� ����%2't �H%1p   ��    ��� �B�����B�$,B�S��t|+�@� K�N�OZ3��T0 k� �#��'�%2't �H%1p   ��    ��� �B�����B�,-B�[��t|+�@�(J�N�OZ3��T0 k� �3��7�%2't �H%1p   ��    ��� �B�����B�8-B�c��t|+�@ �0I�N�PZ3��T0 k� �C��G�%2't �H%1p   ��    ��� �B�����B�@-B�k��t|+�@$�4H�N�PZ3��T0 k� �S��W�%2't �H%1p   ��    ��� �B�����B�L-B�s��t|+�@,�<H�N�QZ3��T0 k� �g��k�%2't �H%1p   ��    ��� �B������B�T-B�{��t|+�@0�@G�N�QZ3��$T0 k� �w��{�%2't �H%1p   ��    ��� �B������B�\-B����t|+�@4�HF�N�RZ3��(T0 k� ������%2't �H%1p   ��    ��� �B������B�h-B����x|+�@<@LE�N�RZ3��0T0 k� ������%2't �H%1p   ��    ��� �B������B�p.B����x|+�@@@TE�N�SZ3��4T0 k� ������%2't �H%1p   ��    ��� �B������B�x.B����x|+�@D@XD�N�SZ3��<T0 k� ������%2't �H%1p   ��    ��� �B������B��.Bͣ��x|+�@L@\C�N�TZ3�� @T0 k� ������%2't �H%1p   ��    ��� �E�����B��.Bͫ��x|+�@P@dCN�TZ3�� HT0 k� ������%2't �H%1p   ��    ��� �E�����B��.Bͳ��x|+�@T@hBN�UZ3�� LT0 k� ������%2't �H%1p   ��    ��� �E����B��.Bͻ��x|+�@X@lAO UZ3�� PT0 k� ������%2't �H%1p   ��    ��� �E����B��.B����x|+�@\@t@OVZ3�� XT0 k� ����%2't �H%1p   ��    ��� �E���B��.B����x|+�@d@x@OVZ3�� \T0 k� ����%2't �H%1p   ��    ��� �E#���E��.B����x|+�@h@|?OVZ3�� `T0 k� �/��3�%2't �H%1p   ��    ��� �E+���E��.B����x|+�@l@�?OWZ3�� hT0 k� �?��C�%2't �H%1p   ��    ��� �E3���E��.B����||+�@p@�>OWZ3�� lT0 k� �O��S�%2't �H%1p   ��    ��� �E7��#�E��.B����||+�@t@�=OXZ3�� pT0 k� �_��c�%2't �H%1p   ��    ��� �E?��+�E��.B����||+�@x@�=�OXZ3�� tT0 k� �o��s�%2't �H%1p   ��    ��� �B�G��3�E��-B����||+�@|@�<�OXZ3�� xT0 k� �����%2't �H%1p   ��    ��� �B�O��?�E��-B���||+�@�@�;�OYZ3�� �T0 k� ������%2't �H%1p   ��    ��� �B�W��G�B� -B���||+�@�@�;�O YZ3�� �T0 k� ������%2't �H%1p   (�    ��� �B�_��O�B�-B���||+�@�@�:�O$ZZ3�� �T0 k� 4�����%2't �H%1p   -�    ��� �B�c��W�B�,B�#��||+�@�@�:�O$ZZ3�� �T0 k� 4�����%2't �H%1p   ��    ��� �@k��_�B�,B�+��||+�@�@�9�O(ZZ3�� �T0 k� 4�����%2't �H%1p   ��    ��� �@s��g�B�$+B�7��||+�@�@�9�O,[Z3�� �T0 k� 4�����%2't �H%1p   ��    ��� �@w��o�B�0+B�?��||+�@�@�8�O,[Z3�� �T0 k� 4�����%2't �H%1p   ��    ��� �@��w�B�8+B�G��||+�@�@�8LO0[Z3�� �T0 k� ������%2't �H%1p   ��    ��� �@����B�@*B�O��||+�@�@�7LO4\Z3�� �T0 k� ������%2't �H%1p  ��   ��� �K������B�L*B�W���|+�@�@�7LO4\Z3�� �T0 k� �����%2't �H%1p  ��    ��� �K������B�T)B�_���|+�@�@�6LO8\Z3�� �T0 k� �{���%2't �H%1p  ��    ��� �K������B�\)B�k���|+�@�@�6LO<]Z3�� �T0 k� �w��{�%2't �H%1p  ��    ��� �K������B�h(B�s���|+�@�@�5LO<]Z3�� �T0 k� �s��w�%2't �H%1p  ��    ��� �K������Cp'B�{��|+�@�@�5LO@]Z3�� �T0 k� �o��s�%2't �H%1p  ��    ��� �K������Cx'B����|+�@�@�4LOD^Z3�� �T0 k� �k��o�%2't �H%1p  ��    ��� �K������C�&B����|+�@�@�4LOD^Z3�� �T0 k� �g��k�%2't �H%1p  ��    ��� �K������C�&B����|+�@�@�3LOH^Z3�� �T0 k� �c��g�%2't �H%1p  ��    ��� �K������C�&B����|+�@�@�3LOH^Z3�� �T0 k� D_��c�%2't �H%1p   ��    ��� �K������C�%B����|+�@�@�2LOL_Z3�� �T0 k� D[��_�%2't �H%1p   ��   ��� �K������C�%B����|+�@�@�2LOP_Z3�� �T0 k� DW��[�%2't �H%1p   ��    ��� �K������C�%B����|+�@�@�1LOP_Z3�� �T0 k� DS��W�%2't �H%1p   ��    ��� �K������C�%B����|+�@�@�1LOT`Z3�� �T0 k� DO��S�%2't �H%1p   ��    ��� �K������C�$B���L�|+�@�@�1LOT`Z3�� �T0 k� $K��O�%2't �H%1p   ��    ��� �K������C�$B���L�|+�@�@�0LOX`Z3�� �T0 k� $G��K�%2't �H%1p   /�   ��� �K�����C�$B���L�|+�@�@�0LOX`Z3�� �T0 k� $C��G�%2't �H%1p   ��    ��� �K�����C�#B���L�|+�@�@�/LO\aZ3�� �T0 k� $?��C�%2't �H%1p   ��    ��� �K�����C�#B���L�|+�@�@�/LO\aZ3�� �T0 k� $;��?�%2't �H%1p   ��    ��� �K����#�C�#B���L�!�+�@�A /LO`aZ3�� T0 k� �7��;�%2't �H%1p   ��    ��� �K����+�C�"B���L�!�+�@�A .L O`aZ3�� T0 k� �3��7�%2't �H%1p   ��   ��� �K����3�C�"B��L�!�+�@�A.L OdbZ3�� T0 k� �/��3�%2't �H%1p   ��    ��� �K����;�C�"B��L�!�+�@�A.L OdbZ3�� T0 k� �+��/�%2't �H%1p   ��    ��� �K���C�C�"B���!�+�@�A-L OhbZ3�� T0 k� �'��+�%2't �H%1p   ��    ��� �K���K�C�!B���!�+�@�A-L OhbZ3��  T0 k� �#��'�%2't �H%1p   ��    ��� �K���S�C�!B�+��!�+�@�A-L OlcZ3�� $T0 k� ���#�%2't �H%1p   ��    ��� �K���[�C� B�3��!�+�@�A,L OlcZ3�� ,T0 k� ����%2't �H%1p   ��    ��� �K���g�C/� B�;��!�+�@�A,L OpcZ3�� 0T0 k� ����%2't �H%1p   ��    ��� �K���o�C/� B�C� ��!�+�@�A,L OpcZ3�� 8T0 k� ����%2't �H%1p   ��    ��� �K���w�C/� B�K� ��!�+�@�A+L OpcZ3�� <T0 k� ����%2't �H%1p   ��    ��� �K����C  B�W� ��|+�@�A+L OtdZ3�� DT0 k� ����%2't �H%1p   ��    ��� �K�#���C B�_� ��|+�@�A +L OtdZ3�� HT0 k� ����%2't �H%1p   ��    ��� �K�'���C B�g� ��|+�@ A *L OxdZ3�� PT0 k� ����%2't �H%1p   ��    ��� �K�+���C B�o� l�|+�@ A$*L OxdZ3�� TT0 k� ����%2't �H%1p   ��    ��� �K�/���C B�w� l�|+�@A(*L O|dZ3�� \T0 k� �����%2't �H%1p   ��    ��� �K�3���C  Bσ� l�|+�@A()L O|eZ3�� `T0 k� ������%2't �H%1p   ��    ��� �K�7���C (K��� l�|+�@A,)L O|eZ3�� dT0 k� ������%2't �H%1p   $�    ��� �K�;���C ,K��� l�|+�@A,)L O�eZ3�� lT0 k� ������%2't �H%1p   ��
    ��� �K�;���B�4K�����|+�@A0(L O�eZ3�� pT0 k� ������%2't �H%1p   ��
    ��� �K�?����B�4K�����|+�@A0(L O�eZ3�� xT0 k� ������%2't �H%1p   ��
    ��� �K�C����B�8K�����|+�@A4(L O�fZ3�� |T0 k� ������%2't �H%1p   ��
    ��� �K�G����B�@K�����!�+�@A4(L O�fZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�K����B�DK�����!�+�@A8'L O�fZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�O����B�LK�����!�+�@A<'L O�fZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�O����B�PK�����!�+�@A<'L O�fZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�S����B�XK�����!�+�@A@'L O�gZ3�� �T0 k� ������%2't �H%1p   ��
   ��� �K�W���B�\K�����!�+�@A@&L O�gZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�[���K�dK�����!�+�@AD&L O�gZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�_���K�hK�����!�+�@ AD&L O�gZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�_���K�hK�����!�+�@ AD&L O�gZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�c��'�K�lK�����!�+�@ AH%L O�gZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�g��/�K�pK�����!�+�@$AH%L O�gZ3�� �
T0 k� ������%2't �H%1p   ��
    ��� �K�k��7�K�xK����|+�@$AL%L O�hZ3�� �
T0 k� ������%2't �H%1p   ��
    ��� �K�k��?�K�|K����|+�@(AL%L O�hZ3�� �	T0 k� ������%2't �H%1p   ��
    ��� �K�o��G�K��K����|+�@(AP%L O�hZ3�� �	T0 k� ������%2't �H%1p   ��
    ��� �K�s��S�K��K����|+�@(AP$L O�hZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�s��[�K��K����|+�@,AT$L O�hZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�w��c�K��K�#���|+�@,AT$L O�hZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�{��k�K��K�+���|+�@0AT$L O�iZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K�{��s�K��K�/���|+�@0AX$L O�iZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K���{�K��
K�7���|+�@0AX#L O�iZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �@���K��	K�;���|+�@4A\#L O�iZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �@����K��	K�C���|+�@4A\#L O�iZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �@����K��K�G���|+�@4A\#L O�iZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �@����K��K�K���|+�@8A`#L O�iZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �@����K��K�S���|+�@8A`"L O�iZ3��  T0 k� ������%2't �H%1p   ��
    ��� �@����K��K�W���|+�@8Ad"L$O�jZ3�� T0 k� ������%2't �H%1p   ��
    ��� �@����K��K�[���|+�@<Ad"L$O�jZ3�� T0 k� ������%2't �H%1p   ��
    ��� �@����K��K�c���|+�@<Ad"L$O�jZ3�� T0 k� ������%2't �H%1p   ��
    ��� �@��q��K��K�g���|+�@<Ah"L$O�jZ3�� T0 k� ������%2't �H%1p   ��
    ��� �@��q��K��K�k���|+�@@Ah"L$O�jZ3�� T0 k� ������%2't �H%1p   ��
    ��� �@��q��K��K�s���|+�@@Ah!L$O�jZ3�� T0 k� ������%2't �H%1p   ��
    ��� �@��q��K��K�w���|+�@@Al!L$O�jZ3�� T0 k� ������%2't �H%1p   ��
    ��� �@��q��K��K�{���|+�@DAl!L$O�jZ3��  T0 k� ������%2't �H%1p   ��
    ��� �@��q��K��K����|+�@DAl!L$O�jZ3�� $T0 k� ������%2't �H%1p   ��
    ��� �@��q��K��K�����|+�@DAp!L$O�kZ3�� (T0 k� ������%2't �H%1p   ��
   ��� �@��q��K��K�����|+�@HAp!L$O�kZ3�� , T0 k� ������%2't �H%1p   ��
    ��� �@��q��K�� K�����|+�@HAp L$O�kZ3�� 0 T0 k� ������%2't �H%1p   ��
    ��� �@��r�K�� K�����|+�@HAp L$O�kZ3�� 4 T0 k� ������%2't �H%1p   ��
    ��� �@��r�K���K�����|+�@HAt L$O�kZ3�� ;�T0 k� ������%2't �H%1p   ��
    ��� �@����K���K�����|+�@LAt L$O�kZ3�� ?�T0 k� ������%2't �H%1p   ��
    ��� �@����K���K�����|+�@LAt L$O�kZ3�� ?�T0 k� ������%2't �H%1p   ��
    ��� �@����K���K�����|+�@LAx L$O�kZ3�� C�T0 k� ������%2't �H%1p   ��
    ��� �@���#�K���K�����|+�@LAx L$O�kbs�� G�T0 k� ������%2't �H%1p   ��
    ��� �@���'�K���K�����|+�@PAxL$O�lbs�� K�T0 k� ������%2't �H%1p   ��
    ��� �K����+�K���K�����|+�@PAxL$O�lbs�� O�T0 k� ������%2't �H%1p   ��
    ��� �K����3�K��K�����|+�@PA|L$O�lbs�� S�T0 k� ������%2't �H%1p   ��
    ��� �K����7�K��K�����|+�@PA|L$O�lbs�� S�T0 k� ������%2't �H%1p   ��
    ��� �K����?�K��K�����|+�@TA|L$O�lbs�� W�T0 k� ������%2't �H%1p   ��
    ��� �K����C�K��K�����|+�@TA�L$O�lbs�� [�T0 k� ������%2't �H%1p   ��
   ��� �K����K�K��K�����|+�@TA�L$O�lbs�� _�T0 k� ������%2't �H%1p   ��
   ��� �K����O�K��K�����|+�@TA�L$O�lbs�� _�T0 k� ������%2't �H%1p   ��
    ��� �K����[�K��K�����|+�@XA�L$O�lbs�� g�T0 k� ������%2't �H%1p   ��
    ��� �K����_�K��K�����|+�@XA�L$O�lZ3�� k�T0 k� ������%2't �H%1p   ��
    ��� �K����c�K��K�����|+�@XA�L$O�lZ3�� k�T0 k� ������%2't �H%1p   ��
    ��� �K����g�K��K�����|+�@XA�L$O�mZ3�� o�T0 k� ������%2't �H%1p   ��
    ��� �K����o�K��B�����|+�@\A�L$O�mZ3�� s�T0 k� ������%2't �H%1p   ��
    ��� �K����s�K�#�B�����|+�@\A�L$O�mZ3�� s�T0 k� ������%2't �H%1p   ��
    ��� �K����w�K�'�B�����|+�@\A�L$O�mZ3�� w�T0 k� ������%2't �H%1p   ��
    ��� �K����{�K�'�B�����|+�@\A�L$O�mZ3�� {�T0 k� ������%2't �H%1p   ��
    ��� �K�����K�+�B�����|+�@`A�L$O�mZ3�� {�T0 k� ������%2't �H%1p   ��
    ��� �K������K�+�B�����|+�@`A�L$O�mZ3�� �T0 k� ������%2't �H%1p   ��
    ��� �K������K�/�B�����|+�@`A�L$O�mZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K������K�3�E�����|+�@`A�L$O�mZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K������K�3�E�����|+�@`A�L$O�mb��� ��T0 k� ������%2't �H%1p   ��
    ��� �K������K�7�E����|+�@`A�L$O�mb��� ��T0 k� ������%2't �H%1p   ��
   ��� �K������K�7�E����|+�@dA�L$O�mb��� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�;�E����|+�@dA�L$O�mb��� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�;�E����|+�@dA�L$O�nb��� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�?�E����|+�@dA�L$O�nb��� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�C�E����|+�@dA�L$O�nb��� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�G�E����|+�@hA�L$O�nb��� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�K�E����|+�@hA�L$O�nb��� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�S�E����|+�@hA�L$O�nb��� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�W�E�'���|+�@hA�L$O�nb��� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�[�E�+���|+�@hA�L$O�nZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�_�E�/���|+�@hA�L$O�nZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�_�B�7���|+�@hA�L$O�nZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K������B�c�B�;���|+�@lA�L$O�nZ3�� ��T0 k� ������%2't �H%1p   ��
   ��� �K������Cg�B�?���|+�@lA�L$O�nZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K���r��Ck�B�?���|+�@lA�L$O�nZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K���r��Co�B�C���|+�@lA�L$O�nZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K���r��Cs�B�G�� |+�@lA�L$O�nZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K���r��Cw�B�O��|+�@lA�L$O�nZ3�� ��T0 k� ������%2't �H%1p   ��
   ��� �K���r��C�B�S��|+�@pA�L$O�oZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K���r��C��C[��|+�@pA�L$O�oZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K������C��C_��|+�@pA�L$O�oZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K������C��Cc��|+�@pA�L$O�oZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K������C��Ck��|+�@pA�L$O�oZ3�� ��T0 k� ������%2't �H%1p   ��
   ��� �K������C��Co��|+�@pA�L$O�oZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �K������C��Cw�� |+�@pA�L$O�oZ3�� ��T0 k� ������%2't �H%1p   ��
    ��� �EqBC�C�H<C����9|(E���ќp��`;Z3��XT0 k� ������%2't �H%1p   ��8    � +  EqB?�C�@:C����8|(E���јp��`;Z3��WT0 k� ������%2't �H%1p   ��8    � +  EqB3�C�07C��}�6|(E���ѐp��`;Z3��UT0 k� ������%2't �H%1p   �8    � +  EqB/�C�,5C��}�5|(E����`��`;Z3�� TT0 k� �����%2't �H%1p   ��8    � +��Eq B'�C�$4C��}�4|(Eѻ��`��`;Z3���ST0 k� �����%2't �H%1p   ��8    � +��D�$B#�E�2C��}�4|(Eѳ��`��`;Z3���RT0 k� �����%2't �H%1p   ��8    � +��D�$B�E�0C��}�3|(Eѫ��|`��`:Z3���QT0 k� �����%2't �H%1p   ��8    � +��D�,��E�-C��}�1|(E���p`��`:Z3���NT0 k� �����%2't �H%1p   ��8    � *��D�,��E�+C��}�/|(E���l`� �`9Z3���MT0 k� ������%2't �H%1p   ��8    � )��D�0��E��*C��}�.|(E���d`���`9Z3���LT0 k� ������%2't �H%1p   ��8    � (��D�4���E��(C��}�-|(E���``���`9Z3��JT0 k� ������%2't �H%1p   ��8    � '��D�4���E��&C��m�,|(E���XP���`8Z3��IT0 k� ������%2't �H%1p   ��8    � &��D�8��E��%C��m�+|(E�{��TP���`8Z3��GT0 k� ������%2't �H%1p   ��8    � %��D�<��E��!C��m�(|(E�k��DP���`6Z3��ET0 k� ������%2't �H%1p   ��8    � $��                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \���� ]�' &� � �����  � �
     � z��    ��#o zL�    ��;             c �� �           �    ���   0	          �Ǣ)   M M     � �D�    ��	� �Zs    �Ra               q�� �         H�b     ���  @
"	         ��D  1 1      f�[    ���� e}�    �+             #�� �         ��  	  ���   		'          �م+  0 0        ]`�    �ځ. [�     ��2              �� �          �p�    ���   8	
           &u   ,
	    .�H��     &u�Gy�      B              / �� �           ��  	  ���  X	
         ��}�  ��	      B�
)    ��}��
)                          �����              �  ���    00
           #�  �
     V���     #��ܬg      �                 �          p     ��@   (
           ��  $ $     j hd     � g��    �             � �         ��     ��@   8�		          g"  $/
   ~�	|n     f�	|n                    	    � $          bp     ��B   0

 
 
          oWB  $ $     ���F�     oJO��.�     �n             
     Y         	 P     ��B   P
B 
         ��(��     � ���    ��( ���                              �� �       
      �  ��H    8		 1 	            ���          � q�\    ��� p�b    �	Z                �� �          �     ��@   (
                 ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��.  ��        � �`�    ��. �`�                          x                j  �    
   �                         ��    ��        � �      ��   �           "                                                 �                          z � f ]�H�
�� h�	�� � q�� � � 
           	     
  �   it� ~ �K        ``� � a� � a� ��  _� Є _� Ф _� 
�< W� 
�\ W� �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À���� ����� ����� ����� � 
�< W� 
�� W� 
�\ W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���� � �����C  ������  
�fD
��L���"����D" � j  "  B   J jF�"     "�j  " ��
��
��"    B�j l �  B �
� �  �  
� ��   ��     � �      ��    ��     � z      ��   ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �
 1 1      �� �T ���        �*T ���        �        ��        �        ��        �     ��    ��������        ��                         T�) , ��� �                                     �                 ����            
�� �
���%��  �� � 2               16 Pat LaFontaine y    5:21                                                                        2  2     �8K �/K �G K �G K �+cj; cr#c� �J� �	J� � �
J� � �B� � � � � �k� � �k� � �k� � � k� � �	� � �	�  �� � �� �"� � � "� � �� � �
� �>"� �> "� �."� �.*� � �"� � � "� � �� � � 
� � �!� � � 
� � � 
� � �$� � � 
� � � 
� � �'� � � 
� � � 
� � �*� � � 
� �n ,"�"^-�^ 
�V/�V 
�S 1"�"C2�C 
�94
�^  "D qR  "I q`  *Py^ *2t` *2t[ * |^ *:} |<"" |=*$B |>*4Z � "Z                                                                                                                                                                                                                         �� R @       �    @ 
        �     g P E g  ��         
            �������������������������������������� ���������	�
��������                                                                                          ��    �;�   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, 7  $ G�@,@����� ����                                                                                                                                                                                                                                                                                                                                      �� ��A���                                                                                                                                                                                                                                      >    -    � �  4�J     ��  	                           ������������������������������������������������������                                                                     	 	                                                                 �  ��^                        �^ (             	 
     �������� ��� ��������  ����� ��� �� ���������������������  ���  �� � � �� ������������ ��� ��� ���������������������������� ������ ����� ����������������� ��� ��������� ���� ������������ �� ���������������������� �           �             	    A  	  '     ��  L�J                                     �������������������������������������������������������                                                                                                                      	                  �    �c                         � �             	 	  ��������� ��������� �������������� �� ������� �������� ������������������ ����� ������ ������� � ���������������������������� ��� ��������� �� �������� ��� ��� ������������� ������� ����   ��� ���������������� ���� ����             (                                                                                                                                                                                                                                                                                                           �             


           �   }�    �                                                           R�  '�                     ������������       ����������������������������   &��������������������  'r����  'r���������������������ww�ww333wwwwwwww�ww�ww�ww�ww333wwww 4 H <                                 � Uei� �\                                                                                                                                                                                                                                                                                    �
  	��                                            m                                           ��                                                                                                                                                                                                                                                                                                                                                                 ( `  (`  @`  � 0��  � (��  EZm( ��d�� �N �����������������������������������                ���A :�� 9 
         �   & AG� �  �   
              �                                                                                                                                                                                                                                                                                                                                      p N I   �     p                 !��                                                                                                                                                                                                                            Y   �� �� ����      �� 8   	 
�������� ��� ��������  ����� ��� �� ���������������������  ���  �� � � �� ������������ ��� ��� ���������������������������� ������ ����� ����������������� ��� ��������� ���� ������������ �� ���������������������� � ��������� ��������� �������������� �� ������� �������� ������������������ ����� ������ ������� � ���������������������������� ��� ��������� �� �������� ��� ��� ������������� ������� ����   ��� ���������������� ���� ����              $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    8      5     ��                       8     �   �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p����      � �N     `d     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@       �      �     ��        # � ��� �� � ��� 1G� � �  �� �  �      �      3�������2����   g���   �     f ^�         ��M��      3      �������2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                          �      �  a r!   f�"""""*��**"*�"�""�""v""*f   "  ""- ��"�"*"-""z"""""����            n   �  "  q  ��                          �  �                                 � gv"!g�vg�vggfvv|�b��r""gb"�vr�rgb��v���g���v���***�*q!q�"!a�!vwfqqr~� qw��q�~~q�����~~~�w~~w�w            �   ~   ��  ~~  �w      v    �                ggj�vvggvvgg!vg�g֪vvg�r�r��⢪rq**gjb�v�q*gjj*vv��gg�z�/�"!�"�*�""*z����qw�~q~ww��q~qwvq�w�`� ��� �w �~p w�p  ��                    �                        lggz�v��g        �       ggbvvrgggavvvqggav� �      ���w!z�w"""�!""*�"! ��        q� q�        `               �        �                      wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                               s   D   O   w   w   v   u   f   T   �   �              3@  DDp ��4 ��tp��wpO�tpdfwGfeTwfeWwfUFwdUFweTfp�DDp���p���@�w�p   C   D   O   D   w   u   U   U  F  d  f   f   D   �   �   �DD ���7���uP��e`O�V ffg ffG Ufw UU� FUN dFw ffp DDp ��p ��@ w�p  C4 4D@O�C���O�Dt�GVfeVfdFfdFfdUfffUfffwFff�DDD���� ���                    0   G   W   W   U   E   E   w   �   �   @    fg D� O�� �� w�}�w��}����������M���M���M��������y�                    �   �   �   �   �   �   �   �   ~   w       ���w���w���~���~�DMw�������������y�                        w���w}��wt��wt��w}M�����������   M   M   ~�  p�  p   p   p      �   �   �   �               vd  eVp ffpw�Op���w���G���M�}�                                     v   ub  ub  f   `   P               "  f  U` wfP        p   p   p   p   p   p   p   p                               C4 �y�                              f  vU`vf`D�O������p}�w�  ?�  ?�  ?�  33  3#                                      f  Ug	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  " ! " ""                "                                                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  "!  "" "  """ !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  " ! " ""                "                                                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                       ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                      ��  ��  ���              �  �˰ ��� �wp ���                                                                                                                                                                  ˰ ̻ ̻ �� {�  �� 
�� ��� ��� ������
���	��ܻ̍ݻ���"� 8"  8  �  D�  H�  X�  ��  �   �          "  "     �                        ��  ��� �̺�̻����ۻ�˽��̽��̝ ̙� �30 �EP �U@ �T0 EC0 T3  C:  K�  �"  �"/ ����˽� �"� "" �""� � �� ��      �   �� ��  �"  �                   
 "� ""� ""� "                       �                             ���                         �  ��                    �����                       �       �                        �   ��  ���  � �    �                                                                                                                                                     � � ̹ �� �� �� ��� ��� �̻ 9�� EJ� EJ� 4D� 3DJ 4Z 3D �E ɽˠ
� "" �"�"! �"��" ��   �            �  �˰ ̻� ��p �wp ��  ��  ��  ��  ��  �̰ ۻ� ݙ� ݪ� =�� 0�  �   �   �   �   �   �   �   �   �   "   "�    ��  �    �      �   �" �"� "������     �     �� �� ��
��׊��w٪�|��������            "   "   "       �         �        �   �     �       �   �   �   �   �      �                    ��� ���� ��         �  ��� ݼ� w{� �װ vw�    �   ��  �   ��   �       �                                                                                                                                               � � ̹ �� �� �� ��� ��� �̻ 9�� EJ� EJ� 4D� 3DJ 4Z 3D �E ɽˠ
� "" �"�"! �"��" ��   �            �  �˰ ̻� ��p �wp ��  ��  ��  ��  ��  �̰ ۻ� ݙ� ݪ� =�� 0�  �   �   �   �   �   �   �   �   �   "   "�    ��  �    �          �  ��  �  ��  �            �  �   �   ��  �             ��  ��  �                            �   �    �   �       �   �   �                .          � ��                    ���� �                           �   ��  ���  � �    �                                                                                                                                       � ��~ ��� �}~ g~  ׮  
�  ��  �� ̾��� ��� ��� �� �� ��� �" "  �                           "   ¨�ˋ��˜��̌������ ��������˻�˻�����D���C��ET��EUZ�U ����Z� ��  �   �        "   "   "       �              �       33  DD3�DD;�3C��34��D� �U��� ��̰ �̰  ̊  ɫ  ��  ""  ""��"� �                                              �   �  �  �     �   �   �   �   �   �   �   �"" ""!! ��� �          �  �  ��  �   �   �         ���� �                                                                                                                                                                                              �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �           �   �     �   �               �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                                        	�  ���+��"+��-��  �  	�  X� U� EU 4U 4U  EU UU ̵Z��Uʜ��̨� ��  �"/ ""/�/���"���"�� ��           ˰ �� ̽ �����ך��pə���˙��̻���ݻ̽݉��ت��ۘ��ݰ��  U�  U�  Z�  �   �                       ��  ��� ��                     �   �   �                              �   �   ��   �    �     �                              "��" �"  �"     ��   �          ���� ��� ����               �  �  �  �                   ��   �  ��  �  �  �         � �������������  �       �  �   �   �   �                                                                                                                 �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   �   �"  ""  !� �� ��  �               �   ������  ��   "   "   "  �� ��                   ����������                          �  �� ��  �    � ���                                  � �������������  �                                                                                                                                       �UCD�UTE
EUT �T8 �D�  ��  �  �   �   �      �  �  �� �� ��EO  TO  C�� ��� ��� ������̻�̻�̻�w˙�b��v&���}��ۻ����ȯ����                       �ϻ��̋��̨���z������ ��  ��  ��  ��  �                           ��  "   "/  ./� "�� �   �   ��     �                    �   ��  �  �   ��  �  �  �� �� ��  �� �,� �"/�""�"/� "/  �         "  "  ""  "+� �� � ��   �  "   "�  +�  
�� ��� D�D 4ETO3    �   �   �   D   E�  U�  UO                         "  "  "                                                                                                                                                                      �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   ɪ  ��� ټ� �̰ �̰ ��� ��  ��                              ��                     �   �                      �������  ���    �                    ��  ��  ���                         ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                                            �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                               � ����ݼ� ����                                                                                                                                                                  �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �   �   �   ˰  ˙  ɪ  ��� ټ� �̰ �̰ ��� ��  ��                              ��  �   �   �                                      �������  ���    �                            � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                               �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��   �  �   
�  �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                             "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`����������������  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq:K �0K �,cj< cr$c� �J� �J� � �J� � �	B� � � 
B� � � � � � � � �k� � �k� � �k� � � k� � �	� � �	�  �� � �� �"� � � "� � �� � �
� �>"� �> "� �."� �.*� � �"� � � "� � �� � � 
� � �!� � � 
� � � 
� � �$� � � 
� � � 
� � �'� � � 
� � � 
� � �*� � � 
� �n ,"�"^-�^ 
�V/�V 
�S 1"�"C2�C 
�94
�^  "D qR  "I q`  *Py^ *2t` *2t[ * |^ *:} |<"" |=*$B |>*4Z � "Z3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3�������������������������������������������,�X�K�T�Z��<�[�Z�Z�K�X� � � � � � � � �-�2�3�����������������������������������������!��9�G�Z��6�G�0�U�T�Z�G�O�T�K� � � � � � �,�>�0�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�2�3� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�A�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                