GST@�                                                            \     �                                               T���      �               ���2�����	 J�������������������        �g     #    ����                                d8<n    �  ?     �����  �
fD�
�L���"����D"� j   " B   J  jF�"    
 �j� � 
 ���
��
�"     "�j��   * ��
   �                                                                              ����������������������������������      ��    =b 0Qb 4 114  4c  c  c        	 
      	   
       ��G �� � ( �(                 �nn 	)1         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                �   T       �   @  &   �   �                                                                                 '      	�)n1n  �    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE T �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    QtpTDs� �BA�@��|/�K�����#Cs�:	��K���c�-T0 k� �����e2$ 4r1'TP ��    ��� QtlTDs� �BA�@��|/�K�����$CC�9
�K���c�,T0 k� C�����e2$ 4r1'TP ��    ��� QtlTDs� �BA�@��|/�K�����$CC�8
�K��c�,T0 k� C�����e2$ 4r1'TP ��    ��� QtlTDs� �BA�@��|/�K�����%CC�7
�K��c�+T0 k� C�����e2$ 4r1'TP  ��    ��� QtlTDs� �BA�@��|/�K�����%CC�5
�K��c�*T0 k� C�����e2$ 4r1'TP  ��    ��� QtlTDs� �BA�@��|/�K�����&CC�4
�K��c�*T0 k� C�����e2$ 4r1'TP  ��    ��� QtlUDs� �BB @��|/�K�����&CC�2	��K��c�)T0 k� �����e2$ 4r1'TP  ��    ��� QthUDw� �BB@��|/�K����'CC�/	��K��c�(T0 k� �����e2$ 4r1'TP  ��    ��� QthUDw� �BB@��|/�K����(CC�.	��K��c�'T0 k� �����e2$ 4r1'TP  ��    ��� QthUDw� �BBA�|/�K����(CC�,	��K��c�'T0 k� �����e2$ 4r1'TP  ��    ��� QthUDw� �BBA�|/�K����(CC�*
�K��c�&T0 k� #�����e2$ 4r1'TP  ��    ��� QthUDw� �BBA�|/�K����)CC�)
�K��c�&T0 k� #�����e2$ 4r1'TP  ��    ��� QthVDw� �BBA�|/�K����)CS�'
�K��c�&T0 k� #�����e2$ 4r1'TP  ��    ��� QthVDw� �BB A�|/�K����*CS�%
�K��c�&T0 k� #�����e2$ 4r1'TP  ��    ��� QtdVDw� �BB$A�|/�K����*CS�#
�K��c�&T0 k� #�����e2$ 4r1'TP  ��    ��� QtdVDw� �BB(A�|/�K����+CS|!	��K��c�&T0 k� �����e2$ 4r1'TP  ��    ��� QtdVDw� �BB,A�|/�K����+CS|	��K��c�&T0 k� �����e2$ 4r1'TP  ��    ��� QtdVD{� �BB0A�|/�K����,CSx	��K��c�&T0 k� �����e2$ 4r1'TP  ��    ��� QtdVD{� �BB4A�|/�K����,CSx	��K��c�&T0 k� �����e2$ 4r1'TP  ��    ��� QtdWD{� �BB8A#�|/�K����,CSt	��K��c�&T0 k� �����e2$ 4r1'TP  ��    ��� QtdWD{� �BB8A#�|/�K����-CStD�K��c�&T0 k� �����e2$ 4r1'TP  ��    ��� QtdWD{� �BB<A'�|/�K����-CSpD�K��c�&T0 k� �����e2$ 4r1'TP  ��    ��� QtdWD{� �BB@A+�|/�K����-CSpD�K��c�&T0 k� �����e2$ 4r1'TP  ��    ��� Qt`WD{� �BBDA/�|/�K��� .CclD�K��c�&T0 k� �����e2$ 4r1'TP  ��    ��� Qt`WD{� �BBHA/�|/�K���.CclD�K��c�'T0 k� �����e2$ 4r1'TP  ��    ��� Qt`WD{� �BBLA3�|/�K���/Cch �K��c�'T0 k� �����e2$ 4r1'TP  ��    ��� Qt`WD{� �BBLA7�|/�K���/Cch
 �K��c�'T0 k� �����e2$ 4r1'TP  ��    ��� Qt`XD� �BBPA7�|/�Kӯ�/Ccd �K��c�'T0 k� �����e2$ 4r1'TP  ��    ��� Qt`XD� �BBTA;�|/�Kӯ�0Ccd �K��c�'T0 k� �����e2$ 4r1'TP  ��    ��� Q�`XD� �BBXA?�|/�Kӫ�0Cc` �K��c�'T0 k� �����e2$ 4r1'TP  ��    ��� Q�`XD� �BBXA?�|/�Kӫ�0Cc` �K��c�'T0 k� �����e2$ 4r1'TP  ��    ��� Q�`XD� �BB\AC�|/�Kӫ�0Cc_� �K��c�'T0 k� �����e2$ 4r1'TP  ��   ��� Q�\XD� �BB`AG�|/�Kӫ�� 0Cc_� �K��c�'T0 k� �����e2$ 4r1'TP  ��    ��� Q�\XD� �BBdAG�|/�E3���(1Cc[� d�K��c�(T0 k� �����e2$ 4r1'TP  ��    ��� Q�\XD� �BBdAK�|/�E3���,1Cs[� d�K��c�(T0 k� �����e2$ 4r1'TP  ��    ��� Q�\XD� �BBhAK�|/�E3���01CsW� d�K��c�(T0 k� �����e2$ 4r1'TP  ��    ��� Q�\YD� �BBlAO�|/�E3���41CsW� d�K��c�(T0 k� �����e2$ 4r1'TP  ��    ��� Q�\YD� �BBlAS�|/�E3���80CsW� d�Kӣ�c�(T0 k� �����e2$ 4r1'TP  ��    ��� U$\YD� �BBpAS�|/�Kӧ��<0CsS� d�Kӣ�c�(T0 k� �����e2$ 4r1'TP  ��    ��� U$\YD� �BBtAW�|/�Kӧ��@0E3S� d�Kӣ�c�(T0 k� �����e2$ 4r1'TP  ��    ��� U$\YD�� �BBtAW�|/�Kӣ��D0E3O� d�Kӣ�c�(T0 k� �����e2$ 4r1'TP  ��    ��� U$\YD�� �BBxA[�|/�Kӣ��H/E3O� d�Kӣ�c�(T0 k� �����e2$ 4r1'TP  ��    ��� U$\YD�� �BB|A[�|/�Kӣ��L/E3O� d�Kӟ�c�(T0 k� �����e2$ 4r1'TP  ��    ��� U$\YD�� �BB|A_�|/�Kӣ��P/E3O� d�@���c�(T0 k� �����e2$ 4r1'TP  ��    ��� U$XYD�� �BB�A_�|/�Kӣ��T.E#O� d�@���c�)T0 k� �����e2$ 4r1'TP  ��    ��� U$XYD�� �BB�Ac�|/�Kӣ��X.E#K� ��@���c�)T0 k� �����e2$ 4r1'TP  ��    ��� U$XYD�� �BB�Ac�|/�Kӣ��\-E#K� ��@���c�)T0 k� �����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�Ag�|/�Kӟ��`,E#K� ��@���c�)T0 k� ����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�Ag�|/�Kӟ��d,E#K� ��Kӟ�c�)T0 k� �����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�Ak�|/�K㟺�d+B�K� ��Kӟ�c�)T0 k� �����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�Ak�|/�K㟹�h*B�O� ��Kӛ�c�)T0 k� �����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�Ao�|/�K㟹�l)B�O� ��Kӛ�c�)T0 k� �����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�Ao�|/�K㟸�p)B�O� ��Kӛ�c�)T0 k� �����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�As�|/�K㟸�t(B�O� ��Kӛ�c�)T0 k� �����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�As�|/�K㛷Sx'E#O� ��Kӛ�c�)T0 k� �����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�Aw�|/�K㛷Sx&E#S� ��Kӛ�c�)T0 k� �����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�Aw�|/�K㛶S|%E#S� ��Kӛ�c�)T0 k� �����e2$ 4r1'TP  ��    ��� @dXZD�� �BB�Aw�|/�K㛶S|%E#S��Kӛ�c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dTZD�� �BB�A{�|/�K㛵S|%E#W��Kӛ�c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[D�� �BB�A{�|/�K㛵S�%E#W��Kӗ�c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[D�� �BB�A�|/�K㛴S�$EW��Kӗ�c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[D� �BB�A�|/�K㛴S�$E[��Kӗ�c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[D� �BB�A�|/�K㛴S�#E[��K��c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[D� �BB�A��!�/�K㟴S�#E[��K��c�*T0 k� �����e2$ 4r1'TP  ��   ��� @dT[D� �BB�A��!�/�K㟳S�#E[��K��c�*T0 k� �����e2$ 4r1'TP  ��   ��� @dT[D{� �BB�A��!�/�K㣳S�"B�[���K��c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[D{� �BB�A��!�/�K㣲S�"B�[���K��c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[D{� �BB�A��!�/�K㣱c�"B�[���K��c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[D{� �BB�A��!�/�K㧱c�"B�_���K��c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[D{� �BB�A��!�/�K㧰c�"B�_���K��c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[Dw� �BB�A��!�/�K㧰c�"B�c���K��c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[Dw� �BB�A��!�/�K㫯c�"K�c���K��c�*T0 k� �����e2$ 4r1'TP  ��    ��� @dT[Dw� �BB�A��!�/�K㫯c�!K�c���K��c�+T0 k� �����e2$ 4r1'TP  ��    ��� @dT[Dw� �BB�A��!�/�K㫮c�!K�g���K��c�+T0 k� �����e2$ 4r1'TP  ��    ��� @dT\Dw� �BB�A��|/�K㯮c�!K�g���K��c�+T0 k� �����e2$ 4r1'TP  ��    ��� @dT\Ds� �BB�A��|/�K㯭c�!K�k���K��c�+T0 k� �����e2$ 4r1'TP  ��    ��� @dT\Ds� �BB�A��|/�K㯭c� K�k���K��c�+T0 k� �����e2$ 4r1'TP  ��    ��� @dT\Ds� �BB�A��|/�K㳬c� K�k���K��c�+T0 k� �����e2$ 4r1'TP  ��    ��� @dP\Ds� �BB�A��|/�K㳬c� K�o���K��c�+T0 k� �����e2$ 4r1'TP  ��    ��� @dP\Ds� �BB�A��|/�K㳫c� K�o��K��c�,T0 k� �����e2$ 4r1'TP  ��    ��� @dP\Do� �BB�A��|/�K㷫c� K�s��K��c�,T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Do� �BB�A��|/�K㷪c� K�s��K��c�,T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Do� �BB�A��|/�K㷪c�K�s��K��c�,T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Do� �BB�A��|/�K㻩c�K�w��K��c�,T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Do� �BB�A��|/�K㻩c�K�w��K��c�,T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Do� �BB�A��!�/�K㻨c�K�w��K��c�-T0 k� ����e2$ 4r1'TP  ��   ��� @dP\Dk� �BB�A��!�/�K㻨c�K�{��K��c�-T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Dk� �BB�A��!�/�K㿧c�K�{��K��c�-T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Dk� �BB�A��!�/�K㿧c�K�{��K��c�-T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Dk� �BB�A��!�/�K㿧c�K���K㏿c�-T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Dk� �BB�A��!�/�Kӿ�c�K���K㏿c�-T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Dk� �BB�A��!�/�K�æc�K���K㏿c�-T0 k� ����e2$ 4r1'TP  ��    ��� @dP\Dk� �BB�A��!�/�K�åc�K����K㏿c�.T0 k� ����e2$ 4r1'TP  ��    ��� @dP]Dg� �BB�A��!�/�K�åc�K����K㏾c�.T0 k� ����e2$ 4r1'TP  ��    ��� @dP]Dg� �BB�A��!�/�K�åc�K����K㏾c�.T0 k� ����e2$ 4r1'TP  ��    ��� @dP]Dg� �BB�A��!�/�K�Ǥc�K����K㏾c�.T0 k� ����e2$ 4r1'TP  ��    ��� @dP]Dg� �BB�A��|/�E#Ǥc�K����K㏾c�.T0 k� ����e2$ 4r1'TP  ��    ��� @dP]Dg� � BB�A��|/�E#ǣc�K����K㏾c�.T0 k� ����e2$ 4r1'TP  ��    ��� @dP]Dg� � BB�A��|/�E#ˣc�K����K㏽c�/T0 k� ����e2$ 4r1'TP  ��    ��� @dP]Dg� � BB�A��|/�E#ˢc�K����K㋽c�/T0 k� ����e2$ 4r1'TP  ��    ��� @dP]Dc� �!BB�A��|/�E#ϡc�K����K㋽c�/T0 k� ����e2$ 4r1'TP  ��    ��� @dP]Dc� �!BB�A��|/�E#ϡc�K����K㋼c�/T0 k� �����e2$ 4r1'TP  ��    ��� @dP]Dc� �!BB�A��|/�E#Ӡc�K����KӋ�c�/T0 k� �����e2$ 4r1'TP  ��    ��� @dP]Dc� �!BB�A��|/�E#Ӡc�K����KӋ�c�/T0 k� �����e2$ 4r1'TP  ��    ��� @dP]Dc� �!BB�A��|/�E#ןc�K����KӋ�c�0T0 k� �����e2$ 4r1'TP  ��    ��� @dP]Dc� �!BB�A��|/�E#מc�K����KӋ�c�0T0 k� �����e2$ 4r1'TP  ��    ��� @dP]Dc� �!BB�A��|/�E#۞c�K����KӋ�c�0T0 k� �����e2$ 4r1'TP  ��    ��� @dP]Dc� �!BB�A��|/�E۝S�K����KӋ�c�0T0 k� �����e2$ 4r1'TP  ��    ��� @dL]D_� �!BB�A��|/�EߜS�K����@���c�0T0 k� �����e2$ 4r1'TP  ��    ��� @dL]D_� �"BB�A��|/�EߜS�K����@���c�0T0 k� �����e2$ 4r1'TP  ��    ��� @dL]D_� �"BB�A��|/�E�S�K����@���c�1T0 k� �����e2$ 4r1'TP  ��    ��� @dL]D_� �"BB�A��|/�E�S�K����@���c�1T0 k� �����e2$ 4r1'TP  ��    ��� @dL]D_� �"BB�A��|/�E�S�K����@���c�1T0 k� �����e2$ 4r1'TP  ��    ��� @dL]D_� �"BB�A��|/�E���K����@���c�1T0 k� �����e2$ 4r1'TP  ��    ��� @dL]D_� �#BB�A��|/�E����K����@���c�1T0 k� �����e2$ 4r1'TP  ��    ��� @dL]D_� �#BB�A��|/�E����K����@���c�1T0 k� �����e2$ 4r1'TP  ��    ��� @dL]D_� �#BB�A��|/�E����K����@���c�1T0 k� �����e2$ 4r1'TP  ��    ��� @dL^D_� �#BB�A��|/�E����K����@���c�1T0 k� �����e2$ 4r1'TP  ��    ��� @dL^D[� �#BB�A��|/�E�����K����@���c�2T0 k� �����e2$ 4r1'TP  ��    ��� @dL^D[� �$BB�A��|/�E�����K�����@���c�2T0 k� �����e2$ 4r1'TP  ��    ��� @dL^D[� �$BB�A��|/�E�����K�����@���c�2T0 k� �����e2$ 4r1'TP  ��    ��� @dL^D[� �$BB�A��|/�Et���K�����@���c�2T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^D[� �$BB�A��|/�Et���K�����@���c�2T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^D[� �$BB�A��|/�Et���K�����@���c�2T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^D[� �$BB�A��|/�Et���K�����@���c�2T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^D[� �%BB�A��|/�Et���K�����@���c�2T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^D[� �%BB�A��|/�Et���K����@���c�3T0 k� �w��{�e2$ 4r1'TP  ��    ��� @dL^D[� �%BB�A��|/�Et���K����KӇ�c�3T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^D[� �%BB�A��|/�Et���K����KӇ�c�3T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^D[� �%BB�A��|/�Et���K����KӇ�c�3T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �%BB�A��|/�Ed���K����KӇ�c�3T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �%BB�A��|/�Ed���B���T�KӇ�c�3T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �&BB�A��|/�Ed#���B���T�KӇ�c�3T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �&BB�A��|/�Ed#���B���T�KӇ�c�3T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �&BB�A��|/�Ed'���B���T�KӇ�c�3T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �&BB�A��|/�D4'���B���T�KӇ�c�4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �&BB�A��|/�D4'���
E��T�KӇ�c�4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �&BB�A��|/�D4'���	E��T�KӇ�c�4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �&BB�A��|/�D4+���E��T�KӇ�c�4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �'BB�A��|/�D4+���E��T�KӇ�c�4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �'BB�A��|/�D4+���E���KӇ�c�4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �'BB�A��|/�D4/���E����Kㇷc�4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �'BB�A��|/�D4/���E�É�Kㇷc�4T0 k� �{���e2$ 4r1'TP  ��   ��� @dL^DW� �'BB�A��|/�D4/���E�Ǌ�Kㇷc�4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DW� �'BB�A��|/�D4/����E�ˊ�Kㇶc�4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DS� �'BB�A��|/�D43����E�ϊ�Kㇶc�4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DS� �'BB�A��|/�D43����D�Ӌ�Kㇶc�5T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DS� �(BB�A��|/�DD3����D�׋�Kㇶ��5T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DS� �(BB�A��|/�DD3����D�ی�Kㇶ��4T0 k� �{���e2$ 4r1'TP  ��    ��� @dL^DS� �(BB�A��|/�DD3����D�ߍ�Kㇶ��4T0 k� �{���e2$ 4r1'TP  ��   ��� E���T7���#C�,��|#�G�P(��LDC��⇂EC<I3�T0 k� �<�<e2$ 4r1'TP  ��/    � &��E���T3���#C�(��|#�G�P)��LDC���EC8I3�T0 k� ��<� <e2$ 4r1'TP  ��/    � &��D3��T/���#C� ��|#�G�L)��LDC{��w�EC4I3�T0 k� ��=��=e2$ 4r1'TP  ��/    � &��D3��T+���#C���|#�C�H)��LDCw��o�EC4H3�T0 k� ��>��>e2$ 4r1'TP  ��/    � &��D3���'�a�"C���|#�C�D)иLDSs��g�E30H3�T0 k� ��?��?e2$ 4r1'TP  ��/    � &��D3���#�a�"C���|#�C�@)�KDSo��_�E3,G3�T0 k� ��@��@e2$ 4r1'TP  ��/    � &��D3����a�"C���|#�C�<)�KDSk��W�E3,G3�T0 k� �A��Ae2$ 4r1'TP  ��/    � &��D3����a�"C���|#�C�8*�KDSg��O�E3(F3�T0 k� �B��Be2$ 4r1'TP  ��/    � &��D3����a�!C� ��|#�C�4*�KDSc��G�E3$E3�T0 k� �C��Ce2$ 4r1'TP  $�/    � &��D3����a�!C�� ��|#�C�0*��JES_��?�E#$E3�T0 k�  �B��Be2$ 4r1'TP  ��/    � &��D3����a� C�����|#�C�,*0�JESW��7�E# D3�T0 k�  �@��@e2$ 4r1'TP  ��/    � &��D3����a| C�����|#�C�(*0�JESS��/�E# C3�T0 k�  �?��?e2$ 4r1'TP  ��/    � &��D3�����QxC�����|#�C�$*0�IESO��'�E#C3�T0 k�  �=��=e2$ 4r1'TP  ��/    � &��D3�����QpC�����|#�C� *0xIESG���E#B3�T0 k�  �<��<e2$ 4r1'TP  ��/    � &��DC����QhC�����|#�C�*0tHESC���EA3�T0 k� �;��;e2$ 4r1'TP  ��/    � &��DC����QdC����|#�C�*0lHES?���E@3�T0 k� �9��9e2$ 4r1'TP  ��/    � &��DC����Q\D��w�|#�C�*0dGC�7���E@3�T0 k� �8��8e2$ 4r1'TP  ��/    � &��DC{����TD��o�|#�C�*0\GC�/����E?3�T0 k� �6��6e2$ 4r1'TP  ��/    � &��DCs��۸�PD��Qg�|#�C�*0TFC�'���E>3�T0 k� �5��5e2$ 4r1'TP  ��/    � &��DCk��׸�HD��Q_�|#�C�*0LEC����E=3�T0 k� �4��4e2$ 4r1'TP  ��/    � &��DCg��Ϸ�@D��QW�|#�C�*@DEC����E=3�T0 k� �2��2e2$ 4r1'TP  ��/    � &��DC_��Ƕ�8D��QO�|#�C�*@<DC���ۄE<3�T0 k� �1��1e2$ 4r1'TP  ��/    � &��DCW���0D��QG�|#�C�*@4CC��υE;3�T0 k� ��0��0e2$ 4r1'TP  ��/    � &��DCO���(D��AC�|#�C�*@,BC���ǅE;3�T0 k� ��.��.e2$ 4r1'TP  ��/    � &��DCG����D��A;�|#�C�*@$BC�����E�:3�T0 k� ��-��-e2$ 4r1'TP  ��/    � &��DS?����D��A3�|#�C�*@AC�����E�:3�T0 k� ��+��+e2$ 4r1'TP  ��/    � &��DS7���� D��A+�|#�D*@@C�����E�93�T0 k� ��*��*e2$ 4r1'TP  ��/    � &��DS3�����D��A#�|#�D*@?C�����E� 93�T0 k� ��)��)e2$ 4r1'TP  ��/    � &��DS+�����D{�A�|#�D*@>C�����E� 83�T0 k� ��'��'e2$ 4r1'TP  ��/    � &��DS#�����Ds�1�|#�D*O�=C�����E� 83�T0 k� ��&��&e2$ 4r1'TP  ��/    � &��ES�����Dk�1�|#�D*O�<C�����E�$83�T0 k� ��%��%e2$ 4r1'TP  ��/    � &��ES�{���Dc�1�|#�D*_�;C���E�$73�T0 k� �� �� e2$ 4r1'TP  ��"    � &��ES�s�дD[�0��|#�D*_�:C��w�E�(73�T0 k� �t�xe2$ 4r1'TP  ��"    � &��ER��k�ШDS�0��|#�J�*_�:C��o�E�(73�T0 k� �h�le2$ 4r1'TP  ��"    � &��ER��c�МDK�0��|#�J�*_�9E��g�D�,73�T0 k� �\�`e2$ 4r1'TP  ��"    � &��ER��[�АDC�0��|#�J�*_�8E��_�D�073�T0 k� �P�Te2$ 4r1'TP  ��"    � &��ER��S�ЄD;�0��|#�J�*_�7E��S�D�073�T0 k� �D�He2$ 4r1'TP  ��"    � &��ER��K��xD3�0��|#�J�*_�6E��K�D�473�T0 k� �8�<e2$ 4r1'TP  ��"    � &��E���C��lC�'����|#�J�*_�5E��QC�D�873�T0 k� �0�4e2$ 4r1'TP  ��"    � &��E���;��`C�����|#�J�*_�4E�s�Q;�D�873�T0 k� �$�(e2$ 4r1'TP  ��"    � &��E���3��XC�����|#�J�*_�3E�k�Q3�D�<73�T0 k� ��e2$ 4r1'TP  ��"    � &��E��+��LC�����|#�J�*_�2E�c�Q'�D�@73�T0 k� ��e2$ 4r1'TP  ��"    � &��E��#��@C�����|#�J�*_�1E�[�Q�D�D73�T0 k� ��e2$ 4r1'TP  ��"    � &��E����8C������|#�J�*_�0E�O�A�D�D73�T0 k� ����e2$ 4r1'TP  ��"    � &��E����,C������|#�J�*_�/D2G�A�D�H73�T0 k� ����e2$ 4r1'TP  ��"    � &��E����$C������|#�J�*_�.D2?�A�D�L73�T0 k� ����e2$ 4r1'TP  ��"    � &��E������C������|'�J�*_x-D27�@��D�L73�T0 k� ����e2$ 4r1'TP  ��"    � &��E������C������|'�J�*_p,D2/�@�D�P73�T0 k� ����e2$ 4r1'TP  ��"    � &��D2�����C������|'�J�*_h+D2'���D�P73�T0 k� ����e2$ 4r1'TP  ��"    � &��D2{�����C���Ѓ�|'�J� *_`+D2���D�T73�T0 k� ����e2$ 4r1'TP  ��"    � &��D2s��ߤo�C����{�|'�Eb *_X*D2��׊D�T73�T0 k� ����e2$ 4r1'TP  ��"    � &��D2k��ףo�C���s�|'�Eb$*_P)D2��ϊD�T73�T0 k� ����e2$ 4r1'TP  ��"    � &��D2c��ˣo�C���k�|'�Eb(*OH(D2��ǊD�X73�T0 k� ����e2$ 4r1'TP  ��"    � &��ER[��âo�C���g�|'�Eb()O@(D1��п�D�X73�T0 k� ����e2$ 4r1'TP  ��"    � &��ERS�⻢o�C���_�|'�Eb,)O8'D1��з�D�X73�T0 k� ����e2$ 4r1'TP  ��"    � &��ERK�ⳡ	��C���W�|'�Eb0)O0&D1��Ы�D�X73�T0 k� ����e2$ 4r1'TP  ��"    � &��ERC�⫡	��C����O�|'�K4)O(&DA��࣋D�X73�T0 k� ����e2$ 4r1'TP  ��"    � &��ER7�⣠	��C����G�|'�K8(O%DA�����D�X73�T0 k� ����e2$ 4r1'TP  ��"    � &��ER/��	��C�{��C�|'�K8(O%DA�����D�X73�T0 k� �|��e2$ 4r1'TP  ��"    � &��ER'��	��C�s��;�|'�K<(�$DA�����D�X73�T0 k� �x�|e2$ 4r1'TP  ��"    � &��C���	��C�k��3�|'�K@'�$DA����D�X73�T0 k� �t�xe2$ 4r1'TP  ��"    � &��C����	��D c��+�|'�KD'��$E���w�D�X73�T0 k� �p�te2$ 4r1'TP  ��"    � &��C���w�	��D W��#�|'�KH&��#E���o�BCX73�T0 k� �l�pe2$ 4r1'TP  ��"    � &��C���o�	��D O���|'�KL&��#E���g�BCX73�T0 k� �d�he2$ 4r1'TP  ��"    � &��C����g�	��D G���|'�KP%��#E���[�BCX73�T0 k� �`�de2$ 4r1'TP  ��"    � &��E����_�	��D G���|'�KT%��"E���S�BCX73�T0 k� �X�\e2$ 4r1'TP  ��"    � &��E����W�	�|D ?���|'�KX$��"E���K�BCX73�T0 k� �T�Xe2$ 4r1'TP  ��"    � &��E����K�	�xD 7����|'�KX$��"E���C�A�X73�T0 k� �P�Te2$ 4r1'TP  ��"    � &��E����C�	�tD /����|'�K\#��!E�{��7�A�X73�T0 k� �H�Le2$ 4r1'TP  ��"    � &��E�� ;�	�pD '����|'�K`"޸!E�s��/�A�X73�T0 k� �D�He2$ 4r1'TP  ��"    � &��E��3�	�lD ����|'�Kh"ެ!E�k��'�A�X73�T0 k� �@�De2$ 4r1'TP  ��"    � &��E��+�	�hD ����|'�Kl!ޤ E�g���A�X73�T0 k� �L�Pe2$ 4r1'TP  �"    � &��D1�#�	�`E�����|'�Kp!� E�_���A�X73�T0 k� �\�`e2$ 4r1'TP ��/    � &��D1��	�\E�����|'�E�t � E�W�@�A�X73�T0 k� �h�le2$ 4r1'TP ��/    � &��D1��	�XE������|'�E�x �E�O�@�A�X73�T0 k� �t�xe2$ 4r1'TP ��/    � &��D1���TE���߻�|'�E�|�E�G�O��A�X73�T0 k� ����e2$ 4r1'TP ��/    � &��D1����PE���߳�|'�EҀ�|E�?�O�A�X73�T0 k� ����e2$ 4r1'TP ��/    � &��D1�	���LE�����|'�E҈�pE�8O�A�X73�T0 k� ����e2$ 4r1'TP ��/    � &��D1�
��HE�����|'�EҌ�hE�0OߐA�X73�T0 k� ����e2$ 4r1'TP ��/    � &��D1���DE�����|+�EҐ�`E�(OבA�X73�T0 k� ����e2$ 4r1'TP ��/    � & D1xۘ�@E�����|+�JҔ�XF$�ϑA�X73�T0 k� ����e2$ 4r1'TP ��/    � & 	D1pӗ�<E�����|+�JҜ�PF�ǑA�X73�T0 k� ����e2$ 4r1'TP ��/    � & D1d˗�<K��o��|+�JҠ�HF	���A�X73�T0 k� ����e2$ 4r1'TP ��/    � & D1\×�8K��o�|+�JҤ�@F���A�X73�T0 k� ����e2$ 4r1'TP ��/    � & DALQ���0K��os�|+�ER��0FO��A�X73�T0 k� �"�"e2$ 4r1'TP ��/    � & !DADQ���,K��ok�|/�ER��(F O��A�X73�T0 k� �$�$e2$ 4r1'TP ��/    � & &DADQ���(E��oc�|/�ER�� F �O��A�X73�T0 k� �$%�(%e2$ 4r1'TP ��/    � & +DA@Q���$E��o_�|/�ER��F �O��ASX73�T0 k� �0'�4'e2$ 4r1'TP  ��/    � & 0DA8Q��� E��W�|/�ER��F �O��ASX73�T0 k� �@(�D(e2$ 4r1'TP  ��/    � & 5DA4Q��� E��S�|/�ER��F �Ow�ASX73�T0 k� �L*�P*e2$ 4r1'TP  ��/    � & :DA,Q��E��K�|/�EB�� F �Oo�ASX73�T0 k� �X+�\+e2$ 4r1'TP  ��/    � & ?DA(Aw��E��G�|/�EB���E��Og�ASX73�T0 k� �h-�l-e2$ 4r1'TP  /�/    � & DDA$Ak��E��C�|/�EB���E��?_�C�T73�T0 k� �t.�x.e2$ 4r1'TP  ��/    � & IDAAc��E��;�|/�EB��E��?W�C�T73�T0 k� ��0��0e2$ 4r1'TP  ��/    � & NDQA[��E��7�|/�EB��E��!?O�C�T73�T0 k� �1��1e2$ 4r1'TP  ��/    � & RDQAS��E�{�/�|/�E���E��"?G�C�P73�T0 k� �3��3e2$ 4r1'TP  ��/    � & VDQAK��E�s�+�|/�E���E��$??�C�P73�T0 k� �4��4e2$ 4r1'TP  ��/    � & ZDQA?��E�o�'�|/�E���E��&?7�C�L73�T0 k� �6��6e2$ 4r1'TP  ��/    � & ^DQ A7��E�g���|/�E���E��'?/�C�L73�T0 k� ��7��7e2$ 4r1'TP  ��/    � & \E�!A/�� E�c���|/�E���
E��)?'�C�H73�T0 k� ��8��8e2$ 4r1'TP  ��     � & ZE�!A���E�W���|/�E��M�E��-?�C�D73�T0 k� ��9��9e2$ 4r1'TP  ��  	   � & YE� "A���E�O���|/�E��M�E��.?�C�@73�T0 k� ��:��:e2$ 4r1'TP  ��  	   � & XE��#A���E�G���|/�C��M�E��0/�C�<73�T0 k� ��:��:e2$ 4r1'TP  ��  	   � & WE��%1���E�C����|/�C��M�E��1/�C�873�T0 k� ��;��;e2$ 4r1'TP  ��  	   � & VE��&0����E�;����|/�C��M�E��2.��C�473�T0 k� ��<��<e2$ 4r1'TP  ��  	   � & UE��(0���E3����|/�C��M�E��4.��C�073�T0 k� ��=��=e2$ 4r1'TP  ��  	   � & UE��)0���E+����|/�C��M� E��5.�C�,73�T0 k� ��?��?e2$ 4r1'TP  ��  	   � & UE��+0���E'����|/�C����E �6.�C�(73�T0 k� ��@��@e2$ 4r1'TP  ��  	   � & TE��+0ӗ��E��� |/�C����E �9.�C� 73�T0 k� ��C��Ce2$ 4r1'TP  ��  	   � & TE��,0˗��E��|/�C����E �:.۬D73�T0 k� ��C��Ce2$ 4r1'TP  ��  	   � & TE��.0Ø��E��|/�C����E �;.׮D73�T0 k� ��D��De2$ 4r1'TP  ��  	   � & TE��/0����E���|/�C�����E�=.ӯD73�T0 k� ��E��Ee2$ 4r1'TP  ��  	   � & TE��10����E���|/�C�����E�>.ϰD73�T0 k� ��G��Ge2$ 4r1'TP  ��     � & TE��3 ����E���|/�C�����E�?˲D73�T0 k� ��H��He2$ 4r1'TP  ��     � & TE��4 ����E���|/�C��
���E�@ǳD73�T0 k� ��J��Je2$ 4r1'TP  ��     � & TE��6 ����E���|/�C��
���E�AôD 73�T0 k� ��L��Le2$ 4r1'TP  ��     � & TF �8 ����E.��
�|/�C��
��B��B��D�73�T0 k� ��L��Le2$ 4r1'TP  ��     � & TF �; ����E.��
�|/�C��	��B��D��D�73�T0 k� ��M��Me2$ 4r1'TP  ��     � & TF �= ����E.��
�	!�/�C���{�B��E��D�73�T0 k� ��N��Ne2$ 4r1'TP  ��     � & TF �= ����E.��
�
!�/�C���{�B��F���D�73�T0 k� ��N��Ne2$ 4r1'TP  ��     � & UF �> ���JN��
�
!�/�C���{�B��G���D�73�T0 k� ��N��Ne2$ 4r1'TP  ��     � & VF �@ {���JN��
|!�/�C��{�B��H���D�73�T0 k� ��O��Oe2$ 4r1'TP  ��     � & WF �B w���JN��
t!�/�C��{�B��J���D�7"s�T0 k� ��P� Pe2$ 4r1'TP  ��     � & XF �C s���JN��
l!�/�D��{�E�K���D�7"s�T0 k� � Q�Qe2$ 4r1'TP  ��     � & YF �Eo���JN��
d!�/�D��{�E�L���D�7"s�T0 k� � R�Re2$ 4r1'TP  ��     � & ZF �Gk���JN��
\!�/�D��{�E�M���D�7"s�T0 k� � T�Te2$ 4r1'TP  ��     � & [E��Ig���JN{�
T!�/�D��{�E�N���D�7"s�T0 k� ��R� Re2$ 4r1'TP  ��     � & \E��Jc�N�JNs�
.L!�/�D��{�E�O���D�7"s�T0 k� ��Q� Qe2$ 4r1'TP  ��     � & ]E��Lc�N�JNk�
.H!�/�D��{�E�P���D�7"s�T0 k� ��P��Pe2$ 4r1'TP  ��     � & ^E��N_�N�JNc�
.@|/�D���E�Q���D�7"s�T0 k� ��P��Pe2$ 4r1'TP  ��     � & _E��O[�N�JN[�
.8|/�D���E�R���I��7"s�T0 k� ��Q��Qe2$ 4r1'TP  ��     � ' `E��Q[�N�J^O�
.0|/�D����E�S���I��7"s�T0 k� ��Q� Qe2$ 4r1'TP  ��     � ( aE��RW���J^G�
.(|/�D����E�S���I��7"s�T0 k� � R�Re2$ 4r1'TP  ��     � ) bE��T�W���J^?�
. |/�D����E��T���I��73�T0 k� � S�Se2$ 4r1'TP  ��     � * cE��U�W���J^7�
.|/�D����E��U���I�|73�T0 k� �T�Te2$ 4r1'TP  ��     � + dE��W�S���J^/�
.|/�D����E��V���I�t73�T0 k� �U�Ue2$ 4r1'TP  ��     � , eE��X�S���J^'�
.|/�D����E��W���I�p73�T0 k� �W�We2$ 4r1'TP  ��     � - fE��Z�S���J^�
.|/�D����E��X���I�h73�T0 k� �T�Te2$ 4r1'TP  ��     � . gE��[�S���J^�
�|/�Dx���E��Y���I�d73�T0 k� �S�Se2$ 4r1'TP  ��     � / hE��\�S���J^�
�|/�I�t���E��Z���I�`73�	T0 k� �R�Re2$ 4r1'TP  ��     � 0 iE� ^�S���J^�
�!�/�I�p���E��Z���I�\73�	T0 k� �R� Re2$ 4r1'TP  ��     � 1 jE�_�S���J]��
�!�/�I�l���E��[���I�X73�	T0 k� � R�$Re2$ 4r1'TP  ��     � 2 l@qa�S���JM��
�!�/�I�h���E��\ο�I�P73�	T0 k� �(Q�,Qe2$ 4r1'TP  ��     � 3 n@qb�S�� JM��
�!�/�I�d���E��]ο�I�L7"��	T0 k� �0P�4Pe2$ 4r1'TP  ��     � 4 p@qc�S��JM��
�!�/�I�`���B��]���I�H7"��	T0 k� �4O�8Oe2$ 4r1'TP  ��     � 5 r@qd�S��JM��
�!�/�I�\���B��^���I�D7"��	T0 k� �8O�<Oe2$ 4r1'TP  ��     � 6 t@q d�S��JM��
�!�/�I�X���B��^���I�@7"��	T0 k� �<O�@Oe2$ 4r1'TP  ��     � 7 v@q$e�W��JM��
�!�/�I�X���B��_���I�<7"��	T0 k� �DO�HOe2$ 4r1'TP  ��     � 8 x@q,f�W��JM��
=�!�/�I�T���B��_���I�87"��	T0 k� �HO�LOe2$ 4r1'TP  ��     � 9 z@q0f�W��JM��
=�!�/�I�T���B��_���I�87"S�	T0 k� �LO�POe2$ 4r1'TP  ��     � : |@q4g�[��JM��
=�|/�I�P��E�_���I�47"S�	T0 k� �TO�XOe2$ 4r1'TP  ��     � ; ~@q<g�[�� JM��
=�|/�I�P��E�_���I�07"S�	T0 k� �XP�\Pe2$ 4r1'TP  ��     � < �@q@h�[��$Jm��
=� |/�I�L��E `���I�07"S�	T0 k� �`P�dPe2$ 4r1'TP  ��     � < �@qHh�_��(Jm��
=� |/�I�L��E`���I�,7"S�	T0 k� �dQ�hQe2$ 4r1'TP  ��     � < �@�Lh�_��,Jm��
=�!|/�I�H��E`���I�,7�	T0 k� �hR�lRe2$ 4r1'TP  ��     � < �@�Ti�c��4Jm��
=�!|/�I�H��E`���I�(7�	T0 k� �pS�tSe2$ 4r1'TP  ��     � < �@�Xi�g��8Jm��
=�"|/�I�H��Ea���I�(7�	T0 k� �xT�|Te2$ 4r1'TP  ��     � < �@�`i�g��<Jm��
=�"|/�I�H��E a���I�(7�	T0 k� �|T��Te2$ 4r1'TP  ��     � < �@�di�k��DE���|#|/�I�D��E(a���I�$7�	T0 k� �T��Te2$ 4r1'TP  ��     � < �@�li�o��HE���x#|/�I�D��E0a��I�$7�
T0 k� �T��Te2$ 4r1'TP  ��     � < �@�ti�o��LE���t#|/�I�D��E�4a��I�$7�
T0 k� �T��Te2$ 4r1'TP  ��     � < �@�xi�s��TE���p$|/�I�D��E�<b��I�$7�
T0 k� �T��Te2$ 4r1'TP  ��     � < �@��i�w��`E���h%|/�I�D���E�<b��I�$7�
T0 k� �T��Te2$ 4r1'TP  �     � < �@��i�{��hE���d%|/�I�D���E�Dc��I�$7�
T0 k� �T��Te2$ 4r1'TP  ��     � < �@��i���lE���`&|/�I�D���PLd�#�I�$7�
T0 k� �T��Te2$ 4r1'TP  ��     � < �@��i����tE���`&|/�I�D���PTd�+�I�$7�
T0 k� ��T��Te2$ 4r1'TP  ��  	   � < �@��i����|E���\&|/�I�D���P\e�3�I�$7�
T0 k� ��T��Te2$ 4r1'TP  ��  	   � < �@��i���߄B����\'|/�I�D���Pdf�7�I�$7�T0 k� ��T��Te2$ 4r1'TP  ��  	   � < �@��i���߈B����X'|/�A�D���Plf�?�I�$7�T0 k� ��S��Se2$ 4r1'TP  ��  	   � < �@��h���ߐB����X(|/�A�D���Ptg�C�A�$7�T0 k� ��S��Se2$ 4r1'TP  ��  	   � < �@��h���ߘB����T(|/�A�D���Pxg�K�A�$7�T0 k� ��S��Se2$ 4r1'TP  ��  	   � < �@��h���ߠB����T(|/�A�D��P�h�S�A�$7�T0 k� ��S� Se2$ 4r1'TP  ��  	   � < �@��h���ߨB����T)|/�A�D��P�i�[�A�$7�T0 k� �R�Re2$ 4r1'TP  ��  	   � < �@��g���߰B����T)|/�A�D��P�i�_�A�$7�T0 k� �R�Re2$ 4r1'TP  ��  	   � < �@��g�����B����T)|/�A�D��P�j�g�BB$7�T0 k� �R�Re2$ 4r1'TP  ��  	   � < �@��g�����B����T*|/�A�D��P�j�o�BB$7�T0 k� �S�Se2$ 4r1'TP  ��  	   � < �@�f�����B����T*|/�A�D�#�P�k�w�BB$7�T0 k� � T�$Te2$ 4r1'TP  ��  	   � < �@�f�����B����T*|/�A�D�+�P�k��BB$7�T0 k� �$T�(Te2$ 4r1'TP  ��  	   � < �@�e�����B����T+|/�D�D�/�P�l���BB$7�T0 k� �(T�,Te2$ 4r1'TP  ��  	   � < �@�$e�Ǩ��B����T+|/�D�D�7�P�l���@$7�T0 k� �4T�8Te2$ 4r1'TP  ��  	   � < �@�,d�˧��B����T+|/�D�H�?�P�m���@$7�T0 k� �<T�@Te2$ 4r1'TP  ��  	   � < �@�4d�ӧ��B����X,|/�D�H�C�P�m���@$7�T0 k� �DS�HSe2$ 4r1'TP  ��  	   � < �@�<c�צ��B����X,|/�D�H�K�P�n���@$7�T0 k� �LS�PSe2$ 4r1'TP  ��  
   � < �@�Hc�ߦ� B����X,|/�D�H�S�P�n���@$7�T0 k� �XR�\Re2$ 4r1'TP  ��  
   � < �@�Pb���B����\-|/�D�L�W�P�o��@b$7�T0 k� �`Q�dQe2$ 4r1'TP  ��  
   � < �@�Xa���B����\-|/�D�L�_�P�o��@b$7�T0 k� �hQ�lQe2$ 4r1'TP  ��  
   � < �@r`a���B����`-|/�D�L�g�P�p��@b$7�T0 k� �tN�xNe2$ 4r1'TP  ��  
   � < �@rh`����$B����`.|/�D�P�k�P�p��@b$7�T0 k� �L��Le2$ 4r1'TP  ��  
   � < �@rt_����,B����d.|/�D�P�s�P�q��@b$7�T0 k� �J��Je2$ 4r1'TP  ��  
   � < �@r|_���4B����h.|/�D�P�{�E��q��@$7�T0 k� �H��He2$ 4r1'TP  ��  
   � < �@r�^���<B����l/|/�D�T���E��r��@$7�T0 k� �G��Ge2$ 4r1'TP  ��  
   � < �@r�]���HB����l/|/�D�T���E��r��@$7�T0 k� �F��Fe2$ 4r1'TP  ��  
   � < �@r�]���PB����p/|/�D�X���E� r��@$7�T0 k� �E��Ee2$ 4r1'TP  ��  
   � < �@r�\�'��XB����t/|/�D�X���E�s��@$7�T0 k� �D��De2$ 4r1'TP  ��  
   � < �@r�[�/��`B����x0|/�D�\���E�s��B�$7�T0 k� ��C��Ce2$ 4r1'TP  ��  
   � < �@r�Z�7��hB���|0|/�D�\���E�t��B�(7�T0 k� ��C��Ce2$ 4r1'TP  ��  
   � < �@r�Y�?��pB��݀0|/�D�`���E�t��B�(7�T0 k� ��B��Be2$ 4r1'TP  ��  
   � < �@r�Y�G��xB��݄0|/�D�`	��E� t�#�B�,7�T0 k� ��A��Ae2$ 4r1'TP  ��  
   � < �@��X�O���B��݈1|/�D�d	��E�(u�+�B�,7�T0 k� ��A��Ae2$ 4r1'TP  ��  
   � < �@��W�W���B��݌1|/�Fh
��E�0u�7�B�07�T0 k� ��A��Ae2$ 4r1'TP  ��  
   � < �@��V�_���B�#�ݐ1|/�Fh
��E�8u�?�B�07�T0 k� ��@� @e2$ 4r1'TP  ��  
   � < �@��T�o���B�/�ݜ2|/�Fp��E�Dv�O�B�47�T0 k� �?�?e2$ 4r1'TP  ��  
   � < �@��S�w���B�3���2|/�Fp��E�Lv�W�B�87�T0 k� �>�>e2$ 4r1'TP  ��  
   � < �@��R����B�;���2|/�Ft��E�Tv�c�B�<7�T0 k� �=� =e2$ 4r1'TP  ��  
   � < �@�R�����B�?���2|/�Fx��E�\v�k�B�@7�T0 k� �$<�(<e2$ 4r1'TP  ��  
   � < �@�Q�����B�G���2|/�E�|��Edv�s�B�D7�T0 k� �0;�4;e2$ 4r1'TP  ��  
   � < �@�P�����B�O���3|/�E���Elv�{�B�H7�T0 k� �8:�<:e2$ 4r1'TP  ��     � < �@� O�����B�W���3|/�E���EtvЃ�B�L7�T0 k� �@9�D9e2$ 4r1'TP  ��     � < �@�(N�����B�[���3|/�E����E|vЏ�B�P7�T0 k� �H8�L8e2$ 4r1'TP  ��     � < �@�0M�����B�c���3|/�E����E�vЗ�B�T7�T0 k� �P7�T7e2$ 4r1'TP  ��     � < �@�8Lѿ���B�k���4|/�B���'�E�vП�B�X7�T0 k� �X6�\6e2$ 4r1'TP  ��     � < �@�@K�ǚ��B�s���4|/�B���/�E�vЧ�B�\7�T0 k� �`5�d5e2$ 4r1'TP  ��     � < �E�TI�ך�B�����4|/�B���?�E�vл�B�d7�T0 k� �t4�x4e2$ 4r1'TP  ��     � < �E�\H�ߙ�B�����4|/�B���G�E�v���B�h7�T0 k� �|4��4e2$ 4r1'TP  ��     � < �E�dG���B�����5|/�B���O�E�v���B�p7�T0 k� �4��4e2$ 4r1'TP  ��     � < �E�lF���$B�����5|/�B���W�E��v���B�t7�T0 k� �4��4e2$ 4r1'TP  ��     � < �E�tE����,B���� 5|/�B���c�E��v���B�x7�T0 k� �3��3e2$ 4r1'TP  ��     � < �E�|D���8B����5|/�B���k�E��v���B7�T0 k� �2��2e2$ 4r1'TP  ��     � < �E��B���@B�� �5|/�B���s�E��v���B7�T0 k� �1��1e2$ 4r1'TP  ��     � < �E��A���HB�� �5|/�B���{�E��u���B7�T0 k� �-��-e2$ 4r1'TP  �     � < �F��?�'��XB�� �$5|/�B�����I��u��B7�T0 k� �%��%e2$ 4r1'TP ��    � < �F��>�/��`B�� �,5|/�B�����I�u��B7�T0 k� �!��!e2$ 4r1'TP ��    � < F��=�7��hB���44|/�B�����I�u��B¤7�T0 k� ���e2$ 4r1'TP ��    � < F��<�?��tB���<4|/�E�����I�t�#�BҬ7�T0 k� ���e2$ 4r1'TP ��    � < F��;�G��|B���D4|/�E�����I� t�+�BҰ73�T0 k� ���e2$ 4r1'TP ��    � < F��:�O���B���L4|/�E�����I�$t�3�BҸ73�T0 k� ���e2$ 4r1'TP ��    � ; F��9�[���B���T3|/�E�����J,t�;�B��73�T0 k� ���e2$ 4r1'TP ��    � : F��8�c���B��\3|/�E�����J4t�C�B��73�T0 k� �
��
e2$ 4r1'TP ��    � 9 F��7�k���B��d3|/�E�����J<t�K�B��73�T0 k� ���e2$ 4r1'TP ��    � 8 F��6�s���B��l2|/�E�����J@t�W�B��7d T0 k� ���e2$ 4r1'TP ��    � 7 F��5�{���B� �t2|/�E�� ���JHt�_�B��7dT0 k� �����e2$ 4r1'TP ��    � 6 F��4ҋ���B�0ބ1|/�E�!���I�Tt�o�B��7dT0 k� �����e2$ 4r1'TP ��    � 4 F��3җ���B�8ވ0|/�E�!���I�\t�w�I�7dT0 k� �����e2$ 4r1'TP ��    � 2 F� 2ҟ���B�@ސ0|/�E�"��I�`t��I�7d T0 k� �����e2$ 4r1'TP ��    � 0 F�1����B�Lޘ/|/�E�"��I�dt���I7d!T0 k� �����e2$ 4r1'TP ��    � . F�1����B�T�/|/�E�$"��I�lt���I7�$"T0 k� �����e2$ 4r1'TP �    � , QT2����B�\�.|/�E�("��Jpt���I7�(#T0 k� �����e2$ 4r1'TP ��    � * QT3����Ed�.|/�E�0#�'�Jtt���I7�0#T0 k� �����e2$ 4r1'TP ��    � ' QT4�Ӓ�Ex��-|/�E�<#�7�J|t���I# 7�<%T0 k� �����e2$ 4r1'TP ��    � $ QT 5�ۑ�E���,|/�E�D#�?�J�t���I#(7�@%T0 k� �����e2$ 4r1'TP ��    � ! QT$6���E���,|/�E�H#�G�I�t���I#,7�D%T0 k� �����e2$ 4r1'TP ��    �  QT(6���E���+|/�E�P$�O�I�t���I#07�L%T0 k� �����e2$ 4r1'TP ��    �  QT,7���$E���+|/�E�X$�W�I�t���I#47�P%T0 k� �����e2$ 4r1'TP  ��    �  Qd08����0E���*|/�E�\$�_�I�t���E�<7�X%T0 k� �����e2$ 4r1'TP  ��    �  Qd48���8E���*|/�E�d$�k�I�t���E�@7�\%T0 k� �����e2$ 4r1'TP  ��    �  Qd<:���HE�� )|/�E�p#�{�J�t���E�L7�h%T0 k� ����e2$ 4r1'TP  .�    �  Qd@:���PE���(|/�E�x#���J�t��E�P6�p%T0 k� ����e2$ 4r1'TP  ��    �  QdD;���XE���(|/�E�|#���J�t��E�X6�t%T0 k� ����e2$ 4r1'TP  ��    �  QdH<�'��`E���'|/�E��#��J�t��E�\6�|%T0 k� ����e2$ 4r1'TP  ��    �  QtL<�/��lE���'|/�E��"��J�t��E�d5�%T0 k� ����e2$ 4r1'TP  ��    �   QtP=�7��tE���$&|/�E��"��I�t�#�E�h5D�%T0 k� ����e2$ 4r1'TP  ��    ��� QtT=�;��|E���,&|/�E��"��I�t�/�E�p5D�%T0 k� ����e2$ 4r1'TP  ��    ��� Qt\>�K�ҌE� �<%|/�E��! ��I�t�?�E�|4D�%T0 k� ����e2$ 4r1'TP  ��    ��� Qt`?�S�ҔE��D$|/�E��  ��I�t�G�E��3D�%T0 k� ����e2$ 4r1'TP  ��    ��� Qt`@�W�ҜE��L#|/�E��  ��J�t�O�E��2Ę%T0 k� ����e2$ 4r1'TP  ��    ��� Qtd@�_�ҤE��T#|/�E�� ��J�t�W�E��2Ę$T0 k� ����e2$ 4r1'TP  ��    ��� QthA�c�	�B�$�\"|/�Eô ��J�t�_�E��1Ĕ$T0 k� ����e2$ 4r1'TP  ��    ��� QtlA�k�	�B�,�d!|/�Eü ��J�t�g�E��0Ĕ#T0 k� ����e2$ 4r1'TP  ��    ��� QttB�w�	�B�@�p |/�E�� ��I�t�{�E��/Ԑ"T0 k� ����e2$ 4r1'TP  ��    ��� QttC��	�B�H�x|/�E�� ��I�t҃�E��.Ԑ"T0 k� �~��~e2$ 4r1'TP  �    ��� QtxCネ	�B�P߀|/�C���I�t���E��-Ԍ!T0 k� ����e2$ 4r1'TP  ��    ��� Qt|D㋍	"�B�X߈|/�C���I�t���E��,Ԉ!T0 k� ����e2$ 4r1'TP ��    ��� Qt�D㏍	"�B�`ߐ|/�C���I�t���E��+Ԅ T0 k� ��Íe2$ 4r1'TP ��    ��� Qt�E�	"�B�lߘ|/�C���@�t���Eü*�� T0 k� �Ò�ǒe2$ 4r1'TP ��    ��� Qt�F�	"�B�|ߤ|/�C��+�@�t���E��(�x!T0 k� �˝�ϝe2$ 4r1'TP ��    ��� Qt�F�	�B��߬|/�C��3�@�t���E��&�x!T0 k� �Ϣ�Ӣe2$ 4r1'TP ��    ��� Qt�G�	 B���|/�C��;�@�t���E��%�t"T0 k� �ӧ�קe2$ 4r1'TP ��    ��� Qt�G	��	B���|/�C��C�@c�t���E��$�p"T0 k� �׬�۬e2$ 4r1'TP ��    ��� Qt�H	��	B����|/�C��K�@c�t���C��#�l"T0 k� �۱�߱e2$ 4r1'TP ��    ��� Qt�I	Ï	B����|/�C��X@c�tr��C��#�d#T0 k� ����e2$ 4r1'TP ��    ��� Qt�I	Ǐ	#E����|/�C��!`@c�tr��C��"�`$T0 k� ������e2$ 4r1'TP ��    ��� Qt�I	ˏ	#E����|/�C��!hCC�tr��C��!�`$T0 k� ������e2$ 4r1'TP �    ��� Qt�ICϐ	# E��O�|/�C��!pCC�tr��C�� �\$T0 k� ������e2$ 4r1'TP �    ��� Qt�JCې	#,E��	O�|/�E3�!�CC�s�C���T%T0 k� ������e2$ 4r1'TP ��    ��� Qt�JC� 0E��	O�|/�E3��CC�s�C���T&T0 k� ������e2$ 4r1'TP ��    ��� Qt�KC� 4E��	@|/�E4 
�CC�r�C���P&T0 k� �����e2$ 4r1'TP ��    ��� Qt�K��� 8B@�	@|/�E4	�CC�q#�C���L&T0 k� ����e2$ 4r1'TP ��    ��� Qt�K�� @BA 
@|/�E4�
CC�p3�C���H'T0 k� ����e2$ 4r1'TP ��    ��� Qt�L�� DBA
@ |/�E4�CC�o;�C���D'T0 k� ����e2$ 4r1'TP ��    ��� Qt�L�� HBA
@$|/�E4 �CC�o�C�C���@(T0 k� ����e2$ 4r1'TP �    ��� Qt�L�� LBA
@,|/�CD �CS�n�K�C���<(T0 k� $���e2$ 4r1'TP ��    ��� Qt�M�� PBA 
@0|/�CC���CS�m�S�C���8)T0 k� $���e2$ 4r1'TP ��    ��� Qt�M�� XBA0
@<
|/�CC���CS�k�_�C��d0)T0 k� $���e2$ 4r1'TP ��    ��� Qt�M�#� \BA4@D	|/�CC� ��CS�j�g�C��d,)T0 k� $���e2$ 4r1'TP ��    ��� Qt�N�'� \BA<@H|/�E3����CS�i�o�C��d(*T0 k� #� �  e2$ 4r1'TP ��    ��� Qt�N�+� `BAD@P|/�E3����CS�h�w�C��d$*T0 k� ����e2$ 4r1'TP ��    ��� Qt�N�+� dBAL@T|/�E3����CS�f��C��d *T0 k� ����e2$ 4r1'TP ��    ��� Qt�N�/� hBAP@\|/�E3����CS�e	�E3�d*T0 k� ����e2$ 4r1'TP ��    ��� Qt�O�7� pBA\@h|/�K����CS�b	�E3�	d+T0 k� ����e2$ 4r1'TP ��    ��� Qt�O�;� tBAd@l|/�K����Cc�a	�E3�d+T0 k� 3�����e2$ 4r1'TP ��    ��� Qt�O�;� xBAl@p|/�K����Cc�_	�E3�d+T0 k� 3�����e2$ 4r1'TP ��    ��� Qt�O�?� xBAp@x|/�K���� Cc�^	�E3�d,T0 k� 3�����e2$ 4r1'TP ��    ��� Qt|P�C� |BAx@||/�K����$Cc�\
��E3�d,T0 k� 3�����e2$ 4r1'TP ��    ��� Qt|P�G� �BA�@�|/�K����4Cc�Y
��E3�d ,T0 k� 3�����e2$ 4r1'TP ��    ��� Qt|P�K� �BA�@�|/�K����8Cc�W
��K��c�-T0 k� ������e2$ 4r1'TP ��    ��� Qt|Q�O� �BA�@� |/�K����@Cc�V
ǫK��c�-T0 k� ������e2$ 4r1'TP ��    ��� QtxQDO� �BA�@� |/�K����DCc�T	�˫K���c�-T0 k� ������e2$ 4r1'TP ��    ��� QtxQDS� �BA�@��|/�K����LCc�R	�ϪK���c�-T0 k� ������e2$ 4r1'TP  ��    ��� QtxQDW� �BA�@��|/�K����XCc�N	�שK���c�.T0 k� ������e2$ 4r1'TP  -�    ��� QtxRD[� �BA�@��|/�K����\Cs�L	�۩K���c�.T0 k� #�����e2$ 4r1'TP  ��    ��� QttRD_� �BA�@��|/�K����dCs�J
�K���c�.T0 k� #�����e2$ 4r1'TP  ��    ��� QttRD_� �BA�@��|/�K����hCs�H
�K���c�.T0 k� #�����e2$ 4r1'TP  ��    ��� QttRDc� �BA�@��|/�K����pCs�F
�K���c�.T0 k� #�����e2$ 4r1'TP  ��    ��� QttSDg� �BA�@��|/�K����x Cs�B
�K���c�/T0 k� #�����e2$ 4r1'TP ��    ��� QtpSDk� �BA�@��|/�K����� Cs�?	��K���c�/T0 k� ������e2$ 4r1'TP ��   ��� QtpSDk� �BA�@��|/�K�����!Cs�=	���K���c�/T0 k� ������e2$ 4r1'TP ��    ��� QtpSDo� �BA�@��|/�K�����!Cs�=	���K���c�/T0 k� ������e2$ 4r1'TP ��    ��� QtpSDo� �BA�@��|/�K�����"Cs�=	���K���c�.T0 k� ������e2$ 4r1'TP ��    ���                                                                                                                                                                             � � �  �  �  c A�  �J����  �      � \��9
 ]�$�$� � � ^�$         �]�     ^�`     a��                  8          O      ���   			          ��R   $ $     ���    ����y    ��1   	                      �      ���   0	&          (;�            �z     ( �7    �                �          .�  �  ���   8
	            $ $      ��     	1 ��@     :�                A�$           �      ���   @	           ���   $ $     . rӨ    ��() r��    �p�                 �$          ��     ���   84         ����  ��	      B�Av    �����Av                             ���I               }  ���     

 0            ��� D D     Vo�    ���h�    _��              	��          &P�    ��@  H          ���S  K K     j ���    ��|� ���    �� h               		�� �         � �    ��@  8
          �� M M       ~ �:r    ��s� �+-    	V�               ��          {b     ��@  

'           ����  � � 	  ��8    ���g�     A��             	��         	 ��     ��`   X
         ��q � �	   � �Dv    ���� �I>    ����               c��          
 ���    ��h   8

           4�j ��     � �\     4�� �r(    ���                     ���r              �  ��@   0 0                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         ���  ��        � �m�    ��,; �ri    ���� "                x                j  �    
   �                         ��    ��        � �      ��   �           "                                                �                          � � r� � � � ��� � �         	   
     
 ~    y �� 1��       1� m@ 1� m` 1� `m� S� `w@ Td x  T� x  T� x@ )� `j� *D k� �D  k� ��  k� 
�� V  
�| V  @  \� @D  ]  :d q  >D `[� ? @\� ?� ]  / `^@ /� _  /� _  0 _@ �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �d �Q` �� �R����� ����� � 
�� W� 
�| W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����   �����   ������  
�fD
��L���"����D" � j  "  B   J jF�"     
�j � � 
��
��
��"     "�j��   * �
� �  �  
� ����  ��     � �      ��    ��     �      ����  ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �&      �� �) ���        �6T ���        �        ��        �        ��        �   *�     ���g�        ��                         5�$ 8  80� ��                                     �                ����            
�� �
���%��  ��  2����           14 Theoren Fleury      0:01                                                                        5  5     �dC.t C6 �K:' K"J � �
 � � �k� � �k� � 	k� �
k� � �k� � cj � ck �cl �CM �k~ � � k� � �c�U � c�U � c�P � c�e �c� � � c� � �kV � � k\ � �	� �	�+ �� ��= �J�� �J�q � B�
 � !B�""� � #"� �
$� �
%
� � �&"� � '"� �("� �)*�*"� � +"� �
,� �
-
� � � ."H � �/" � � 0!� � � 1"K � �2"( � � 3"O � �4"* | �5"8 | � 6" � �7!� � �8" � �9" � �:" �;!� �<"D �=*d � >"E t �  "G �                                                                                                                                                                                                                         �� P   �     �     @ 
             W P E ^  ��        
            �������������������������������������� ���������	�
��������                                                                                          ��    �?�   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, /� * � ��@�@���@q�@����                                                                                                                                                                                                                                                                                                                                � ��]�                                                                                                                                                                                                                                     
     X  	  &    ��  :�J      U  	                           ������������������������������������������������������                                                                      	                                                                   �    6    �        g,      C�       C          
     ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� �������            �             	     �    4     �  4�J       �                             ������������������������������������������������������                                                                     
                                                                   �  �           �             �   �           	 
     ��  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���             C                                                                                                                                                                                                                                       	                                                              
        �             


             �  }�  � �    ������������  '���������  +	����������������       ������������  'q������������������������������������                                                 N�     Ry  'w                     ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" R > / 	                                � �&p �\                                                                                                                                                                                                                                                                                      	�)n1n  �        k      c                              `      l                                                                                                                                                                                                                                                                                                                                                                               j                        0 �  
>�  J�  2�  2�  J`�  ����(���Z��� ���:����(�_����������c�����J                      �% q           �   & AG� �  r   
              �                                                                                                                                                                                                                                                                                                                                     S H                         !��                                                                                                                                                                                                                            Y   �� �� Ѱ�      �� 7  �� 
����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� ���������  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���             $������������������������������������������������������eU���U����������������l��lfl�l�ff�Uw��U��f���������ˊ����ff�lf�l���f��˚�˛�����������l����fj�l���l���ƛ�̩���������������������������i������������������������������������lw�vffl�fjfl���Ōj��lf�|�w�yx��l�ll���lfffefff�ffff�fffk�ff�l��ƥWˆk���f��fl��flf���l�l�llff�̼gu���U\l�ʉƬ�U�l������l�ll����f�������[ʩ�U���uW���U��luz��ǚ����������������������������������x���ywU����Y����i���f���ǬƇ�\f��˺yflˈ�fl�W�f̗U����[f˘wff��ffl̬��lk��f����ff��f��̶��̖������l��Ƽ�̦�f̶��fl�����l��l�l��lk��l�ʩ�̺��˚�ll��lʫ�̺��̻�����������������������������������wZf�Wu��ww{���x��j�W�ʉx��zX�x��k����w�ɇ�w�����������������y�xvjll�eVk��[��UZU�u�u�uWx��xx�UX��k�l���l��lk�x�ʖgƻ��l�u{k�uvk��ɪ��ɛ�������������ʚ��ɚ������������������������ɚ�������̗x��|l��z�f�W��kX���w����xy�������������x��x�xxy�x�y�������z������x��Ux��U{��u\l��YƗ�Ux���Uˇu�jwU�xffh�ff�fu��hY̪Uff�Vf��ffl�flƵ�����������������������������xx�u{��X��̼�����������������������ʈ���Ǌ��ɇ��̸���iU̶hY���X�ƺw���f��f��˅U�uU�Uw������������ʊ�x�ywy�[X�wY��xW���{�������ȫ���fff�f�Ƹl[��Ō�̈���|�����������Wxyw��UUgWx�ƵXZ�Ɨw��ky���g�������    4   !   D     ��                       7     �   �����J����    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �΀ �� �    � �N ^$    ��H     ��   i  ��   �   ���t����������J������    # ��     ^   ��  ^ >�������� J  ^ ^   ��  ^   i  ��   �    >   �����   �z � �N ^$  �   �   
              [� � ��  o� � ��� �� � ��� �$ #  ��T  �      �       �������2����   g���        f ^�         ��m��            ��9l���2�������J������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                               	                 �  ��� �UU���U              �	���UUU�UUUUUU      	� ��U�UUUUUUUUUUUUUUUUUUU    ��� U^��UUU�UUU^UUUUUUUUUUUU            �   �   ^�  U�  UY�    � 	UU 	��  	�  	�  �^ 	��    �	UY�������UUUUUUU��UU��UU�U�UUUUUUUUUUUUUUUUUUUUUUUUUUUU^UUUYUU^�U^� U� ^�  �  ��  �   �   ��UU ��U �U  �U  ��            U^� UU� UU� UU� ���                    	   �       	   	   	    �UUU�UU���U  	�� �����U�UUU�UUUUUUYUUUYUUUYUUU^UUU^UUUUUUUUUUUU�   �   �   �   �   � �^���U^��            	����UUU�UUU�UUUUUU^            ��  U�  Y�  �  �      �   �   �   	                ���Y���U��Y�^�U��U ��^ 	� 	� UUUU�UUUUUUUU^�U^����� �        UUUUUUUUUUUUUUUUUUUU�������    UUU�UU^�UU�U� Y�  ��          �                               wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                                    �����   �   �   �   ����                                     	�  		  	 � 	 	 	   	   	   	   	  ��                  ��   	   	   	   	   	   	 	 	 � 		  	�                 �   	    �   	    �   	    �   	   	   �  	   �  	   �  	   �                                      
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            "! "   "      ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ ""   "! " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       "! "   "      ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                              	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                         �   �     �   �        �   �"/� ����                                     ��  ��  �                  �  ������� ��                                                                                                                                                                                                            �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �                  ���� ���  ��    �            �   ������  ��                      �   �                      �������  ���    �                    ��  ��  ���  �  �  �   �   ��  �                            �   ���                            �   �                                                                                                    �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   2 1220!2 #!0 #        �   �   �   �   �   �   �     �     �     �   "   "                                      �       ����������                                ��  ��  ���                                                                                                                                                                                                       �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   ɪ  ��� ټ� �̰ �̰ ��� ��  ��              �   ������  ��                   �                        ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                      �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                        �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �   �" �!  �  �� �   �                �  �� Ș ��  ��  �                �   �                                                                                                                                                                                                                ̰ ˻ ���wݛk}�gz� w��  ��  ��  ��  ��  ,�  "�  �  ,�  "�  ..  ..  �  �   �                        �   �   ̰  ��  ��  ��� ��� �ܘ �ل@�؊@�4�@�H�@�D �@ �H� "H�""C�"ˋ" �" ��" "��� �  �                     ��  �                                         �   �   ��  ��  ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����            �  �  ��  �   �   �                         ���                � ���� ��   � � �                                                                                                                                  �  �  ��� �                     �  �˰ ˻� w�� k}� gw� z�� ��� ��� ��� ��� ��  �� ���"�ȍ�̽�"��4  4H H� D�� X�D X� Ą  ��" 
��  "  "" ""  ��    �   ��  ��  ��  ��  ��  ̐  ��  �0  �0  �0  T   C   3   �   ��  +�  ""  ""� /�� / �    ��                 �   �                           �   �  "������"    /   �  �   ��               ����                         � "            � "�",�"+� ",                       "  .���"    �     �                         � ���� ��   � � �                           �   �                                                                                                    ˰ ̻ ̻ �� {�  �� 
�� ��� ��� ������
���	��ܻ̍ݻ���"� 8"  8  �  D�  H�  X�  ��  �   �          "  "     �                        ��  ��� �̺�̻����ۻ�˽��̽��̝ ̙� �30 �EP �U@ �T0 EC0 T3  C:  K�  �"  �"/ ����˽� �"� "" �""� � �� ��      �   �� ��  �"  �            �   �"  ""  !� �� ��  �               �   ������  ��           �   �    �   �       �   �   �                .                      ��  ��  ���       +  "  "     �  �                                                                                                                                                                       �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                        � ��                  �  �˰ ��� �wp ���                                                                                                                                                                               � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �         ��                                 � ���� ��   � � �                           �   �                                                                                                   ����������ݼ������ى����.(����M���M D � ��� �"( ��� �� �� �  �  �   �   �  �   ��  ��� ؼ̰ڛ�˺������ɪ�۸��Ȕ͙̄̄͜Mڜ��̩U�̴@��ݿ��������ɉ��ɋ�������������𻻲  "/  ��   �   �   �   �           ��  �     �  �  �      �   �   �   ��      �   ��          ��  ��� ��  �                                        �� ��  �� ��  "/������ � �               �   �                     �     �                                      � ����ݼ� ����                                                                                                                                                                             �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""��������������������""""������DDM�D��""""�������MM�M�M""""��������DD�A��""""�������MAA�MA""""��������AA�A""""����������M�MA""""������������M���M���M���"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUQUUQUUUUUUQUUUUUUUU3333DDDDUUUUDEEDDTEUUUU3333DDDDAEAEQQUDTDUUUU3333DDDDQUQUQDUDDUUUU3333DDDDAADAUAUEDUTUUUU3333DDDDADAEAQAUEDUTUUUU3333DDDDUDUQEUQUUQUEUDUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��           	 
          
        ((((((( 
	(((( """"��������AA�A             ! " # $ % & '   ( $ % ) ! " # * ('(&(%($(#("(! (((ADA�LL��L�D����3333DDDD + , -   . / 0 1  	 2         3       4 (((((((2	10/(.(-(,(+LL����������D����3333DDDD 5 6   7   8 9 1 :   $ % ) ! " #   ; ) ! " # $ % ) (#("(!()(%($ :198(((7(6(5""""����������A������    <     = 8 0 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>108(=((( (<""""�������I�I������ L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L""""�������I��D���I�������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7�D�M�D���M������3333DDDD  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`D�M�A�����MD�����3333DDDD 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
""""�����AMAD������ w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw""""������������������ w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xwwfFfFDfFFfFffdFffff3333DDDD + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+DDFFDfFFfdFffff3333DDDD � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(�""""wwwwwwwGGD � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(�""""wwwwwwqwAqwAwA �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(�""""wwwwqwqAwAqAqAq = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=A�A�A�A��LD�����3333DDDD    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( �A�LDL�L�D�L�����3333DDDD x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx""""wwwwwwDGAD w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww""""wwwwqqDAAq  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(""""wwwwwwwGGwGGwGwGw �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((�UQUUQUUQUUQUUUDUUUUU3333DDDD ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`DEQQUUDUTEUUUU3333DDDD M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M""""������������������������ � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(�""""�������DAADAI � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(��A�AM�M�DM��M334CDDDD 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5DD����M��DM�����3333DDDD x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x""""wwwwwwDGqGq w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwwGwwDGwwwwwwww + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+ADAH�DJ�H�H�����3333DDDD � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(��H��J�AD�DH�D����3333DDDD333333333333333333333333333333333333333333333333333333333333����  
�fD
��L���"���""""�������DD������D" � j  "  B   J jF� ����
��� �����
���� ����
��� �����
��� 0 q""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqdC.t C6 �K:' K"J � �
 � � �k� � �k� � 	k� �
k� � �k� � cj � ck �cl �CM �k~ � � k� � �c�U � c�U � c�P � c�e �c� � � c� � �kV � � k\ � �	� �	�+ �� ��= �J�� �J�q � B�
 � !B�""� � #"� �
$� �
%
� � �&"� � '"� �("� �)*�*"� � +"� �
,� �
-
� � � ."H � �/" � � 0!� � � 1"K � �2"( � � 3"O � �4"* | �5"8 | � 6" � �7!� � �8" � �9" � �:" �;!� �<"D �=*d � >"E t �  "G �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3�����������������������������������������#��<�Z�K�\�K��6�G�X�S�K�X� � � � � � � � �-�2�3�������������������������������������������=�N�K�U�X�K�T��0�R�K�[�X�_� � � � � � �-�1�B�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������-�2�3� �� �������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�1�B� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            