GST@�                                                            \     �                                               ��a      �     ?         ����e ����J�������������������        �g     #    ����                                d8<n    �  ?     l�����  �
fD�
�L���"����D"� j   " B   J  jF�"     "�j  " ���
��
�"    
 �j�
�
  
  ��
  Y                                                                               ����������������������������������       ��    =o 0b 4o 1 4  +c  c 'c      �     	  
     �	G �7� �V( �	(                 nn 	1         :8�����������������������������������������������������������������������������������������������������������������������������=  0b  4  11                                         �  �  �  �                  �  
1          = �����������������������������������������������������������������������������                                ��  �       _�   @  #   �   �                                                                                '    	n1n  
1�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    �P#���L�/�D�ӊ#3�Mg�A��PA��� d����"s��T0 k� �C��G�"�2't ��1"t'!  ��F    ������L"���L�+�D�Ӌ#3�M_�A��PA��� d#����"s��T0 k� �;��?�"�2't ��1"t'!  ��F    ������D ���L�'�D�ό#3�mW�A��PA��� d#����"s��T0 k� �3��7�"�2't ��1"t'!  ��F    ������@���L��D�ό#3�mO�A��PA��� d#����"s��T0 k� �+��/�"�2't ��1"t'!  ��F    ������<���L��D�ˍ#3�mG�A��PA��� d#����"s��T0 k� �#��'�"�2't ��1"t'!  ��F    ������4���L��D�ˎ#3�m?�A��QA��� d#����"s��T0 k� ����"�2't ��1"t'!  ��F    ������0���L��L^Ǐާ�#3�m7�A��QA��� d'����"s��T0 k� ����"�2't ��1"t'!  ��F    ������,���E>�L^Ǐާ�#3�]/�A��QA��� d'���3��T0 k� ����"�2't ��1"t'!  ��F    ������$���E>�L^ǐާ�#3�]'�A��QA��� d'���3��T0 k� ����"�2't ��1"t'!  ��F    ������ b��E>�L^Ñޫ�#3�]#�A��QA��� d'���3��T0 k� �����"�2't ��1"t'!  ��F    ������b��E>�L^Òޫ��3�]�A��QA��� d'���3��T0 k� ������"�2't ��1"t'!  ��F    ������b��E=��L^��ޫ��3�]�A��QA� d'���3��T0 k� ������"�2't ��1"t'!  ��F    ������b��E-��L^�� ����3�M�A��QA� d'���3��T0 k� ������"�2't ��1"t'!  ��F    ������b��E-��L^�� ����3�M�A��QA� d+���3��T0 k� ������"�2't ��1"t'!  ��F    ������
b��E-��L^�� ����3�L��A��RA�� d+���3��T0 k� ������"�2't ��1"t'!  ��F    �����_b��E-�L^�� ����3�L��A��RA�� d+���3��T0 k� ������"�2't ��1"t'!  ��F    �����_ b��E-�L^�� ����3�L��A��RA�� d+���3��T0 k� ������"�2't ��1"t'!  ��F    �����^�b��E-�L^�� ����3�l��A��RA�� d+���3��T0 k� ������"�2't ��1"t'!  ��F    �����^�R��E-�L^�� ����3�l��A��RA�� d+���"���T0 k� ������"�2't ��1"t'!  ��F    �����^�R��E�L^�� ����3�l��A��RA�� d/���"���T0 k� ������"�2't ��1"t'!  ��F   �����^��R��E�Ln�� ����3�l��A��RA�� d/���"���T0 k� ������"�2't ��1"t'!  �F    �����^��R��E�Ln�� ����3�l��A��RA�� d/���"���T0 k� ������"�2't ��1"t'! ��O    �����^��R��E�Ln�� ����3�|��A��RA�� d/���"���T0 k� ������"�2't ��1"t'! ��O    �����^����E�Ln�� ����3�|��A��RA�� d/���"���T0 k� ������"�2't ��1"t'! ��O    �����^����E�Ln�� ����3�|��A��SA�� d/���"���T0 k� �w��{�"�2't ��1"t'! ��O    �����^����E�Ln�� ����3�|��A��SA�� d/���"���T0 k� �k��o�"�2't ��1"t'! ��O    �����^����E�Ln�� ����3�|��A��SA�� d/���"���T0 k� �[��_�"�2't ��1"t'! $�O    �����^����B��Ln�� ����3����A��SA�� d3���"���T0 k� ,_��c�"�2't ��1"t'! ��O    �����^����B��Ln�� ����3����A��SA�� d3���"���T0 k� ,c��g�"�2't ��1"t'! ��O    �����n����B��Ln�� ����3����A��SA�� d3���3��T0 k� ,c��g�"�2't ��1"t'! ��O    �����n����B��Ln�� ����3����A��SA�� d3���3��T0 k� ,g��k�"�2't ��1"t'! ��O    �����n����B��Ln�� ����3����A��SA�� d3���3��T0 k� ,k��o�"�2't ��1"t'! ��O    �����n����B��Ln�� ����3����A��SA�� d3���3��T0 k� ,k��o�"�2't ��1"t'! ��O    �����n��"��B��Ln�� ����3����A��SA�� d3���3��T0 k� �o��s�"�2't ��1"t'! ��O    �����n��"��B��Ln�� ����3����A��SA�� d3���3��T0 k� �s��w�"�2't ��1"t'! ��O    �����n��"��B��Ln�� ����3����A��SA�� d7���3��T0 k� �w��{�"�2't ��1"t'! ��O    �����n��"��E��Ln�� ����3����A��TA�� d7���3��T0 k� �w��{�"�2't ��1"t'! ��O    �����n��"��E��Ln�� ����3����A��TA�� d7���3��T0 k� �{���"�2't ��1"t'! ��O    �����n��"��E��Ln�� ����3���A��TA�� d7���3��T0 k� <����"�2't ��1"t'! ��O    �����n��"��E��Ln�� ����3��{�A��TA�� d7���3��T0 k� <����"�2't ��1"t'!  ��O    �����n��"��E�Ln�� ����3��w�A��TA�� d7���3��T0 k� <�����"�2't ��1"t'!  ��O    �����n��"��K��Ln�� ����3��s�A��TA�� d7���3��T0 k� <�����"�2't ��1"t'!  ��O    �����n��"��K��Ln�� ����3��o�A��TA�� d7���3��T0 k� <�����"�2't ��1"t'!  .�O    �����n��"��K��Ln�� ����3��k�A��TA�� d7���3��T0 k� ������"�2't ��1"t'!  ��O    �����n��"��K��Ln�� ����3��g�A��TA�� d7���3��T0 k� ������"�2't ��1"t'!  ��O    �����n��"��K��Ln�� ����3��c�A��TA�� d;���3��T0 k� ������"�2't ��1"t'!  ��O    �����n��"��K��Ln�� ����3��_�A��TA�� d;���3��T0 k� ������"�2't ��1"t'!  ��O    �����n��"��K��Ln�� ����3�[�A��TA�� d;���3��T0 k� ������"�2't ��1"t'!  ��O    �����n��"��K��Ln�� ����3�W�A��TA�� d;���3��T0 k� ,�����"�2't ��1"t'!  ��O    �����n��"��K��Ln�� �î�3�S�A��TA�� d;���3��T0 k� ,�����"�2't ��1"t'!  ��O    �����n��"��K��Ln�� �î�3�O�A��TA�� d;���3��T0 k� ,�����"�2't ��1"t'!  ��O    �����n��"��K��Ln�� �ï�3�O�A��UA�� d;���3��T0 k� ,�����"�2't ��1"t'!  ��O    �����n��"��K��Ln�� �ï�3�K�A��UA�� d;���3��T0 k� ,�����"�2't ��1"t'!  ��O    �����n��"��K�#�Ln�� �ï�3�G�A��UA�� d;���3��T0 k� ������"�2't ��1"t'!  ��O    �����n��"��K�'�Ln�� �ï�3�C�A��UA�� d;���3��T0 k� ������"�2't ��1"t'!  ��O    �����n�"��K�'�Ln�� �ï�3�?�A��UA�� d;���3��T0 k� ������"�2't ��1"t'!  ��O    �����n�"��K�+�Ln�� �ï�3�;�A��UA�� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����n{�"��K�/�Ln�� �ǰ�3�7�A��UA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����nw�"��K�/�Ln�� �ǰ�3�3�A��UA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����ns�"��K�3�Ln�� �ǰ�3�/�A��UA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����ns�"��K�7�L^�� �ǰ�3�+�A��UA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����no�"��K�7�L^�� �Ǳ�3�'�A��UA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����no�"��K�;�L^�� �Ǳ�3�'�A��UA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����nk�"��K�;�L^�� �Ǳ�3�#�A��UA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����nk�"��K�?�L^�� �Ǳ�3��A��UA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����ng�"��K�?�L^�� �Ǳ�3��A��UA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O   �����ng�"��K�C�D��� �˱�3��A��UA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����nc�"��K�C�D��� �˱�3��A��VA��� d?���3��T0 k� ������"�2't ��1"t'!  ��O    �����nc�"��K�C�D��� �˲�3��A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    �����^_�"��K�G�D��� �˲�3��A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    �����^_�"��K�G�D��� �˲�3��A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    �����^[�"��K�K�D��� �˲�3��A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    �����^[�"��K�K�D��� �˲�3��A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    �����^W���K�O�D��� �˲�3��A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    �����^W���K�O�D��� �˲�3��A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������S�ǿK�S�A��� �˳�3��A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������S�ǿK�S�A��� �˳�3���A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������S�ǿK�S�A��� �ϳ�3���A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������O�ǿK�W�A��� �ϳ�3���A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������O��ǿK�W�A��� �ϳ�3���A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������K��ÿK�[�A��� �ϳ�3���A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������K��ÿK�[�A����ϳ�3���A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������K��ÿK�[�A����ϳ�3���A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������G��ÿK�_�A����ϴ�3���A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������G�⿿K�_�A����ϴ�3���A��VA��� dC���3��T0 k� ������"�2't ��1"t'!  ��O    ������C�⿿K�_�A����ϴ�3���A��VA��� dG���3��T0 k� ������"�2't ��1"t'!  ��O    ������C�⻿K�c�A����ϴ�3���A��VA��� dG���3��T0 k� �����"�2't ��1"t'!  ��O    ������C�⻿K�c�A����ϴ�3���A��VA��� dG���3��T0 k� �����"�2't ��1"t'!  ��O    �����?�ⷿK�c�A����ϴ�3���A��VA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    �����?�ⷿK�g�A����ϴ�3���A��VA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    �����?�⳾K�g�A����ϴ�3���A��WA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    �����?��K�g�A����Ӵ�3���A��WA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    �����?��K�k�A����ӵ�3���A��WA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    �����;��K�k�A����ӵ�3���A�|WA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    �����;��K�k�A����ӵ�3���A�|WA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    �����;��K�o�A����ӵ�3���A�|WA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    �����;��K�o�A����ӵ�3���A�|WA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    �����;��K�o�A����ӵ�3���A�|WA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    ������?��K�s�A����ӵ�3���A�|WA��� dG���3��T0 k� ����"�2't ��1"t'!  ��O    ������?��Es�A����ӵ�3���A�|WA��� dG���3��T0 k� ���#�"�2't ��1"t'!  ��O    ������?��Es�A����ӵ�3���A�|WA��� dG���3��T0 k� ���#�"�2't ��1"t'!  ��O    ������?��Ew�A����ӵ�3���A�|WA��� dG���3��T0 k� �#��'�"�2't ��1"t'!  ��O    ������C���Ew�A����ӵ�3���A�xWA��� dG���3��T0 k� �#��'�"�2't ��1"t'!  ��O    ������C���E{�A����Ӷ�3���A�xWA��� dG���3��T0 k� �'��+�"�2't ��1"t'!  ��O    ������C��E�{�A����Ӷ�3���A�xWA��� dG���3��T0 k� �+��/�"�2't ��1"t'!  ��O    ������G�w�E��A����Ӷ�3���A�xWA��� dK���3��T0 k� �+��/�"�2't ��1"t'!  ��O    ������G�s�E���A����׶�3���A�xWA��� dK���3��T0 k� �/��3�"�2't ��1"t'!  ��O    ������K�o�E���A����׶�3���A�xWA��� dK���3��T0 k� �/��3�"�2't ��1"t'!  ��O    �����}2PR,'D��F ���|0 �S�F(nDB6��@�r�T0 k� �8x�<x"�2't ��1"t'!  ��    � < �B ~"LR0(D��I ���|0 �S�F$oDB7��@�r�T0 k� �Tv�Xv"�2't ��1"t'! ��    � < �B ~"LR0(D��K ���|0 �S�F$oDB7��@�r�T0 k� �dt�ht"�2't ��1"t'! ��    � < �A�"HR0(D��M ���|0 �S�E�$pDB7�'�0�r�T0 k� �ps�ts"�2't ��1"t'! ��    � < �A��"HR0(Eq�N ���|0 �S�E�$qDB7�+�0�r�T0 k� ��r��r"�2't ��1"t'! ��    � < �A�"HR0(Eq�P ���|0 �S�E�(rDB7�3�0�s�T0 k� ��p��p"�2't ��1"t'! ��    � < �Q��DR0(Eq�R ���|0 �S�E�(rDB8�7�0�s�T0 k� ��o��o"�2't ��1"t'! ��    � < �Q��DR0(Eq�T ���|0 �S�E�(sDB8�?�0�r�T0 k� ��n��n"�2't ��1"t'! ��    � < �Q��D	UD0(Eq�V ���|0 �S�E�,tDB8�C�0�r�T0 k� ��m��m"�2't ��1"t'! ��    � < �Q�~�D
UD0)Eq�W ���|0 �S�E�,uDB8�G�0�r�T0 k� ��k��k"�2't ��1"t'! ��    � < �Q�~�DUD0)Eq�Y ���|0 �S�E�0vDR8CO�0�r�T0 k� ��j��j"�2't ��1"t'! ��    � < �a�~�DUD0)Eq�[ ���|0 �S�E�0wDR8CS�0�r�T0 k� ��i��i"�2't ��1"t'! ��    � < �a�~�@UD0)Ea�] ���|0 �S�B�4xDR8CW�0�r�T0 k� ��g��g"�2't ��1"t'! ��    � < �a�~�@UD0)Ea�_ ���|0 �S�B�4yDR8C_�0|r�T0 k� � f�f"�2't ��1"t'! ��    � < �a�}�@UD0)Ea�c a��|0 �S�B�<zA�8Cg� pr�T0 k� �d� d"�2't ��1"t'! ��    � < �a�}"@UD0)Ea�e a��|0 �S�B�@{A�8Co� lr�T0 k� �(b�,b"�2't ��1"t'! ��    � < �a�}"@UD0)Ea�g a��|0 �S�E�D|A�8Cs� hr�T0 k� �8a�<a"�2't ��1"t'! ��    � < �a�|"@UD0*Ea�i a��|0 �S�E�D|A�8Cw� ds�T0 k� �D`�H`"�2't ��1"t'! ��    � < �a�|"@UD0*Ea�j a��|0 �S�E�H}A�8C{� `s�T0 k� �T^�X^"�2't ��1"t'! ��    � < �a�|"@UD4*Ea�j a��|0 �S�E�L}A�8S�� \s"C�T0 k� �`]�d]"�2't ��1"t'! ��    � < �a�}"@UD4*Ea�k a��|0 �S�E�P~A�8S�� Xs"C�T0 k� �p\�t\"�2't ��1"t'! ��    � < �a�~"DUD4*Ea�l a��|0 �S�E�T~A�8S�� Tt"C�T0 k� �|[��["�2't ��1"t'! ��    � < �a�"DUD4*Ea�m a��|0 �S�E�X~A�8S��Pt"C�T0 k� ��Y��Y"�2't ��1"t'! ��    � < �a�"DUD4*Ea�n a��|0 �S�E�\A�8S��Pu"C�T0 k� ��X��X"�2't ��1"t'!  ��    � < �aԀ"DUD4*EQ�o a��|0 �S�E�`A�8S��Lu"�T0 k� ��W��W"�2't ��1"t'!  ��    � < �aԀHUD4*EQ�p ��|0 �S�E�dA�8S��Hu"�T0 k� ��U��U"�2't ��1"t'!  ��    � < �aЀHUD4+EQ�q ��|0 �S�E�hA�8S��Hv"�T0 k� ��T��T"�2't ��1"t'!  /�    � < �aЀL UD4+EQ�q ��|0 �S�E�lA�8S��Dv"�T0 k� ��S��S"�2't ��1"t'!  ��    � < �aЁL!UD4+EQ�r ��|0 �S�E�pA�8S��Dw"�T0 k� ��R��R"�2't ��1"t'!  ��    � < �àP#UD4+EQ�r ��|0 �S�E�tA�8S��Dw��T0 k� ��P��P"�2't ��1"t'!  ��    � < �̀P$UD4+EQ�r ��|0 �S�E�x~A�8c��Dw��T0 k� ��O� O"�2't ��1"t'!  ��    � < �ȀT%UD4+EA�rA��|0 �S�E�|~A�8c���@x��T0 k� �N�N"�2't ��1"t'!  ��    � < �ȀX'UD4+EA�rA��|0 �S�CB�}A�8c���@x� T0 k� �(K�,K"�2't ��1"t'!  ��    � < ��\)UD4+EA�sA��|0 �S�CB�}BB8c���@y�T0 k� �4J�8J"�2't ��1"t'!  ��    � < ����`*UD4+EA�sA��|0 �S�CB�|BB8c���@y�T0 k� �DI�HI"�2't ��1"t'!  ��    � < ����d+UD4,C��sA��|0 �S�CB�|BB8c���@y�T0 k� �PG�TG"�2't ��1"t'!  ��    � < ����h,UD4,C��s��|0 �S�CB�{BB8c���Dz�T0 k� �\F�`F"�2't ��1"t'!  ��    � < ����l-UD4,C��r��|0 �S�CB�zBB8c���Dz�T0 k� �lE�pE"�2't ��1"t'!  ��    � < ���~�p.UD4,C��r��|0 �S�E��z@8c���Dz�T0 k� �xD�|D"�2't ��1"t'!  ��    � < ���~�t/UD8,C��r��|0 bS�E��y@8c���H{� T0 k� ��B��B"�2't ��1"t'!  ��    � < ���~�x0UD8-C��r��|0 bS�E��x@8s���H{� T0 k� ��A��A"�2't ��1"t'!  (�    � < �A�~�|1UD<.C��q���|0 bS�E��w@8s���H{�!T0 k� Đ@��@"�2't ��1"t'!  .�    � < �A�}��2UD<.C��q���|0 bS�E��v@8s���L{�!T0 k� Đ?��?"�2't ��1"t'!  ��    � < �A�}��3UD</C��q���|0 bS�EB�u@b8s���P|�"T0 k� Č=��="�2't ��1"t'!  ��    � < A�}��4UD@/C��p���|0 S�EB�t@b8s���P|t"T0 k� Ĉ<��<"�2't ��1"t'!  ��    � < �}��6UD@0C��o���|0 S�EB�r@b8����X}t#T0 k� Ā:��:"�2't ��1"t'!  ��    � < �}��7UDD1C��n���|0 S�EB�q@b8����X}t#T0 k� �|9��9"�2't ��1"t'!  ��    � < �}��8UDD1C��n���|0 S�E2�pCB7����\}t$T0 k� �x7�|7"�2't ��1"t'!  ��    � < �}��9UDD2C��m���|0�W�E2�nCB7����`}t$T0 k� �x6�|6"�2't ��1"t'!  ��    � < �|��:UDH2C��l���|0�W�E2�mCB7�� �d~t%T0 k� �t5�x5"�2't ��1"t'!  ��    � < ��|��;UDH3C��l���|0�W�E2�lCB63��h~t%T0 k� �p4�t4"�2't ��1"t'!  ��    � < ��|��<UDL3EA�k���|0�[�E2�jCB63��l~t%T0 k� �l3�p3"�2't ��1"t'!  $�    � < ��{��=UDL4EA�i���|0�_�E2�gCB54�tt&T0 k� �p3�t3"�2't ��1"t'!  ��    � < ��{��>E�P5EA�h���|0�_�E2�fCB44�xt'T0 k� �t3�x3"�2't ��1"t'!  ��    � < ��{��?E�P5EA�g���|0�c�E"�dCB44�|t'T0 k� �t3�x3"�2't ��1"t'!  ��    � < ��{��@E�P6E1�f���|0�g�E"�cCB34��t'T0 k� �x3�|3"�2't ��1"t'!  ��    � < ��z��AE�P7E1�d���|0�k�E"�_CB24���t(T0 k� �|3��3"�2't ��1"t'!  ��    � < ��z��BE�P7E1�c���|0�o�E"�^CR1$����(T0 k� ��3��3"�2't ��1"t'!  ��    � < �z��CE�P8E1�b���|0�s�E"�\CR0$��� )T0 k� ��3��3"�2't ��1"t'!  ��    � < �z��DE�L8CA�a���|0�w�E"�ZCR/$��� )T0 k� ��3��3"�2't ��1"t'!  ��    � < �y�EE�L9CA�^���|0��E"�WCR-$����)T0 k� ��3��3"�2't ��1"t'!  ��    � < �y�FE�L:CA�]���|0���E"�UCR,$а~��*T0 k� ��3��3"�2't ��1"t'!  ��    � < ��yGE�H:CA�[���|0���E"�SCR*$д~��*T0 k� ��3��3"�2't ��1"t'!  ��    � < ��x HE�H:CA�Z���|0���E"�QCR)$м~��*T0 k� ��3��3"�2't ��1"t'!  ��    � < ��x(HE�H;CA�Y���|0���E"�OIR($ ��~��*T0 k� ��3��3"�2't ��1"t'!  ��    � < ��x0IE�H;CA�W���|0�E�MIR'$ ��}��*T0 k� ��3��3"�2't ��1"t'!  ��    � < ��w@JE�H;CA�T���|0£�E�JIR%$ ��}��*T0 k� ��3��3"�2't ��1"t'!  ��    � < � wHKE�H<CQ�R���|0§�E�HIR$(!��}��*T0 k� ��3��3"�2't ��1"t'!  ��    � < �wPLE�H<CQ�Q���|0¯�E�FIR#,"��|��*T0 k� ��3��3"�2't ��1"t'!  ��    � < �wXLAH<CQ�O���|0³�B��DIb"0#��|��*T0 k� ��3��3"�2't ��1"t'!  ��    � < �w`MAH<CQ�N���|0»�B� CIb!0$��|��*T0 k� ��3��3"�2't ��1"t'!  ��    � < �whNAH<CQ�M���!�0�×B�AIb �4%��|��*T0 k� ��3��3"�2't ��1"t'!  ��    � < �v�pNAH<IQ�K���!�0�ǗB�?Ib�8&�|��)T0 k� ��3��3"�2't ��1"t'!  ��    � < �v�tOAH<IQ�J���!�0�ϗB�>Ib�<&�{��)T0 k� ��3��3"�2't ��1"t'!  ��    � < � w�|OC4H:IQ�I���!�0�חE<IR�<'�{��(T0 k� ��3��3"�2't ��1"t'!  ��    � < �(w��PC4H9IQ�H���!�0�ۗE:IR�@(�{��(T0 k� ��3��3"�2't ��1"t'!  ��    � < �,w��PC4H9IQ�G���!�0��E 9IR�D(�${��'T0 k� ��0��0"�2't ��1"t'!  �	    � < �8w��QC4H9Ia�E���!�0��E,6IR�D'�4z��&T0 k� ��-��-"�2't ��1"t'!  ��	    � < "<w��QO4H9Ia�D���!�0���I44Ib�H'�8z��&T0 k� ��+��+"�2't ��1"t'!  ��	    � < "@x��QO4H9Ia�C��!�0���I83Ib�H'�@z��%T0 k� ��*��*"�2't ��1"t'!  ��	    � < "Hx��RO4H8Ia�B��!�0	�I@2Ib�H'�Hz��%T0 k� �|)��)"�2't ��1"t'!  ��	 	   � < "Lx��RO4L8Ia�A��|0	�ID0Ib�L'�Pz��$T0 k� �|(��("�2't ��1"t'!  ��	 	   � < "Ty��RO4L8IQ�@��|0	�IH/Ib�L'�Xz��$T0 k� �|(��("�2't ��1"t'!  ��	 	   � < "Xx��RO4L8IQ�?��|0	�IP.IR�L'�`y��#T0 k� �|(��("�2't ��1"t'!  ��	 	   � < "`x��RO4L8IQ�>���|0	#�I#T-IR L'�hy� #T0 k� ��&��&"�2't ��1"t'!  ��	 	   � < dx��RO4L8IQ�>���|0	'�I#X,IR P'�py� #T0 k� ��%��%"�2't ��1"t'!  ��	 	   � < lx��RO4L7IQ�=���|0	#/�I#\+IR P'�ty� #T0 k� ��$��$"�2't ��1"t'!  ��	 	   � < xw��RO4L7E��;���|0	#7�I#d)IR T'�y� "T0 k� ��#��#"�2't ��1"t'!  ��	 	   � < �w� RO4L7E��:���|0	#?�Ih(@�P'�x� "T0 k� ��"��""�2't ��1"t'!  �� 	   � < �w�RO4L7E��9Q��|0	#C�Ih'@�P'�x� !T0 k� �|!��!"�2't ��1"t'!  �� 	   � < �v�RO4L7E��8Q��|0	G�Il&@�P'�x� !T0 k� �t!�x!"�2't ��1"t'!  �� 
   � < �v�QO4L7E��7Q��!�0	K�Ip&@�P&�x�!T0 k� �p �t "�2't ��1"t'!  �� 
   � < �v� QO4L7C�6Q��!�0	O�It%@�P&�x�!T0 k� �h�l"�2't ��1"t'!  �� 
   � < �v�,QO4P7C�5Q��!�0	S�I#t$C�DP&�x� T0 k� �h�l"�2't ��1"t'!  � 
   � < �v�4QO4P7C�4��!�0	W�I#x$C�DP%�x� T0 k� 4h�l"�2't ��1"t'! �� 
   � < �u�<PO4P7C�3��!�0	#[�I#|#C�DL%��w� T0 k� 4d�h"�2't ��1"t'! �� 
   � < �u�DPO4P7C�2��!�0	#_�I#|#C�DL%��w� T0 k� 4d�h"�2't ��1"t'! �� 
   � < ��uLPO4P7EѠ1��!�0	#c�I#�"C�DL$��w� T0 k� 4`�d"�2't ��1"t'! �� 
   � < ��t\OO4P6Eј/���!�0	#g�E�!C�tL#��v� T0 k� �\�`"�2't ��1"t'! �� 
   � < ��tdOO4P6Eј.���!�0	k�E�!C�tL"��v� T0 k� �\�`"�2't ��1"t'! ��    � < ��tlNO4T6Eє.���!�0	k�E� C� tL"��v�T0 k� �X�\"�2't ��1"t'! ��    � < ��shNAT6Eѐ-���|0	o�E� C� tL!��v�T0 k� �X�\"�2't ��1"t'! ��    � < ��shNAT6E�,���|0	s�E�C��tL ��u�T0 k� �T�X"�2't ��1"t'! ��    � < ��rdMAT6E�+���|0	s�E��C��dL�u�T0 k� �T�X"�2't ��1"t'! ��    � < ��rdMAT6E�+���|0	#w�E��C��dH�t�T0 k� �P�T"�2't ��1"t'! ��    � < �q`LAP5E�|)���|0	#w�E��C��dD �t�T0 k� �L�P"�2't ��1"t'! ��    � < �p�`KATP5EQx)��|0	#{�E��C��dD �$s� T0 k� �L�P"�2't ��1"t'! ��    � < �o�`JATP5EQp(��|0	#{�DӨC��TD �,s� T0 k� DH�L"�2't ��1"t'! ��    � < �$o�`JATP4EQl'�{�|0	{�DӬC��TD �0r� T0 k� DH�L"�2't ��1"t'! ��    � < �,n�\IATL4EQh'�{�|0	�DӰC��T@ �8r� T0 k� DD�H"�2't ��1"t'! ��    � < �4m�\HATL4EQ`&�w�|0	�DӴC��T@ �@q��T0 k� DD�H"�2't ��1"t'! ��/    � < �<lt\GEDH4EQ\%�w�|0	�DӼC��T< �Hq��T0 k� D@�D"�2't ��1"t'! ��/    � < �Pkt\FEDD3EQP$�o�|0	�DӼC��T< �Xp��T0 k� $<�@"�2't ��1"t'! ��/    � < �Xjt\EED@2EQL$�o�|0	#�DӼC���< �\o��T0 k� $<�@"�2't ��1"t'! ��/    � < �`it\DED@2C�D#�k�|0	#�E��C��
�< �do��T0 k� $8�<"�2't ��1"t'! ��/    � < �hht\CED<1C�@"�g�|0	#�E��C��	�< �ln��T0 k� $8�<"�2't ��1"t'! ��/    � < �xgt\AED80C�4!�c�|0	#�E�� C���< �|m��T0 k� �4�8"�2't ��1"t'! ��/    � < �ftX@E440C�,!�_�|0 ��E�� C���<�l��T0 k� �0�4"�2't ��1"t'! $�/    � < �edX?E400C�$ �[�|0 ��E��!C���<�l��T0 k� � �$"�2't ��1"t'! ��+    � < �ddX=E400C�  �W�|0 ��Es�!C���<�k3�T0 k� ��"�2't ��1"t'! ��+    � < �bdX=E4(/C��O�|0 ��Es�"C�� �<�j3�T0 k� ��"�2't ��1"t'! ��+    � < �adX<PT$/C��K�|0 ��Es�#C����<�i3�T0 k� ��� "�2't ��1"t'! ��+    � < ��`dX;PT 0C� �C�|0�Es�#C����8�h3�T0 k� #���"�2't ��1"t'! ��+    � < ���`dX:PT0C���?�|0�Es�$C����8�hs�T0 k� #���"�2't ��1"t'! ��+    � < ���^dX8PT0C���7�|0�Es�%C����8��fs�T0 k� #���"�2't ��1"t'! ��+    � < ���]dX7Pd0C���3�|0�Es�&C����8 ��fs�T0 k� #���"�2't ��1"t'! ��+    � < ���\TT6Pd1C���+�|0�Es�'C����8 ��es�T0 k� ����"�2't ��1"t'! ��+    � < ���[TT5Pd1C���'�|0S�Es�(C����8 ��ds�T0 k� ����"�2't ��1"t'! ��+    � < ���ZTT4Pd1C���#�|0S�Ec�)C����8 ��ds�T0 k� ����"�2't ��1"t'! ��+    � < ���XTP2Pd1C���|0S�Ec�)C�w��8!��b��T0 k� ����"�2't ��1"t'! �+    � < �� W�P2PT1C���|0S�Ec�)C�s��8!��a��T0 k� ����"�2't ��1"t'! ��+    � < �tV�P2PT1C���|0��Ec�*C�k��8!�a��T0 k� ����"�2't ��1"t'! ��+    � < �tU�P2PT1C���|0�{�g�+C�g��8! `��T0 k� ���"�2't ��1"t'! ��+    � < �tT�P3PT2D ����|0�{�g�+C�_��8"_��T0 k� #���"�2't ��1"t'! ��+    � < �t$Q�L3PT3D ����|0�w�g�-C�S��8"]��T0 k� #���"�2't ��1"t'!  ��+    � < �t,P�L3E43D |���|0�s�g�-C�O��8"]��T0 k� #���"�2't ��1"t'!  ��+    � < �t4O�H4E43D t���|0�s�g�-C�G��8"�$\��T0 k� #���"�2't ��1"t'!  �+    � ; �tDL�H4E43D d���|0�k�g�.C�;��8"�0Zs�T0 k� ����"�2't ��1"t'! ��/    � : �tHK�H4E43D \���|0Ck�g�.E�7��8"�8Ys�T0 k� ����"�2't ��1"t'! ��/    � 9 �tPI�H4@�3D T���|0Cg�g�/E�/��8"�@Xs�T0 k� �|	��	"�2't ��1"t'! ��/    � 8 �tXH�H4@�3D L ��|0Cc�g�/E�+�
�8"�DXs�T0 k� �t�x"�2't ��1"t'! ��/    � 7 �d\G�H4@�2D D ��|0C_�g�0E�#�
�8"�LWs�T0 k� �h�l"�2't ��1"t'! ��/    � 6 �dlD�H4@�2D4 ��|0CW�g#�1E��
�<"�XUs�T0 k� �T�X"�2't ��1"t'! ��/    � 5 �dpB�H4@d2D( ��|0CS�g#�1E��
�<"�`T��T0 k� #L �P "�2't ��1"t'! ��/    � 4 �dtA�H4@d2D 	���|03O�g#�2E���<"�hS��T0 k� #C��G�"�2't ��1"t'! ��/    � 3 �d|?�H4@d1D	���|03O�g#�2E���<"slR��T0 k� #7��;�"�2't ��1"t'! ��/    � 2 �d�<�H3@d1D	���|03G�g#�3E����<"s|P��T0 k� ##��'�"�2't ��1"t'! ��/    � 0 �d�;�H3B�0D 	���|03C�g#�4E����<"s�O��T0 k� ����"�2't ��1"t'!	 ��/    � . �d�9�H2B�0D�	��|03?�g#�4E����8"s�N��T0 k� ����"�2't ��1"t'!	 ��/    � , �d�7�H2B�/K�	�w�|0�;�g�5E����8"s�M��T0 k� ����"�2't ��1"t'!	 ��/   � * �d�4dH2B�/K�	�o�|0�3�g�6E����4"s�K��T0 k� ������"�2't ��1"t'!
 ��/    � ( �d�2dH2E�.K�	�g�|0�/�g�6E����4!s�Js�T0 k� ������"�2't ��1"t'!
 ��/    � & �T�1dH2E�.K�	�c�|0�+�g�6E����0!s�Is�T0 k� ������"�2't ��1"t'! ��/    � $ �T�/dH2E�.E�	�_�|0�'�g�7E����0!s�Gs�T0 k� ������"�2't ��1"t'! ��/    � " �T�-dD2E�-E�	�[�|0�#�g�7E����, s�Gs�T0 k� "�����"�2't ��1"t'! ��/    �   �T�*TD1E�-E�	�S�|0��g�6Eг��(s�Fs�T0 k� "�����"�2't ��1"t'! ��/    �  ~T�)T@1E� -E�
	�O�|0��g�6C௿�(c�Fs�T0 k� "�����"�2't ��1"t'! ��/    �  zT�'T@1E� ,E�
	�K�|0��g�6C৾�(c�Es�T0 k� "�����"�2't ��1"t'! ��/    �  vT�&T<0E��,E�		�G�|0��g�5C����(c�Es�T0 k� ������"�2't ��1"t'! ��/    �  rT�$T<0E��,E�	�C�|0��g�5C����$c�Ds�T0 k� ������"�2't ��1"t'! ��/    �  nT�!T40E��+E��	�?�|0���g�4C���� c�Cs�T0 k� �w��{�"�2't ��1"t'! ��/    �  jT| �4/E��*E�|	�;�|0��D3�4C���� 3�Bs�T0 k� �o��s�"�2't ��1"t'! ��/    �  fTx�0/E��*E�t	�7�|0��D3�3C��3�As�T0 k� �c��g�"�2't ��1"t'! ��/   �  bDt�,/E��*E�l	�7�|0��D3�3C�w�3�@s�T0 k� �[��_�"�2't ��1"t'! ��/    �  ^Dp�(/E��)E�h	�3�|0�ߪD3�3E@o�3�@s�T0 k� "O��S�"�2't ��1"t'! ��/    �  ZDl�$/E��)E�`	�/�|0�۪D3�3E@g�3�?s�T0 k� "C��G�"�2't ��1"t'! ��/    � 
 VDh� .E��(E�X 	�/�|0�ӫEc�3E@_�3�>3�T0 k� ";��?�"�2't ��1"t'! ��O    �  SDd�.E��(E�S�	�+�|0�ˬEc�3E@[�3�=3�T0 k� "/��3�"�2't ��1"t'! ��O    �  P�\�.C��'E�C�	�'�|0⿭Ec�3E@K�3�=3�T0 k� ����"�2't ��1"t'!
 ��O    �  L�X�.C��'E�;�	�'�|0ⷮEc�3E@C� 3�=3�T0 k� ����"�2't ��1"t'!
 ��O    �  I�T�-C��&E�7��#�|0⯯ES�3E@;��3�=3�T0 k� ����"�2't ��1"t'!
 ��O    �   F�P�-C�&E/���|0⧯ES�3E@7��3�<3�T0 k� �����"�2't ��1"t'!	 ��O    ��� C�L�,C�&E'���|0⟰ES�3E@/��C�<3�T0 k� �����"�2't ��1"t'!	 ��O    ��� @�L�,C�%E���|0⛱ES�3C�'��C�;3�
T0 k� ����"�2't ��1"t'!	 ��O    ��� =�H�+C�%E���|0⓱ES�3C���C�;3�
T0 k� �߼��"�2't ��1"t'! ��O    ��� :�H� *C�%E���|0⋲C�|3C���C�:3�	T0 k� !׺�ۺ"�2't ��1"t'! ��O    ��� 7�D��*C�$E���|0��C�x3C���C�:3�T0 k� !˸�ϸ"�2't ��1"t'! ��O    ��� 4�@��*C�$E����|0�o�C�p3C����C�93�T0 k� !�����"�2't ��1"t'! ��O    ��� 1�<c�)C�#J����|0�g�C�h3C�����C�93�T0 k� !�����"�2't ��1"t'! ��O    ��� .�<c�(C�#J��?��|0�_�C�d3C�����C�83�T0 k� ������"�2't ��1"t'! ��O    ��� +�8c�(C�x#J��?��|0�W�C�`3C�����83�T0 k� ������"�2't ��1"t'! ��O    ��� (�4c�'C�p#J��?��|0�O�C�X3C�����7c�T0 k� ������"�2't ��1"t'! ��O    ��� %�4c�&C�h"J��?��|0�G�C�T3C��3���7c�T0 k� ������"�2't ��1"t'! ��O    ��� "�0��%C�`"J��?��|0�?�C�L3C�ۛ3���6c�T0 k� �{���"�2't ��1"t'! ��O    ��� �0��%C�X"J�����|0�7�C�H3EOӚ3���5c�T0 k� �o��s�"�2't ��1"t'! ��O    ��� �,��$C�P!J�����|0�/�C�@3EO˘3���5c� T0 k� �g��k�"�2't ��1"t'! ��O    ��� �, ��#C�H!E�����|0'�C�83EOǗ3���4c� T0 k� �[��_�"�2't ��1"t'! ��O    ��� �(!��#D@!E�����|0�C�43EO�����3c��T0 k� !S��W�"�2't ��1"t'!  ��O    ��� �$"��"D8 E�����|0�C�,3EO�����2c��T0 k� !G��K�"�2't ��1"t'!  ,�O    ��� �$#��!D0 E�����|0�C�$3EO�����2c��T0 k� !;��?�"�2't ��1"t'!  ��O    ��� � $��!D( E�����|0�C�3EO���|��1c��T0 k� !3��7�"�2't ��1"t'!  ��O    ��� 
�%�� D  E�����|0��C�3EO���t��1c��T0 k� !'��+�"�2't ��1"t'! ��O    ��� �&��DE�����|0��C�3EO���l��0c��T0 k� ���#�"�2't ��1"t'! ��O    ��� �'��DE{����|0�C�3P���d�/c��T0 k� ����"�2't ��1"t'! ��O    ��� �)��DEs����|0�D 3P���`
�/c��T0 k� ����"�2't ��1"t'! ��O    ������*��D�Ek����|0߾D�3P���X�.c��T0 k� �����"�2't ��1"t'! ��O    ������+��D�E.c����|0׾D�3P���P�-c��T0 k� ������"�2't ��1"t'! ��O    ������,��D�E.[����|0ϿD�3P{��L�-c��T0 k� ����"�2't ��1"t'! ��O    ������-��D�E.S����|0ǿD�3Pw��D�,c��T0 k� ����"�2't ��1"t'! ��O    ������ .ӼD�E.K����|0��D�3P�o��<�,c��T0 k�  ׊�ۊ"�2't ��1"t'! ��O    �������/ӼD�E.C����|0��D�3P�k��8�+c��T0 k�  ω�Ӊ"�2't ��1"t'! ��O    �������0ӸD�E.;����|0��D�3P�c��0 �+c��T0 k�  Ç�Ǉ"�2't ��1"t'! ��O    �������1ӴD�E.3����|0��D�3P�_��/��*c��T0 k�  �����"�2't ��1"t'! ��O    �������2ӴD�E.+����|0��D�3P�W��'��*c��T0 k�  �����"�2't ��1"t'! ��O    �������3ӰD�E#����|0��D�3P�S��#��)c��T0 k� ������"�2't ��1"t'! ��O    �������4ӰD�E����|0��D�3P�O���)c��T0 k� ����"�2't ��1"t'! ��O    �������5ӬD�E����|0��D�3P�G���(c��T0 k� ��}��}"�2't ��1"t'! *�O    �������6ӬD�E����|0{�D�3P�C���(c��T0 k� ��~��~"�2't ��1"t'! ��O    �������7ӨD�E����|0�s�D�3P?���'c��T0 k� �~��~"�2't ��1"t'! ��O    �������8ӨC�|B�����|0�k�D|3P7���'c��T0 k� 0s�w"�2't ��1"t'! ��O    �������9ӤC�tB����{�|0�c�Dp3P3���&c��T0 k� 0k�o"�2't ��1"t'! ��O    �������:ӤC�lB����w�|0�[�Dh3P/����&c��T0 k� 0_��c�"�2't ��1"t'! ��O    ������:ӠC�`B����w�|0�S�D`3P'����%c��T0 k� 0W��[�"�2't ��1"t'! ��O    ������;ӠC�XB���s�|0�G�DT3EO#����%c��T0 k� 0K��O�"�2't ��1"t'!  ��O    ������<ӠEBPE���o�|0�?�DL3EO�����$c��T0 k�  C��G�"�2't ��1"t'!  ��O    ������=ӜEBHE���k�|0�7�DD3EO�����$c��T0 k�  ;��?�"�2't ��1"t'!  ��O    ������>ӜEB@E���g�|0�/�C�83EO�����#c��T0 k�  /��3�"�2't ��1"t'!  .�O    ������?ӘEB4E���c�|0�'�C�03EO�����#c��T0 k�  '��+�"�2't ��1"t'!  ��O    ������?ӘEB,E���c�|0��C�(3E?�����#c��T0 k�  ���"�2't ��1"t'!  ��O    ������@ӔEB$E���_�|0��C�3E?�����"c��T0 k� ����"�2't ��1"t'!  ��O    ������AӔEBE���[�|0��C�3E?����"3��T0 k� ����"�2't ��1"t'!  ��O    ������|BӔEBE���W�|0��C�3E>�����!3��T0 k� �����"�2't ��1"t'!  ��O    ������tBӐEBE���oW�|0���C� 3E>�����!3��T0 k� ������"�2't ��1"t'!  ��O    ������lC�C� E���oS�|0���C��3E.����3� 3��T0 k� ����"�2't ��1"t'!  ��O    ������dD�C��E��oO�|0���C��3E.���3� 3��T0 k� ����"�2't ��1"t'!  ��O    ������\E�C��E��oK�|0���C��3E.���3| 3��T0 k� �׆�ۆ"�2't ��1"t'!  ��O    ������TE�C��E��oG�|0���C��3E.���3|3��T0 k� �χ�Ӈ"�2't ��1"t'!  ��O    �����LF�C��E��/?�|0���C��3E.���3x3��T0 k� �Ǉ�ˇ"�2't ��1"t'!  ��O    �����DG�E��E��/7�|0���C��3E.���3t3��T0 k� ������"�2't ��1"t'!  ��O    �����<G�E��E��//�|0���C��3E.���3t3��T0 k� ������"�2't ��1"t'!  ��O    �����4H�|E��E��/'��0л�C�3E.ߌ����p3��T0 k� ������"�2't ��1"t'!  ��O    �����,I�|EѸE��/��0г�C�3Eی����p3��T0 k� ������"�2't ��1"t'!  ��O    ����� I�xEѰE��/��0 Ы�C�3Eۋ����l3��T0 k� ������"�2't ��1"t'!  ��O    �����J�tEѨE��/��3�У�C�3Eۊ����l3��T0 k� ������"�2't ��1"t'!  �O    �����J�p
EѠE���/��3�Л�C�3E׊����h3��T0 k� ������"�2't ��1"t'!  ��O    �����K�p	C�E���/��3�Г�C�3E׉���sh3��T0 k� �{���"�2't ��1"t'!  ��O    ����� LSlC�E���.���3�Ї�C�3B�ۉ���sd3��T0 k� �o��s�"�2't ��1"t'!  ��O    ������LShC�E���.���3���C�x3B�����s`3��T0 k� �g��k�"�2't ��1"t'!  ��O    ������MSdC�|E���.��3��w�C�l3B����s\3��T0 k� �_��c�"�2't ��1"t'!  ��O    ������MSdC�tE���.��3��o�Dd3B����s\3��T0 k� �S��W�"�2't ��1"t'!  ��O    ������NS`C�hE���.��3��g�D\3B����sX3��T0 k� �K��O�"�2't ��1"t'!  ��O    ������NS`C�`E���.ۘ�3��_�DP3B�����sT3��T0 k� �;��?�"�2't ��1"t'!  ��H    ������Oc\C�XE���.ו�3��W�DH3B�����sP3��T0 k� �;��?�"�2't ��1"t'!  ��H    ������PcX C�PE���.ϓ�3��O�D@3B�����sP3��T0 k� �;��?�"�2't ��1"t'!  ��H    ������Pc[�C�HE��.ˑ�3��C�D43B����sL3��T0 k� �;��?�"�2't ��1"t'!  ��H    ������QcW�C�<E��.Ï�3��;�E�,3B����sH3��T0 k� �?��C�"�2't ��1"t'!  ��H    ������QcS�C�4E��.���3��3�E�$3B�����sH3��T0 k� �C��G�"�2't ��1"t'!  ��H    ������RcS�C�,E��.���3�0+�E�3B�����sD3��T0 k� �G��K�"�2't ��1"t'!  ��H    ������RcO�C�$E��.���3�0#�E�3B�����s@3��T0 k� �K��O�"�2't ��1"t'!  ��H    ������SsO�C�E��.���3�0�E�3B����s@3��T0 k� �O��S�"�2't ��1"t'!  ��H    ������SsK�C�E��.���3�0�E� 4B����s<3��T0 k� �S��W�"�2't ��1"t'!  ��H   ������TsK�C�E��.���3�0�E��4B�#���s8
3��T0 k� �W�["�2't ��1"t'!  ��H    ������tTsG�EA E��.���3�0�E��4B�+���s8	3��T0 k� �[�_"�2't ��1"t'!  ��H    ������lTsG�E@�E��	����3�?��E��4B�/���s43��T0 k� �_�c"�2't ��1"t'!  ��H    ������dUsC�E@�E��	����3�?��E��5B�3���s43��T0 k� �g�k"�2't ��1"t'!  ��H    ������\UsC�E@�
E��	����3�?��D0�5B�7���s03��T0 k� �k�o"�2't ��1"t'!  ��H    ������TVs?�E@�
E�	����3�?��D0�5B�;��#�s,3��T0 k� �o��s�"�2't ��1"t'!  ��H    ������LVs?�E@�	E��	����3�?��D0�6B�?��+�s,3��T0 k� �s��w�"�2't ��1"t'!  ��H    ������@Ws;�E@�	E��	���3�?��D0�6B�C��/�s(3��T0 k� �w��{�"�2't ��1"t'!  ��H    ������8Ws;�C��E��	�{��3�O��D0�7B�G��3�s(3��T0 k� �{���"�2't ��1"t'!  ��H    ������0Ws7�C��E��	�w��3�O��D0�7B�G��;��$3��T0 k� �{���"�2't ��1"t'!  ��H    ������(Xs7�C��E���	�s��3�O��D0�8B�K��?��$3��T0 k� �����"�2't ��1"t'!  �H    ������ Xs3�C��F��	�s��3�O��A��8EO��C��  3��T0 k� �{���"�2't ��1"t'!  �H    ������Ys3�C��F��	�o��3�O��A��9ES��K��#�3��T0 k� �w��{�"�2't ��1"t'!  ��H    ������Ys/�E@�F�	�k��3����A��9EW� cO���3��T0 k� �w��{�"�2't ��1"t'!  ��H    ������Ys/�E@�F�	�k��3����A�x:E_� cS���3��T0 k� �w��{�"�2't ��1"t'!  ��H    �������Zs+�E@�F�	�g��3����A�l:Ec� c[���3��T0 k� �w��{�"�2't ��1"t'!  ��H    �������Zs+�E@|E��	�c��3����A�d:E�g� c_���3��T0 k� �{���"�2't ��1"t'!  ��H    �������[s+�E@tE��	�c��3���A�\;E�k� cc���3��T0 k� �����"�2't ��1"t'!  ��H    �������[s'�E@lE��	�_��3��{�A�T;E�o� cg���3��T0 k� ������"�2't ��1"t'!  ��H    �������[s'�E@dE�#�	�_��3��s�A�L<E�w� ck���3��T0 k� ������"�2't ��1"t'!  ��H    �������\s#�E@\ E�'�	�_��3��k�A�D<E�{� cs���3��T0 k� ������"�2't ��1"t'!  ��H    �������\s#�C�W�E�+�	�[��3��c�A�@=E�� cw���3��T0 k� ������"�2't ��1"t'!  ��H    �������\s#�C�K�E�3�	�[��3��_�A�8=E��� c{���3��T0 k� ������"�2't ��1"t'!  ��H    ������\s�C�C�E�7�	�[��3��W�A�0=E��� c���3��T0 k� ������"�2't ��1"t'!  ��H    ������]s�C�;�E�?�	�[��3��O�A�(>E��� c����3��T0 k� ������"�2't ��1"t'!  ��H    ������]s�C�3�E�C�	�[��3��K�A� >E�� c����3��T0 k� ������"�2't ��1"t'!  ��H    ������]s�C�+�E�K�	�W��3��C�A�?E�� c����3��T0 k� ������"�2't ��1"t'!  ��H    ������]s�C�#�E�O�	�W��3��?�A�?E�� c����3��T0 k� ������"�2't ��1"t'!  ��H    ������]s�C��E�W��W��3��7�A�?E�� c����3��T0 k� ������"�2't ��1"t'!  ��H    ������]s�C��E�_��W��3��3�A�@E�� c����3��T0 k� ������"�2't ��1"t'!  ��H    ������x]s�C��E�c��W��3��+�A� @E�� c����3��T0 k� ������"�2't ��1"t'!  ��H    �����1p]s�C��E�k��W��3��'�A��AE�� c����3��T0 k� �ã�ǣ"�2't ��1"t'!  ��H    �����1d\s�C���E�o��W��3���A��AE�� c����3��T0 k� �Ǥ�ˤ"�2't ��1"t'!  ��H    �����1\\s�C���E�w� W��3���A��AE�� c�����3��T0 k� �˥�ϥ"�2't ��1"t'!  ��H    �����1T\s�C���E�� [��3���A��BEÐ c�����3��T0 k� ������"�2't ��1"t'!  �H    �����1L\s�C���E��� [��3���A��BH�Ǒ c�����3��T0 k� ������"�2't ��1"t'!  ��O    �����1@\s�C���E��� [��3���A��BH�˒ c�����3��T0 k� ������"�2't ��1"t'!  ��O    �����18[s�C���E��� [��3���A��CH�ϓ c�����3��T0 k� ������"�2't ��1"t'!  ��O    �����10[s�C���E����_��3����A��CH�Ӕ c�����3��T0 k� �����"�2't ��1"t'!  ��O    �����1([s�C���E����_��3����A��CH�ו c�����3��T0 k� �o��s�"�2't ��1"t'!  ��O    �����1 Zs�C���E����_��3���A��DH�ߖ cË���3��T0 k� �_��c�"�2't ��1"t'!  ��O    �����1Zs�C���E����c��3���A��DH� cǋ���3��T0 k� �S��W�"�2't ��1"t'!  ��O    �����1Zs�C���E����c��3���A��DH� cǊ���3��T0 k� �C��G�"�2't ��1"t'!  ��O    �����AYs�C���E����c��3���A��EH� cˊ���3��T0 k� �3��7�"�2't ��1"t'!  ��O    �����@�Ys�C���E����g��3���A��EH� cω���3��T0 k� �#��'�"�2't ��1"t'!  ��O    �����@�Xs�C���E�ì�g��3��ۻA��EH� cӉ���3��T0 k� ����"�2't ��1"t'!  ��O    �����@�Xs�C���E�ǫ�g��3��׻A��EHo�� c׈���3��T0 k� ����"�2't ��1"t'!  ��O    �����@�Ws�C���E�Ϫ�k��3��ӻA��FHo�� c׈���3��T0 k� ������"�2't ��1"t'!  ��O    �����@�Ws�C�{�E�өNk��3��ϻA��FHo�� cۇ���3��T0 k� ����"�2't ��1"t'!  ��O    �����@�Vr��C�s�E�רNk��3��˺A��FHo�� c߇���3��T0 k� �ۭ�߭"�2't ��1"t'!  ��O    �����@�Vr��C�k�E�ۦNo��3��ǺA��GH`� c����3��T0 k� �ï�ǯ"�2't ��1"t'!  ��F    �����@�Ur��C�c�E�ߥNo��3�^úA��GH`� c����3��T0 k� ������"�2't ��1"t'!  ��F    �����@�Tr��C�[�E��No��3�^��A��GH`� c����3��T0 k� ������"�2't ��1"t'!  ��F   �����@�Tr��C�S�E���s��3�^��A��GH`� c����3��T0 k� ������"�2't ��1"t'!  ��F    �����P�Sr��C�K�E���s��3�^��A�|HH`� c����3��T0 k� ������"�2't ��1"t'!  ��F    �����P�Sr��C�C�E���s��3�^��A�tHH`� c����3��T0 k� ������"�2't ��1"t'!  ��F    �����P�Rr��C�;�E���s��3�^��A�pHH`� c����3��T0 k� ������"�2't ��1"t'!  ��F    �����P�Qr��C�3�E����w��3�^��A�lHH`� c�����3��T0 k� ������"�2't ��1"t'!  ��F    �����P�Pr��C�+�E����w��3�^��A�hIH`� c�����3��T0 k� ������"�2't ��1"t'!  ��F    �����P|Pr��C�#�E����w��3�^��A�dIH`#� c�����3��T0 k� �{���"�2't ��1"t'!  ��F    �����PtOr��EO�E����{��3�^��A�`IH`'� c�����3��T0 k� �w��{�"�2't ��1"t'!  ��F    �����PlNr��EO�E����{��3�N��A�\IH`+� c�����3��T0 k� �o��s�"�2't ��1"t'!  ��F    �����PdMr��EO�E���{��3�N��A�XIH`+� c�����3��T0 k� �k��o�"�2't ��1"t'!  ��F    �����P\Mr��EO�E���{��3�N�A�TJH`/� c�����3��T0 k� �c��g�"�2't ��1"t'!  ��F    �����PTLr��EN��E�����3�Nw�A�PJH`3� c�����3��T0 k� �_��c�"�2't ��1"t'!  ��F    �����`HKr��EN��E�����3�Ns�A�LJH`7� c�����3��T0 k� �W��[�"�2't ��1"t'!  ��F    �����`@Jr��EN��E�����3��k�A�HJH`7� d����3��T0 k� �O��S�"�2't ��1"t'!  ��F    �����`8Ir��EN��E�����3��c�A�DKA�;� d����3��T0 k� �G��K�"�2't ��1"t'!  ��F    �����`0Ir��E>��E�����3��_�A�@KA�?� d����3��T0 k� �?��C�"�2't ��1"t'!  ��F    �����`(Hr��E>��E���3��W�A�<KA�?� d����3��T0 k� �7��;�"�2't ��1"t'!  ��F    �����` Gr��E>��E���3��O�A�<KA�C� d����3��T0 k� �/��3�"�2't ��1"t'!  ��F    ������Fr��E>��E���3��G�A�8KA�G� d����3��T0 k� �'��+�"�2't ��1"t'!  ��F    ������Er��E>��E���3��?�A�4LA�G� d����3��T0 k� ���#�"�2't ��1"t'!  ��F    ������Dr��E>��D?��3��;�A�0LA�K� d����3��T0 k� ����"�2't ��1"t'!  ��F    ������ Cr��E>��D?��3�n3�A�,LA�O� d����3��T0 k� ����"�2't ��1"t'!  ��F    �������Br��E>��D?��3�n+�A�(LA�O� d����3��T0 k� �����"�2't ��1"t'!  ��F    �������Ar��E>��D?�#,3�n#�A�(LA�S� d����3��T0 k� ����"�2't ��1"t'!  ��F   �������@r��E>��D?�#,3�n�A�$MA�S� d����3��T0 k� �׵�۵"�2't ��1"t'!  ��F    �������?r��Lޛ�D>��#,3�n�A� MA�W� d����3��T0 k� �˵�ϵ"�2't ��1"t'!  ��F    �������>r��Lޗ�D>��#,3�N�A�MA�[� d����3��T0 k� �˺�Ϻ"�2't ��1"t'!  ��F    �������=r��Lޏ�D>��#,3�N�A�MA�[� d����3��T0 k� �˽�Ͻ"�2't ��1"t'!  ��F    �������<r��Lދ�D>��#,3�M��A�MA�_� d����3��T0 k� ������"�2't ��1"t'!  ��F    �������;r��Lރ�D>��#,3�M�A�MA�_� d����3��T0 k� ������"�2't ��1"t'!  ��F    �������:r��L��E���#,3�M�A�NA�c� d����3��T0 k� ������"�2't ��1"t'!  ��F    �������9r��L��E���#,3�M߸A�NA�c� d����3��T0 k� ������"�2't ��1"t'!  ��F    �������8r��L�{�E��#,3�M׸A�NA�g� d����3��T0 k� ������"�2't ��1"t'!  ��F    �������7r��L�s�E��#,3�MϹA�NA�g� d����3��T0 k� ������"�2't ��1"t'!  ��F    �������5r��L�o�E���3�ǹA�NA�k� d����3��T0 k� ������"�2't ��1"t'!  ��F    �������4r��L�k�E���3���A�NA�k� d����3��T0 k� ������"�2't ��1"t'!  ��F    �������3r��L�c�E���3���A� NA�o� d����3��T0 k� ������"�2't ��1"t'!  ��F    �������1r��L�_�E���3���A� OA�o� d����3��T0 k� �w��{�"�2't ��1"t'!  ��F    �������0r��L�W�E���3���A��OA�s� d����3��T0 k� �o��s�"�2't ��1"t'!  ��F   ������|.r��L�S�E���3���A��OA�s� d����3��T0 k� �g��k�"�2't ��1"t'!  ��F    ������t-r��L�O�D���3���A��OA�w� d����3��T0 k� �_��c�"�2't ��1"t'!  ��F    ������p+r��L�G�D�߈�3���A��OA�w� d����3��T0 k� �W��[�"�2't ��1"t'!  ��F    ������h*r��L�C�D�ۈ�3���A��OA�{� d����"s��T0 k� �O��S�"�2't ��1"t'!  ��F    ������d(r��L�?�D�ۉ�3�M�A��OA�{� d����"s��T0 k� �O��S�"�2't ��1"t'!  ��F    ������\'r��L�7�D�׉�3�Mw�A��PA�� d����"s��T0 k� �K��O�"�2't ��1"t'!  ��F    ������X%r��L�3�D�׊#3�Mo�A��PA�� d����"s��T0 k� �G��K�"�2't ��1"t'!  ��F    �����                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��(� ]�#�#� � ����9m   Y Y      �����    ��z����     �	�              J�����          �p�     ���  @
	"         ���   @ V
      � �&�    ��" �{�    �F�   
           N����         ���    ���   8
(         ���'  X X
     ����    ������:�    	   	          ����         I`b      ���  

'          ��I�        ����    ��I�����           
            L	����          ��     ���   8	
	          ��k�   � �	   .���    ��VP�� �    A �              _ ����          %@�    ���   X
	         ����  ��
      B��    ������                               �\              Q  ���    0 0            ���\   x	    V���    ��� ��`�    ����              ����         ��     ��J   8

�          W��   
    j��w     W������     x��               i 6         �     ��@   0

           �Ϯ�       ~ 6��    �Ϛ� 6}�    ,K              �;          �0  �  ��@   (
"
          ���?   ?       �'    ���:v     � �               �� �         	 �     ��@   H	w         ��z,   C      � �HL    ��}� �O4    ����                  �         
 �     ��@   (
         ��X ��     � ��|    ��X ��|                              ���v             �  ��@    0

 2                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         ���  ��        ��K��  ����P��KY�  ���}	                   x                j  �   �   �                         ��    ��        ��L      ��  �L           "                                                 �                         �� ������������ 6 � ����K�L     	    
        
  q  	� �P�G       AD �`� BD  a� B� b  �D  f� ��  f� �  g  �D g` �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0� ���� � � }`���� ����� � Ǥ x@ ��  x` �� @c@ �$ c� �D  c� �� d  �� 0d@ �  d� �D d� -� �`� .� a� .�  a� �D �[� �D \� �d  \� ɤ  ]  �� ]` �� 0}` �$ }����� � ��  z� 
�\ V� 
�� V� 
�\ W  
�\ W� 
�\ W� 
�\ W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ������������ Y  ������  
�fD
��L���"����D" � j  "  B   J jF�"     "�j  " ��
��
��"     
�j
�� 
  
 �
� �  �  
� ��    ��     ��6  �   ����  ��     ���      ��    ��     ���          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �O��      ��! �  ���        �T ��        �        ��        �        ��        �   �    �o	 ��        ��                         ��  0 �� ��                                    �                ����            ������%��  ������               22 Christan Ruuttu     4:48                                                                        2  2     �C
� �E �D � �B� � �K � �K � � K � �K � � 	K" � �
C. � �C1 � � C4 � �C5 � �C7 � Jk~ _ k� �"� � � "� � �"� � �*� � � "K � � "I �7 "& �? ", |": �/ "P �? !� �? !� �/  "G �/ "K �?  "B �?  "B �W  " |{"
� � #"E � �$* | �%!� |&"8 �/ '"E �/  "G �? !� �? !� � � +"& | �,"* | �-"2 | ."@ |/": �/ 0"P �? !� �/ 2"E �/  "G �
  *A� 5*Gx  *Ax  7*Ov  *Kv  *J�.  *E|K ;*Jw[ )�g=**} >*<e( *2u                                                                                                                                                                                                                         `� R @           @ 
      4 	�     a P E b  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    �;�   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, )   c�� �� ��������                                                                                                                                                                                                                                                                                                                                             �"                                                                                                                                                                                                                                         U    0     ��  4�J      -�                             ������������������������������������������������������                                                                                                                                 	       �  ��              �          ��               	 
     �������  ��� ���������������� �������������������� ������� ����� ���� ���� ����������� ����� ���������������������������� ����������������� ������������������������������������� �������� �� ��  �� ������������� ��� ���������������������                                  +         .�J      d�                             ������������������������������������������������������                                                                                                                                          y  ��               �        �    �           	     � ��� ��� ����� ������������������� ����������������� � ��� ����� ������  ������� �� ��������� ��� �������� ��� � ��������������������� �� ����������������������������� ��� �� � �������  ���� �� �� ����������� ������� ����������������            �                                                                                                                                                                                                                             
                     	                                                           �             


           �   }�                                              '�                 +                        ��������  '}  '���������������������������������    ����������������������������  '}���������������������ww�ww333wwwwwwww�ww�ww�ww�ww333wwww E B 6                                 � �� �\        �U�!&R�1U1'                                                                                                                                                                                                                                                           	n1n  
1�        m      b      m      a                        m                                                                                                                                                                                                                                                                                                                                                                                                            C  � (��  � ��  � @��  � #��  EZm4  �N ������������
���������������������o�����ln                �`�? :�A��          �   & AG� �   �   
              �                                                                                                                                                                                                                                                                                                                                      p N K   �     p   $             !��                                                                                                                                                                                                                            Y   �� �~ ���      �� 8      �������  ��� ���������������� �������������������� ������� ����� ���� ���� ����������� ����� ���������������������������� ����������������� ������������������������������������� �������� �� ��  �� ������������� ��� ���������������������� ��� ��� ����� ������������������� ����������������� � ��� ����� ������  ������� �� ��������� ��� �������� ��� � ��������������������� �� ����������������������������� ��� �� � �������  ���� �� �� ����������� ������� ����������������             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    B      4   � ��                       8     �  ���������J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �f ��     �f �$ ^$ �@       �       �     �   n 
� �     �f ��        p����      � �N     `d     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h  y���  ��  y���  �$ ^$    y                      ��� �� � ��� �� � ��� �$  � �  ��  a      �  ��   ?���� e����� g���        f ^�         �� ���      ?      ��)X���2�������J��X����      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                          �      �  a r!   f�"""""*��**"*�"�""�""v""*f   "  ""- ��"�"*"-""z"""""����            n   �  "  q  ��                          �  �                                 � gv"!g�vg�vggfvv|�b��r""gb"�vr�rgb��v���g���v���***�*q!q�"!a�!vwfqqr~� qw��q�~~q�����~~~�w~~w�w            �   ~   ��  ~~  �w      v    �                ggj�vvggvvgg!vg�g֪vvg�r�r��⢪rq**gjb�v�q*gjj*vv��gg�z�/�"!�"�*�""*z����qw�~q~ww��q~qwvq�w�`� ��� �w �~p w�p  ��                    �                        lggz�v��g        �       ggbvvrgggavvvqggav� �      ���w!z�w"""�!""*�"! ��        q� q�        `               �        �                      wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "! " ""                "  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                              """ "!   " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "! " ""                "  !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                              
      �  �  ��  �� �� �� 	�� D� EH EZ  DZ 4J 34Z3EH�T��ʄ
����ܩ���� ""�""�""�"/� �� �  ��� ̽� ��� �w� ��� ��� ��� ˻���ܚ��ة��ی����˻ݼˍ�ۻ���Ѕ" �" R�  B      ��  ��  �     �            � �� �   �       �   ��  ��  ��  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                      "  .���"    �     �                                       �   ���                            �   �                                                                                                                               �   �   �  �  �  �  ���������  �U4"+�B�*�����"/���  ��� �� �  � �     �               ۲  �!  "  �� �� �  ��� ��  �� �                          	ʐ ��� ��� ڝ��ݩ��ݩ��ݩ��ک�̪��̪��̪������̽� ��� ��T �C                �   �   ��  ��  ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                   �   �                      �������  ���    �                    ��� ���� �� �   ��  ��  ��  �  �   ��  ��                    �   ���                            �   �                                                                                                       �� ̽ ̽ ۽�}ک z�� ���
���
��̙�������̽��̘�̙��
� �	�"� �"  .  �
 �  �               �    ���                                    �   ̰  ��  ݚ� ��� ̽� �ͻ ��� �˘ ̸��ˉUP��UZ�UUJETDUDDUU33ET335[3�� ؚ  ��  +   "  �  ��   � �        �   �   @   �   �   �   �   �   �"  ""  !� �� ��  �               �   ������  ��           �   �    �   �       �   �   �                .                       �        �"�!/"�  �                                                                                                                                                                                  �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                    �   �   �   "   "   "  !�    ��                ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                       �   ���                            �   �                                                                                                                 � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �       ���                                                                                                                                                                                                        �  ��� ��� ��� �ݪ�                       �   �    �z� 
�� ������������ ˍ� ��� ���������ˉ����� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��                    ˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                                         �  ��  �� ��  ��                    �   �   ��  ��  ��  ɀ  �   ��  ��  ���   �   �   �                                                                                                                                                                                                                         �� ̚�
���	��������� �ܷ �� +� "� "+  ��UH"+��""��"+���   ��  ̸� ��� �͌��ݩ�g���gz��w���ت��ݚ���ɜЉ��К˽ ȭ� ��9 �UB �UB �T@ ED/ ��� ��� ������   ""  ""� �  �� ��   ��                                         � ��                +��"�"/� ""� "" �   �             ��  ���  �                      � ����  �                                 �              ����������                                ��  ��  ���                        "  "  "                                                                                                                                                                 �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��               � �                 �   �   �    ���                             "��"  �"  "   "                    �  ��  �                   �   �   �   �   P   P   P   P   U   E   ��  �ɠ ��� ���  �"  " ��"�""��"! � �  �   �   �   �                                                                                                           �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���          �     �  ��  ��   �                        �  ��            �   �    �                                ���� ��� ����                      �  �� ��  �    � ���                                                        ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                      	��ˋ����۪��ۚ{Ƚ�g˽˖�-��"�� .� 
�8 
�� 
D> DC �D0 �D 
�C U@ �� 	�� ��" , " "/ "/� �� �   �                    �   ��  ��  w�  k�� g�� w�� ��� �۹ ��� ��� 3̰ �  >�" 2� 2"�DC �3  ��  ��  +   "   "   "/� ��     �                               �  �� �  �  �   �                             �� ̽        �   ��  ��  ��  �   �                 �                        ���� ��� ����               �  �  �  �                            �  �˰ ��� �wp ���                                                                                                                                                                 ̰ ˻����wݩk}�gz� w�� �  �  � ^� UNMTNL�DB,��2"ʪ����� � �" ""/ ���    �    �   ��  ��  ��� ��� ��� ��� ���0۹�0؊�3���3˻�3���C��X��U��T�����  ��  �   �  "��" �"                  �"  ��  ��  �                                         �   �   ��  ��  ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                      �  �� ��  �    � ���                                                �   ���                            �   �                                                                                                                           �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��   �  �   
�  �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                             "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""����������D��M��M""""����������""""�����ADMA����""""����DD�M�""""��������AD�DM�""""�����������A�A�""""������AD�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��M��M�������D����3333DDDD�DD�M�D�������3333DDDDD�������M�DM�D����3333DDDD��A�M�M���M�����3333DDDDMM������D��D����3333DDDDA�A�A�D��M�D�����3333DDDD�������������D������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
� E �D � �B� � �K � �K � � K � �K � � 	K" � �
C. � �C1 � � C4 � �C5 � �C7 � Jk~ _ k� �"� � � "� � �"� � �*� � � "K � � "I �7 "& �? ", |": �/ "P �? !� �? !� �/  "G �/ "K �?  "B �?  "B �W  " |{"
� � #"E � �$* | �%!� |&"8 �/ '"E �/  "G �? !� �? !� � � +"& | �,"* | �-"2 | ."@ |/": �/ 0"P �? !� �/ 2"E �/  "G �
  *A� 5*Gx  *Ax  7*Ov  *Kv  *J�.  *E|K ;*Jw[ )�g=**} >*<e( *2u3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������ �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������.�O�T�U��-�O�I�I�G�X�K�R�R�O� � � � � �.�/�=�����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3�������������������������������������������-�N�X�O�Y�Z�G�T��;�[�[�Z�Z�[� � � � � �-�2�3�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������.�/�=� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�2�3� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�A�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                