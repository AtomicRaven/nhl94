GST@�                                                            \     �                                                ��         f  ��@         � 2�������ʲ���������    ����        ��      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"   "D�j��
� " ��
  B                                                                               ����������������������������������       ��    =b= 0Q0 44 111  4            	 
                    ��� �� � � ��                 nE 
)         8�����������������������������������������������������������������������������������������������������������������������������o  b  o   1  +    '           �                  	  7  V  	                  h  "          := �����������������������������������������������������������������������������                                D   L           @  &   �   �                                                                                 '    
)nE  "h    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E t �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    �l;AS��k��IY|, _�=����d��P $g#��T0 k� �G��K�eA"1�8	e1�D#�  ��?    � ���l;AS��k��IY|, _�-����d��Q g#��T0 k� �G��K�eA"1�8	e1�D#�  ��?    � ���l;AS��k��IY|, _�-����d��Q g#��T0 k� �K��O�eA"1�8	e1�D#�  ��?   � ���l;AS��o��IY|, _�-����d��Q gã�T0 k� �O��S�eA"1�8	e1�D#�  ��?    � ���l;AS��o��IY|, _�-����d�xQ gã�T0 k� �O��S�eA"1�8	e1�D#�  ��?    � ���l;AS��o��IY|, _�-����d�pQ  gã�T0 k� �S��W�eA"1�8	e1�D#�  ��?    � ���l;AS��o��IY|, _������d	�hQ�gã�T0 k� �S��W�eA"1�8	e1�D#�  ��?    � ���l;AS��o��IY|, _������d	�dQ�gã�T0 k� �W��[�eA"1�8	e1�D#�  ��?    � ���l;AS��o��IY|, _������d	�\Q�gã�T0 k� �[��_�eA"1�8	e1�D#�  ��?    � ���l;AS��o��IY|, _������d	�TQ�gã�T0 k� �[��_�eA"1�8	e1�D#�  ��?    � ���l;AS��o��IY|, _������d	�PQ�gã�T0 k� �_��c�eA"1�8	e1�D#�  ��?    � ���l;AS��o��IY|, _������d	�HQ�gã�T0 k� �c��g�eA"1�8	e1�D#�  ��?    � ���l;AS��o��IY|, _�����d	�DQ�gã�T0 k� �c��g�eA"1�8	e1�D#�  ��?    � ���l;AS��o��IY|, _�����d	�<Q�gã�T0 k� �g��k�eA"1�8	e1�D#�  ��?    � ���l;AR���o��IY|, _�����d	�8Q�g#��T0 k� �k��o�eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�� ��d	�4Q�g#��T0 k� �k��o�eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _����d	�,Q�g#��T0 k� �o��s�eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�^�d	�(Q�g#��T0 k� �o��s�eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�^�d	�$Q	��g#��T0 k� �s��w�eA"1�8	e1�D#�  ��?   � ���l;AR���o��JY|, _�^�d	� Q	��g#��T0 k� �w��{�eA"1�8	e1�D#�  ��?   � ���l;AR���o��JY|, _�^�d	�Q	��g#��T0 k� �w��{�eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�^�d�	�Q	��g#��T0 k� �{���eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�	^�d�	�Q	�|g#��T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�^�d�	�Q	�xg#��T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�^�d�	�Q	�pg#��T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _� ^�d�	�Q	�hgç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�$^�d�	�Q	�dgç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�(^�d�	�Q	�`gç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�(^�d�	�Q	�Xgç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�,^�d�	� Q	�Tgç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�0^�d�	� Q	�Pgç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�4n�d	��Q	�Hgç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�8n�d	��Q	�Dgç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�<n�d	��Q	�<gç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��JY|, _�@n�d	��Q�8gç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��KY|, _�Dn�d	��Q�0gç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��KY|, _�Hn�d	��Q�0gç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��KY|, _�P n�d�Q�,gç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��KY|, _�T"n�d�Q�,gç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��KY|, _�.X#n�d�Q(gç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��KY|, _�.\%n�d��Q$gç�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AR���o��KY|, _�.`'n�d��Q$gç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, _�.d(n�d��Q$gç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^��.l*n�d��Q gç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^��.p,n�c��Q hç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^��.t.n�c��Qhç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^��.x/n�c��Qhç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����1n�c��Qhç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����3n�c��Qhç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����4n�c.�Qhç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����6n�c.�Q/hç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����8n�c.�Q/hç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����9n�c.�Q/hç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����;n�b.�Q/hç�T0 k� ������eA"1�8	e1�D#�  ��U   � ���l;AR���o��KY|, ^����<n�b.�Q/hç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����>n�b.�Q/hç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����?n�b.�Q/iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����An�b.�Q/ iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����Bn�b.�Q/ iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����Dn�b.�Q.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^����Dn�b.�Q.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��KY|, ^��θEn�b.�R.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��LY|, ^��θEn�b.�S.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��LY|, ^��θFn�a.�S.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^��μFn�a�.�T.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^��μGn�a�.�T.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^��μHn�a�.�U.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^����Hn�a�.�V.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^����In�a�.�V.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^����In�a�.�W.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^����Jn�a�.�W.�iç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^����Jn�a�.�X.�jç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^����K^�a�.�X.�jç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^����K^�a�.�Y.�jç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��La�, ^����L^�a.�Y.�jç�T0 k� ������eA"1�8	e1�D#�  ��U    � ���l;AR���o��LY|, ^����L^�a.�Z.�jç�T0 k� ������eA"1�8	e1�D#�  ��U    � �����HcO��0��Y|, �7��o��8^�+�s��T3��T0 k� �0�4eA"1�8	e1�D#�  ��    �   �� �HcS��8�'�Y|, �?�w��@^�7�s�X3��T0 k� �8�<eA"1�8	e1�D#�  ��    �   ��R�W��@�/�a�, �K���H^�?�s�X"s��T0 k� �<�@eA"1�8	e1�D#�  ��    �   ��R�_��H�7�a�, �S����P^�G�s'�\"s��T0 k� �D�HeA"1�8	e1�D#�  ��    �   ��R�c��P�;�a�, �_����X^�O�s/�`"s��T0 k� �H	�L	eA"1�8	e1�D#�  ��    �   �(~R�k��d�K�a�, �o����h^�_�;�d"s�T0 k� �T�XeA"1�8	e1�D#�  ��    �   �0~R�o��l�S�a�, �{����p^�g�C��h"s�T0 k� �\�`eA"1�8	e1�D#�  ��    �   �8~R�s��t�[�a�, ������x^�o�G��h"s�T0 k� �`�deA"1�8	e1�D#�  ��    �   �@~R�{��|�c�a�, �������^�{�O��l"s�T0 k� �h�leA"1�8	e1�D#�  ��    �   H}R��͈�k�a�, �������^���S��p"s�T0 k� �l�peA"1�8	e1�D#�  ��    �   P}R���͐�s�a�, �������]���s[��p"s�T0 k� �t�xeA"1�8	e1�D#�  ��    �   �X}R���͘�{�a�, ��������]���s_�t"s�T0 k� �x�|eA"1�8	e1�D#�  ��    �   �h|R���ݨ͋�Y|, ��������]���sk�x3�T0 k� ���eA"1�8	e1�D#�  ��    �   �p|R���ݰ͓�Y|, �ǚ�����]���ss�|3�	T0 k� ���eA"1�8	e1�D#�  ��    �   �x|R���ݼ͗�Y|, �Ӛ�����\����w�|3�
T0 k� ���eA"1�8	e1�D#�  ��    �   ��{R�����͟�Y|, �ۚ�����\������|3�T0 k� ���eA"1�8	e1�D#�  ��    �   ��{R�����ͧ�Y|, ������\���Ӄ���3�T0 k� ���eA"1�8	e1�D#�  ��    �   ��zR�����ͷ�Y|, �����q�[���ӏ�����T0 k� ���eA"1�8	e1�D#�  $�    �   ��zR�����Ϳ�Y|, ����q�[���㓿����T0 k� ���eA"1�8	e1�D#�  ��    �   ��yR��������Y|, ���#�q�Z���㛾����T0 k� ���eA"1�8	e1�D#�  ��    �   ��xR���� ���Y|, 	��3�q�Y���㣼����T0 k� ���eA"1�8	e1�D#�  ��    �   ��xR�������Y|, 	'��?�rX���㧻s���T0 k� ���eA"1�8	e1�D#�  ��    �   r�wR�������Y|, 	/��G�rX��㯺s���T0 k� ���eA"1�8	e1�D#�  ��    �   r�wR�������Y|, 	7�rO��W��ӳ�s���T0 k� ���eA"1�8	e1�D#�  ��    �   r�uR����,���Y|, 	G�r_�� U��ӻ�s�s�T0 k� ���eA"1�8	e1�D#�  ��    �   r�uR����4��Y|, 	#O�rg��(T�'��÷�� s�T0 k� ���eA"1�8	e1�D#�  ��    �   r�tR����<��Y|, 	#W�ro��0S�/��Ƕ�� s�T0 k� ���eA"1�8	e1�D#�  ��    �   s rR����L��Y|, 	#g�r��<Q�?�sϴ���s�T0 k� ���eA"1�8	e1�D#�  ��    �   sqR����X�#�Y|, 	#k�r���DP�G�sӳ���C�T0 k� ���eA"1�8	e1�D#�  ��    �   �spR����`�+�Y|, 	s�r��rLO�O�s۲���C�T0 k� ���eA"1�8	e1�D#�  ��    �   �snR����p�;�Y|, 	�r��rXM�_�s����C�T0 k� ���eA"1�8	e1�D#�  ��    �   �s$mR����x�C�Y|, 	��r��r`L�g�s����C�T0 k� ���eA"1�8	e1�D#�  ��    �   �s,lR������K�Y|, 	��r��rdK�o�s����C�T0 k� ���eA"1�8	e1�D#�  ��    �   �c8iR������[�Y|, 	#��b��rpI��s����C�T0 k� ���eA"1�8	e1�D#�  ��    �   �c@hR������c�Y|, 	#��b��rxG���s�����S�T0 k� ���eA"1�8	e1�D#�  ��    �   �cDgR������k�Y|, 	#��b��r|F���s�����S�T0 k� � �� eA"1�8	e1�D#�  ��    �   �cPdR�����{�Y|, 	#��b��r�C���t����S�T0 k� �#��#eA"1�8	e1�D#�  ��    �   �cTcR�������Y|, 	��2��r�B���d����S�T0 k� �|%��%eA"1�8	e1�D#�  ��    �   �cXaR�������Y|, 	��2��r�@���d�s����T0 k� �t �x eA"1�8	e1�D#�  ��    �   �c\`R�������Y|, 	��2��b�?���d�s���� T0 k� �l�peA"1�8	e1�D#�  ��    �   �ch]R�������Y|, 	Ú2��b�<���d�s����"T0 k� �d�heA"1�8	e1�D#�  ��    �   �cl[R�������Y|, 	#Úb��b�:���$�s����"T0 k� �\�`eA"1�8	e1�D#�  ��    �   �cpZR�������Y|, 	#Úb��b�9���$�s��3�#T0 k� �`�deA"1�8	e1�D#�  ��    �   �3pXR�������Y|, 	#ǚb��b�7���$�s��3�$T0 k� �` �d eA"1�8	e1�D#�  ��    �   �3xUR������Y|, 	#Ǚb��b�4���$�s��3�%T0 k� �`"�d"eA"1�8	e1�D#�  ��    �   �3|SR������Y|, 	Ǚc�b�2���d�s��3�&T0 k� �`$�d$eA"1�8	e1�D#�  ��    �   �3|RR�#�� ���Y|, 	˙c�b�1���d�c��3�&T0 k� �\%�`%eA"1�8	e1�D#�  ��    �   �c�PR�'��(���Y|, 	˙c�b�/���d�c��3|'T0 k� �X%�\%eA"1�8	e1�D#�  ��    �   �c�NR�'��0���Y|, 	˙c�b�.��c��c��3|(T0 k� �X&�\&eA"1�8	e1�D#�  ��    �   �c�KR�+��@���Y|, 	˙c�R�*�c��c��3t)T0 k� �P'�T'eA"1�8	e1�D#�  ��    �  �c�HR�/��H���Y|, 	#˙c�R�)�c��c��3t*T0 k� �P(�T(eA"1�8	e1�D#�  ��    �  �#�ER�/��T��Y|, 	#ǙS�R�'�c��c��3p*T0 k� �L(�P(eA"1�8	e1�D#�  ��    �  �#�BR�3��\��Y|, 	#ǙS�R�%�c��c��3l+T0 k� �H)�L)eA"1�8	e1�D#�  ��    �  �#|@R�3��d��Y|, 	#ǚS�R�$�
c��c��sl+T0 k� �D*�H*eA"1�8	e1�D#�  ��    �  �#x=R�7��l��Y|, 	#ǚS���"�c��c��sh,T0 k� �@+�D+eA"1�8	e1�D#�  ��    �  �#x=R�7��t�#�Y|, �ǚS���!�c��c��sd,T0 k� �<,�@,eA"1�8	e1�D#�  �    �  �Sx=R�;����3�Y|, �ǛS���� c��c��s\-T0 k� �4,�8,eA"1�8	e1�D#�  ��    �  �Sx=R�?����;�Y|, �ǜS����$c��S���X-T0 k� �0*�4*eA"1�8	e1�D#�  ��    �  �St=R�?����C�Y|, �ǜS����$c��S���T-T0 k� �,)�0)eA"1�8	e1�D#�  ��    �  �St=R�C����K�Y|, �ǝ�����(c��S���P-T0 k� �('�,'eA"1�8	e1�D#�  ��    �  �St=R�G����[�Y|, �Ǟ�����(c��S���H-T0 k� � &�$&eA"1�8	e1�D#�  ��    �  �St=R�G����c�Y|, �ǟ�����(c��S��sD-T0 k� �(� (eA"1�8	e1�D#�  ��    �  �St=R�K����k�Y|, �Ǡ�����,c�S��s@-T0 k� �)�)eA"1�8	e1�D#�  ��    �  �ct=R�K����s�Y|, �ǡ�����,c�S��s<-T0 k� �*�*eA"1�8	e1�D#�  ��    �  �ct=R�K����{�Y|, �Ǣ�����,��S��s8.T0 k� �+�+eA"1�8	e1�D#�  ��    �  �ct=R�O���ߋ�Y|, �ä�����,!��S���,.T0 k� � +�+eA"1�8	e1�D#�  ��    �  �ct=R�S��� ߓ�Y|, �å��2��,"��S���(.T0 k� ��+� +eA"1�8	e1�D#�  ��    �  �ct=R�S���!���Y|, �æ��2�
�(#��S���$.T0 k� ��,��,eA"1�8	e1�D#�  ��    �  �ct=R�W���!���Y|, ÿ���2��($S�C��� .T0 k� ��,��,eA"1�8	e1�D#�  ��    �  �st=R�W��"���Y|, ÿ���2�2(&S�C��3.T0 k� ��,��,eA"1�8	e1�D#�  ��    �  �st=R�[��#���Y|, ӻ���R�2$'S�C��3.T0 k� ��,��,eA"1�8	e1�D#�  ��    �  �st=R�[��$	��Y|, ӻ����R�2$(S�C��3.T0 k� ��,��,eA"1�8	e1�D#�  ��    �  �st<R�_��,&	��Y|, ӷ����R��2 *SߓC��3 .T0 k� ��,��,eA"1�8	e1�D#�  ��    �  �st<R�_��4'	��Y|, ӳ����R��R *SߓC��2�.T0 k� ��,��,eA"1�8	e1�D#�  ��    �  �st<R�c��<(	��Y|, ӯ����R��R+C۔C��2�/T0 k� ��-��-eA"1�8	e1�D#�  ��    �  �sp<R�c��D)	/��Y|, ӯ����R��R,CהC��2�/T0 k� ��-��-eA"1�8	e1�D#�  ��    �  �sp<R�c��H*	/��Y|, ӫ����R��R-CӔ3��2�/T0 k� ��-��-eA"1�8	e1�D#�  ��    �  �sp<R�g��X,	/��Y|, 㣬���R��R.Cϔ3��2�/T0 k� ��.��.eA"1�8	e1�D#�  ��    �  �sp<R�g��\-	/��Y|, 㟬��R��R/C˕3��2�/T0 k� ��.��.eA"1�8	e1�D#�  ��    �  �sp<R�k��d.	��Y|, 㛬��B��R0CǕ3��2�/T0 k� �.��.eA"1�8	e1�D#�  ��    �  �sp<R�k��h0	��Y|, 㗬��B��R1CÕC��r�/T0 k� �.��.eA"1�8	e1�D#�  ��    �  sp<R�o��t2	�Y|, S��ÿB����2C��C�r�/T0 k� �.��.eA"1�8	e1�D#�  ��+    �  }sp<R�o��x3	�Y|, S����B����3C��C{�r�/T0 k� �.��.eA"1�8	e1�D#�  ��+    �  {sp<R�o��|5	 �Y|, S����B����4C��Cw�r�/T0 k� �/��/eA"1�8	e1�D#�  �+    �  tsp<R�s���6	 �Y|, S���������4C��Cs�r�/T0 k� �0��0eA"1�8	e1�D#�  ��/    �  nsp<R�s���9	 �Y|, Sw������a�5C��Ck�r�0T0 k� �l1�p1eA"1�8	e1�D#�  ��/    � 	 hsp<R�w�Ќ:	 �Y|, �o�����a�6C��Cg�r�0T0 k� �`2�d2eA"1�8	e1�D#�  ��/    � 
 bsp<R�w�А<	�Y|, �k����{�a�63��Cc�r�0T0 k� �T3�X3eA"1�8	e1�D#� ��/    �  \sp<R�w�Д=	�Y|, �c���Bw�a�73��C_�r�0T0 k� �H4�L4eA"1�8	e1�D#� ��/    �  Vsp<R�{�И>	�Y|, �_���Bo�a�73��S[�r�0T0 k� �84�<4eA"1�8	e1�D#� ��/    �  Psp<R�{�МA	#�Y|, �S�{�Bc�Q�93��SW���0T0 k� � 6�$6eA"1�8	e1�D#� ��/    �  Jsp<R�{�МB	 '�Y|, �K�s�B_�Q�9C��SS���0T0 k� �7�7eA"1�8	e1�D#� ��/    �  Dsp<R��РC	 '�Y|, �C�o�BW�Q�:C��SO���0T0 k� �8�8eA"1�8	e1�D#� ��/    �  ?sp<R��РD	 +�Y|, �;�g�BS�Q�:C��SK���0T0 k� ��8��8eA"1�8	e1�D#�  ��/    �  :sp<R��РF	 +�Y|, �7�_�BO�Q�:C�SG���0T0 k� ��9��9eA"1�8	e1�D#�  ��/    �  5sp<Ră�ФG	 /�Y|, �/�W��G��;C{�SG���0T0 k� ��:��:eA"1�8	e1�D#�  ��/    �  0sp<Ră��H	/�Y|, �'�O��C��;Cw�SC���0T0 k� ��;��;eA"1�8	e1�D#�  ��/    �  +sp<Ră��I	/�Y|, ���G��;��<Cw�S?���0T0 k� ��<��<eA"1�8	e1�D#�  ��/    �  &sp<Ră��J	3�Y|, ���?��3��<Cs�S;�r�0T0 k� �<��<eA"1�8	e1�D#�  ��/    �  !sp<Rć��K	3�Y|, ���7��/��=Co�c;�r�0T0 k� �=��=eA"1�8	e1�D#�  ��/    �  sp<Rć��L	3�Y|, ���/��'��x=Ck�c7�r|0T0 k� �>��>eA"1�8	e1�D#�  ��/    �  sl<Rć��L	 3�Y|, ����#��#��p>Cg�c3�rx1T0 k� �?��?eA"1�8	e1�D#�  ��/    �  sl<Rć��M	 3�Y|, ��������h>Cc�c/�rt1T0 k� �@��@eA"1�8	e1�D#�  ��/    �  sl<Rċ��N	 3�Y|, �������`?S_�c/�rt1T0 k� �t@�x@eA"1�8	e1�D#�  ��/    �  sl<Ut���O	 3�Y|, �������X?S_�c+�rp1T0 k� �hA�lAeA"1�8	e1�D#�  ��/    �  sl<Ut���O	 3�Y|, �ۭ�����P?S[�c'�rl1T0 k� �\B�`BeA"1�8	e1�D#�  ��/    �  sl<Ut���P `3�Y|, �ӭ�����QD@SW�c'�rh1T0 k� �LC�PCeA"1�8	e1�D#�  ��/    �  sl<Ut���P `3�Y|, �˭�����Q<@SS�c#�rd1T0 k� �8E�<EeA"1�8	e1�D#�  ��(    �   sl<Ut���P `3�Y|, �������Q4ASO�c�rd1T0 k� �(F�,FeA"1�8	e1�D#�  ��(    � ��sl<Ut�� �Q `3�Y|, �������Q,ASO�c�r`1T0 k� �G� GeA"1�8	e1�D#�  ��(    � ��sl<Ut�� �Q `3�Y|, ���۬���Q$ASK�s�r\1T0 k� �H�HeA"1�8	e1�D#�  ��(    � ��sl<Ut�� �Q �3�Y|, ���Ӭ���QBSG�s�rX1T0 k� �H�HeA"1�8	e1�D#�  ��(    � ��sl<Ut�� �Q �3�Y|, ���˫���QBSG�s�rX1T0 k� ��I� IeA"1�8	e1�D#�  ��(    � ��sl;A��� �R �3�Y|, ������QBSC�s�rT1T0 k� ��I��IeA"1�8	e1�D#�  ��(    � ��sl;A���РR �3�Y|, ������QCc?�s�rP1T0 k� ��I��IeA"1�8	e1�D#�  ��(    � ��sl;A���РR �3�Y|, �����P�Cc;�s��L1T0 k� ��J��JeA"1�8	e1�D#�  ��(    � ��sl;A���ФR 3�Y|, s�����`�Cc;�s��L1T0 k� ��H��HeA"1�8	e1�D#�  ��(    � ��sl;A���ФR 3�Y|, k�����`�Dc7�s��H1T0 k� �G��GeA"1�8	e1�D#�  ��(    � ��sl;A���ФR 3�Y|, _�����`�Dc7�s��D1T0 k� �G��GeA"1�8	e1�D#�  ��(    � ��sl;A���p�Q 3�Y|, W�����`�Dc3�s��D1T0 k� �F��FeA"1�8	e1�D#�  ��(    � ��sl;A���p�Q 3�Y|, K������`�Dc/�s�rD0T0 k� ��E��EeA"1�8	e1�D#�  �(    � ��sl;A���p�R�3�Y|, C�������Cc/�C�r@0T0 k� �D��DeA"1�8	e1�D#�  ��(    � ��sl;A���p�R�/�Y|, ;�s������Cc+�B��r@0T0 k� �B��BeA"1�8	e1�D#�  ��(    � ��sl;ET��p�R�/�Y|, /�k������Bc'�B��r@0T0 k� �A��AeA"1�8	e1�D#�  ��(    � ��sl;ET�� �S�/�Y|, '�c�����Bc'�B��r@0T0 k� �@��@eA"1�8	e1�D#�  ��(    � ��sl;ET�� �S�+�Y|, �[��{�иBs#�B�r@0T0 k� �?��?eA"1�8	e1�D#�  ��(    � ��sl;ET�� �R�+�Y|, �S��s��As#�2�r@0T0 k� ��:��:eA"1�8	e1�D#�  ��(    � ��sl;ET�� �Q�+�Y|, �K��k��@s�2��@/T0 k� ��5��5eA"1�8	e1�D#�  ��(    � ��sl;ET�� �Q�'�Y|, ��C��c��@s�2��D/T0 k� ��1��1eA"1�8	e1�D#�  ��(    � ��sl;ET����P�'�Y|, ��;��[��?s�2�
�D/T0 k� �|/��/eA"1�8	e1�D#�  ��(    � ��sl;ET����P�#�Y|, ��3��S���>s�2��D/T0 k� �x,�|,eA"1�8	e1�D#�  ��(    � ��sl;ET����O��Y|, ��'��K���=s�2��H/T0 k� �l,�p,eA"1�8	e1�D#�  ��(    � ��sl;C����N��Y|, �׮��C���<s�"��L/T0 k� �`,�d,eA"1�8	e1�D#�  ��(    � ��sl;C����M��Y|, �Ϯ��;���<s�"��L/T0 k� �X,�\,eA"1�8	e1�D#�  ��(    � ��sl;C����M��Y|, �Ǯ��3���;s�"��P/T0 k� �P+�T+eA"1�8	e1�D#�  ��(    � ��sl;C����L��Y|, Ữ��/��x:	S�"��T/T0 k� �H*�L*eA"1�8	e1�D#�  ��(    � ��sl;C�{���K��Y|, ᳮ���'��p9	S�"��X.T0 k� �@)�D)eA"1�8	e1�D#�  ��(    � ��sl;C�w���K��Y|, ᧮�����h8	S�"��\.T0 k� �8(�<(eA"1�8	e1�D#�  ��(    � ��sl;C�s���J��Y|, ៮����`7	S�"��`.T0 k� �4'�8'eA"1�8	e1�D#�  ��(    � ��sl;C�o���J��Y|, ᓮ����\5	S�"��d.T0 k� �,&�0&eA"1�8	e1�D#�  ��(    � ��sl;C�k���I��Y|, ዮۡ���T4	S�"�!�h.T0 k� �$%�(%eA"1�8	e1�D#�  ��(    � ��sl;C�c���H��Y|, �w�ˠ����D2	c�"�%�p-T0 k� �#�#eA"1�8	e1�D#�  ��(    � ��sl;C�[���G��Y|, �o��à����<1	c�"�' Rt-T0 k� �!�!eA"1�8	e1�D#�  ��(    � ��sl;C�W���F��Y|, �c�໠����40	c�"�) R|,T0 k� � � eA"1�8	e1�D#�  ��(    � ��sl;C�S���F��Y|, �[�೟����0/	c�"�+ R�,T0 k� � �eA"1�8	e1�D#�  ��(    � ��sl;C�K���E��Y|, �S�૟���P(.	c�"�- R�+T0 k� ��$� $eA"1�8	e1�D#�  �(    � ��sl;C�G���E_��Y|, �G�������P -����/ R�+T0 k� ��'��'eA"1�8	e1�D#�  �(    � ��sl;C�C���D_��Y|, Q?�P�����P+����1 R�*T0 k� ��)��)eA"1�8	e1�D#�  ��(    � ��sl;AT;���D_��Y|, Q7�P�����P*����3 b�)T0 k� ��*��*eA"1�8	e1�D#�  ��(    � ��sl;AT7���C_��Y|, Q+�P���� P)����5 b�)T0 k� ��+��+eA"1�8	e1�D#�  ��(    � ��sl;AT3���C_��Y|, Q#�P���P(����7 b�(T0 k� ��+��+eA"1�8	e1�D#�  ��(    � ��sl;AT/���B_��Y|, Q�Pw���_�'�����9 b�'T0 k� ��*��*eA"1�8	e1�D#�  ��(    � ��sl;AT'���B_��Y|, Q�Po���_�&�����; b�&T0 k� ��*��*eA"1�8	e1�D#�  ��(    � ��sl;AT#���A_��Y|, Q�Pg���_�%�����= b�%T0 k� ��*��*eA"1�8	e1�D#�  ��(    � ��sl;AT�p�@_��Y|, P��P[���_�$�����? b�$T0 k� ��*��*eA"1�8	e1�D#�  ��(    � ��sl;AT�p�@_��Y|, P��PS���_�#�����B b�#T0 k� ��)��)eA"1�8	e1�D#�  ��(    � ��sl;AT�p�?_��Y|, P�@K���_�"�����D b�"T0 k� ��)��)eA"1�8	e1�D#�  ��(    � ��sl;AT�q >_��Y|, P�@C���_�!�����F b�!T0 k� ��(��(eA"1�8	e1�D#�  ��(    � ��sl;AT�q>_��Y|, P߯@;��|
_� �����H b� T0 k� ��'��'eA"1�8	e1�D#�  ��(    � ��sl;AT�q=_��Y|, Pۯ@3��tO� �����J b�T0 k� ��)��)eA"1�8	e1�D#�  ��(    � ��sl;AT�q<_��Y|, Pӯ@+��lO������L b�T0 k� ��*��*eA"1�8	e1�D#�  ��(    � ��sl;AS��a;_��Y|, P˯@��dO�����N b�T0 k� ��*��*eA"1�8	e1�D#�  ��(    � ��sl;AS��a:_��Y|, Pï@��`O����P b�T0 k� ��+��+eA"1�8	e1�D#�  ��(    � ���l;AS��a9_��Y|, P��@��XO����R b�T0 k� �|+��+eA"1�8	e1�D#�  ��(    � ���l;AS��a8_��Y|, P�����Po����T 3 T0 k� �t*�x*eA"1�8	e1�D#�  ��8    � ���l;AS��a7��Y|, P������Ho����V 3T0 k� �l*�p*eA"1�8	e1�D#�  ��8    � ���l;AS��a6��Y|, P������Do����Y 3T0 k� �d)�h)eA"1�8	e1�D#�  ��8    � ���l;AS��a5��Y|, P�����<o����[ 3T0 k� �\(�`(eA"1�8	e1�D#�  ��8    � ���l;AS��a5��Y|, P�����4ox�	��] 3T0 k� �T(�X(eA"1�8	e1�D#�  ��8    � ���l;AS��a4��Y|, P���ߝ�,op�
��_ 3$T0 k� �L'�P'eA"1�8	e1�D#�  ��8   � ���l;AS��a3O��Y|, P���ם�(_h���a 3(T0 k� �D'�H'eA"1�8	e1�D#�  ��8    � ���l;AS��a2O��Y|, P���ϝ� _`���c 30T0 k� �@&�D&eA"1�8	e1�D#�  ��8    � ��cl;AS��a1O��a�, P��ǝ�_\"���e 38T0 k� �8&�<&eA"1�8	e1�D#�  ��8    � ��cl;AS��a0O�a�, Pw�����_T"���g 3@T0 k� �0%�4%eA"1�8	e1�D#�  ��8    � ��cl;AS���/O{�a�, Ps�����_L"���i 3DT0 k� �(%�,%eA"1�8	e1�D#�  ��8    � ��cl;AS���/Ow�a�, Pk�����_D"���k 3DT0 k� �$$�($eA"1�8	e1�D#�  ��8    � ��cl;AS���.Os�a�, Pg������_@"���n CDT0 k� �$� $eA"1�8	e1�D#�  ��8    � ��cl;AS��� -Oo�a�, Pc������_8"���p CDT0 k� �#�#eA"1�8	e1�D#�  ��8    � ��cl;AS��� ,Ok�a�, P[����� _4"���r CDT0 k� �#�#eA"1�8	e1�D#�  ��8    � ��cl;AS��� +Oc�a�, PW�����"_,"���t CDT0 k� �"�"eA"1�8	e1�D#�  ��8    � ��cl;AS��� +O_�a�, PO�����#o("���v CDT0 k� �"�"eA"1�8	e1�D#�  ��8    � ���l;AS���$*?[�a�, PK�����$o "���x�DT0 k� ��!� !eA"1�8	e1�D#�  ��8    � ���l;AS���$)?W�a�, PG�����%o"��z�DT0 k� ��!��!eA"1�8	e1�D#�  ��8    � ���l;AS���$(?S�Y|, P?�{���&o"��|�DT0 k� �� �� eA"1�8	e1�D#�  ��8    � ���l;AS���((?O�Y|, P;�w���(o"��}�DT0 k� ����eA"1�8	e1�D#�  �8    � ���l;AS���('?K�Y|, P7�o���)"���DT0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS���(&OG�Y|, P/�k���*"��� 3HT0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS���(&OC�Y|, P+�c���+~�"��� 3HT0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS���,%O?�Y|, P'�_���-~�"��� 3HT0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS���,$O;�Y|, P#�W���.~�"��� 3HT0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS���,$O,Y|, P�S���/��"�� 3HT0 k� �l�peA"1�8	e1�D#� ��?    � ���l;AS���,#�$Y|, P�K���0��"�� 3LT0 k� �X�\eA"1�8	e1�D#� ��?    � ���l;AS���0"�Y|, P�G���2��"� "��LT0 k� �H�LeA"1�8	e1�D#� ��?    � ���l;AS���0"�Y|, P�C���3��"�!"�~�LT0 k� �4�8eA"1�8	e1�D#� �?    � ���l;AS���0!�a�, P�;���4��"�""�~�PT0 k� � �$eA"1�8	e1�D#� ��?    � ���l;AS���0!�a�, P�7��|5��"�""�}�PT0 k� ��eA"1�8	e1�D#� ��?    � ���l;AS���0 Oa�, P�3��x7��"�#"�}�PT0 k� ��� eA"1�8	e1�D#� ��?    � ���l;AS���4 Oa�, _��+��p8��"�$"�}�TT0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS���4O	a�, _��'��h9޸"�%"�|�TT0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS���4N�
a�, _��#��d:ް"�%"�|�TT0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS���4N�a�, _���\<ި"�&"�{�TT0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS���4N�a�, _���X=�"�'"�{�X
T0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS���8N�a�, _���P>�"�'"�{�X
T0 k� ����eA"1�8	e1�D#� ��?    � ���l;AS��8N�a�, _���H@�"�("�z�X
T0 k� �x
�|
eA"1�8	e1�D#� ��?   � ���l;AS{��8N�a�, _���DA�"�)"�z�\
T0 k� �d�heA"1�8	e1�D#� ��?    � ���l;AS{��8N�Y|, _߯��<B�"�)"�z�\	T0 k� �T�XeA"1�8	e1�D#� ��?    � ���l;ASw��8N�Y|, _ۯ�	4C�"�*"�y�\	T0 k� �@�DeA"1�8	e1�D#� ��?    � ���l;ASw��<N�Y|, _ׯ��	0E�|"�+"�y�\	T0 k� �,�0eA"1�8	e1�D#� ��?    � ���l;ASs��<N�Y|, _ӯ��	,F�x"�+"�y�`	T0 k� ��eA"1�8	e1�D#� ��?    � ���l;ASs��<N�Y|, _ϯ��	$G�p"�,"�x�`T0 k� ��eA"1�8	e1�D#� ��?    � ���l;ASo��<N�Y|, _ϯ�	 H�l"�,"�x�`T0 k� ����eA"1�8	e1�D#� ��?    � ���l;ASo��<N�Y|, _˯�	I�d"�-"�x�`T0 k� �� �� eA"1�8	e1�D#� ��?    � ���l;ASo��<N�Y|, _ǯ�	�J�`"�."�x�dT0 k� ������eA"1�8	e1�D#� ��?    � ���l;ASk��@N�Y|, _ï�	�K�\�."�w�dT0 k� ������eA"1�8	e1�D#� ��?   � ���l;ASk��@N�Y|, _���	�K�T�/"�w�dT0 k� ������eA"1�8	e1�D#� ��?    � ���l;ASg��@N�Y|, _��ߠ	�L�P�/"�w�dT0 k� ������eA"1�8	e1�D#� ��?    � ���l;ASg��@N�Y|, _��۠	�M�L�0"�v�hT0 k� ������eA"1�8	e1�D#� ��?    � ���l;ASc��@N�Y|, _��נ	 M�D�0"�v�hT0 k� �s��w�eA"1�8	e1�D#� ��?    � ���l;ASc��@N�Y|, _��Ӡ	~�N�@�1"�v�hT0 k� �_��c�eA"1�8	e1�D#� $�?    � ���l;AS_��DN�Y|, _���Ϡ	~�O�<�1"�v�hT0 k� �c��g�eA"1�8	e1�D#� ��?    � ���l;AS_��DΨY|, _���ˠ	~�P�4�2"�u�lT0 k� �g��k�eA"1�8	e1�D#� ��?    � ���l;AS_��DΤY|, _���Ǡ	~�Q�0�2"�u�lT0 k� �k��o�eA"1�8	e1�D#� ��?    � ���l;AS[��DΠY|, _���à>�Q�,�3"�u�lT0 k� �o��s�eA"1�8	e1�D#� ��?    � ���l;AS[��DΜY|, _���à>�R�(�3"�u�lT0 k� �o��s�eA"1�8	e1�D#� ��?    � ���l;ASW��DΘY|, _�����>�S�$�4"�t�lT0 k� �s��w�eA"1�8	e1�D#� ��?    � ���l;ASW��DΔY|, _��N��>�T��4"�t�pT0 k� �w��{�eA"1�8	e1�D#� ��?    � ���l;ASW��HΐY|, _��N��>�U��5"�t�pT0 k� �{���eA"1�8	e1�D#� ��?    � ���l;ASS��HΌY|, _��N��>�W��5"�t�pT0 k� �����eA"1�8	e1�D#� ��?    � ���l;ASS��HΈ Y|, _��N��.�X��6"�s�pT0 k� �����eA"1�8	e1�D#� ��?    � ���l;ASS��H΄!Y|, _��N��.�Y��6"�s�pT0 k� ������eA"1�8	e1�D#� ��?    � ���l;ASO��H�!Y|, _��>��.�Z��7"�s�tT0 k� ������eA"1�8	e1�D#� ��?    � ���l;ASO��H�"Y|, _��>��.�[��7"�s�tT0 k� ������eA"1�8	e1�D#� ��?    � ���l;ASO��H|#Y|, _��>��.�\� �7"�r�tT0 k� ������eA"1�8	e1�D#� ��?    � ���l;ASK��Lx#Y|, _��>��.�^���8�r�tT0 k� ������eA"1�8	e1�D#� ��?    � ���l;ASK��Lt$Y|, _��>��.�_���8�r�tT0 k� �����eA"1�8	e1�D#� ��?    � ���l;ASK��Lp%Y|, _��N��.�`���9�r�tT0 k� �����eA"1�8	e1�D#� ��?    � ���l;ASG��Ll%Y|, _��N��.�b���|9�r�xT0 k� �����eA"1�8	e1�D#� ��?    � ���l;ASG��Ll&Y|, _��N��.�c���x9�q�xT0 k� �����eA"1�8	e1�D#� ��?   � ���l;ASG��Lh&Y|, _�N��.�d���x:�q�xT0 k� �����eA"1�8	e1�D#� ��?    � ���l;ASC��Ld'Y|, _�N���e���p:��q�xT0 k� �����eA"1�8	e1�D#�  ��?    � ���l;ASC��L`'Y|, _{�ޏ��g���l;��q�xT0 k� �����eA"1�8	e1�D#�  ��?    � ���l;ASC��L`(Y|, _{�ދ��h���h;��q�xT0 k� �����eA"1�8	e1�D#�  -�?    � ���l;AS?��P\)Y|, _w�އ��i��d;��q�|T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AS?��PX)Y|, _w�އ��k��`<��p�|T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AS?��PX*Y|, _s�ރ���l��\<��p�|T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AS?��PT*Y|, _s�����m��X<��p�|T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AS;��PP+Y|, _o�����n��P=��p�|T0 k� �����eA"1�8	e1�D#� ��?    � ���l;AS;��PP+Y|, _o��{���o��L=��p�|T0 k� �����eA"1�8	e1�D#� ��?    � ���l;AS;��PL,Y|, _k��{���p��H=��o�|T0 k� ������eA"1�8	e1�D#� ��?    � ���l;AS7��PH,Y|, _k��w���r��D>��oÀT0 k� ������eA"1�8	e1�D#� ��?    � ���l;AS7��PH-Y|, _g��w���s��<>��oÀT0 k� ������eA"1�8	e1�D#� ��?    � ���l;AS7��TD-Y|, _g��s���t��8>��oÀT0 k� ������eA"1�8	e1�D#� ��?    � ���l;AS7��T@.Y|, _c��o���u��0?��oÀT0 k� ������eA"1�8	e1�D#� ��?    � ���l;AS3��T
@.Y|, _c��o���v��,?��oÀ T0 k� ������eA"1�8	e1�D#� ��?    � ���l;AS3��T
</Y|, _c��k���w��$?��oÀ T0 k� ������eA"1�8	e1�D#� ��?    � ���l;AS3��T
</Y|, __��k���x�� @��nÀ T0 k� ������eA"1�8	e1�D#� ��?    � ���l;AS3��T
80Y|, __��g���y��@��nÄ T0 k� ������eA"1�8	e1�D#� ��?    � ���l;AS3��T
40Y|, _[��g���z��@��nÄ T0 k� ������eA"1�8	e1�D#� ��?   � ���l;AS/��T	40Y|, _[��c���{��@�nÄ T0 k� ������eA"1�8	e1�D#� ��?    � ���l;AS/��T	01Y|, _[��c���|��A�nÄ T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS/��T	01Y|, _W��_���}�� A�nÄ T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS/��T	,2Y|, _W��_���~���A�nÇ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS+��T	,2Y|, _S��[������B�mÇ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS+��X(3Y|, _S��[�������B�mÇ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS+��X(3Y|, _S��W������B�mÇ�T0 k� �����eA"1�8	e1�D#�  /�?    � ���l;AS+��X$3Y|, _O��W������B�mË�T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AS+��X$4Y|, _O��S������C�mË�T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AS'��X 4Y|, _O��S������C�mË�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS'��X 4Y|, _K��S���~���C�mË�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS'��X5Y|, _K��O���~���C�mË�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS'��X5Y|, _K��O���~���D�lË�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS'��X6Y|, _G��K���~���D|lË�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS'��X6Y|, _G��K���~���DxlË�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS#��X6Y|, _G��K���}���DplË�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS#��X7Y|, _C��G���}���DllÏ�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS#��X7Y|, _C��G���}��!�EdlÏ�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS#��\7Y|, _C��C���}��!�E`lÏ�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS#��\8Y|, _?��C���|�|!�EXlÏ�T0 k� ���#�eA"1�8	e1�D#�  ��?    � ���l;AS#��\8Y|, _?��C���|�|!�EPlÏ�T0 k� ���#�eA"1�8	e1�D#�  ��?    � ���l;AS��\8Y|, _?��?���|�x!�FLkÏ�T0 k� �#��'�eA"1�8	e1�D#�  ��?    � ���l;AS��\9Y|, _?��?���|�x!�FDkÏ�T0 k� �'��+�eA"1�8	e1�D#�  ��?    � ���l;AS��\9Y|, _;��?���|�t!�F@kÏ�T0 k� �+��/�eA"1�8	e1�D#�  ��?    � ���l;AS��\9Y|, _;��;���{�t!�F8kÏ�T0 k� �+��/�eA"1�8	e1�D#�  ��?    � ���l;AS��\9Y|, _;��;���{�p!�F0kÏ�T0 k� �/��3�eA"1�8	e1�D#�  ��?    � ���l;AS��\:Y|, _;��;���{�p!�G�(kÏ�T0 k� �3��7�eA"1�8	e1�D#�  ��?    � ���l;AS��\:Y|, _7��7���{�l!|G� kÏ�T0 k� �7��;�eA"1�8	e1�D#�  ��?    � ���l;AS��\ :Y|, _7��7���{�l!xG�kÓ�T0 k� �7��;�eA"1�8	e1�D#�  ��?    � ���l;AS��\ ;Y|, _7��7���{�l!tG�kÓ�T0 k� �;��?�eA"1�8	e1�D#�  ��?    � ���l;AS��\ ;Y|, _7��3���z�h!pG�kÓ�T0 k� �?��C�eA"1�8	e1�D#�  ��?    � ���l;AS��\�;Y|, _3��3���z�h!lG�kÓ�T0 k� �C��G�eA"1�8	e1�D#�  ��?    � ���l;AS��\�;Y|, _3��3���z�d!hH��kÓ�T0 k� �C��G�eA"1�8	e1�D#�  ��?    � ���l;AS��\�<Y|, _3��/���z�d!dH��jÓ�T0 k� �G��K�eA"1�8	e1�D#�  ��?   � ���l;AS��\�<Y|, _3��/���z�d!`H��jÓ�T0 k� �K��O�eA"1�8	e1�D#�  ��?    � ���l;AS��`�<Y|, _/��/���z�`!\H��jÓ�T0 k� �O��S�eA"1�8	e1�D#�  ��?    � ���l;AS��`�<Y|, _/��/���y�`!XH�jÓ�T0 k� �O��S�eA"1�8	e1�D#�  ��?    � ���l;AS��`�=Y|, _/��+���y�\!TH�jÓ�T0 k� �S��W�eA"1�8	e1�D#�  ��?    � ���l;AS��`�=Y|, _/��+���y�\!PI�jÓ�T0 k� �W��[�eA"1�8	e1�D#�  ��?    � ���l;AS��`�=Y|, _+��+���y�\!LI�jÓ�T0 k� �[��_�eA"1�8	e1�D#�  ��?    � ���l;AS��`�=Y|, _+��+���y�X!HI�jÓ�T0 k� �[��_�eA"1�8	e1�D#�  ��?    � ���l;AS��`�>Y|, _+��'���y�X!DI�j×�T0 k� �_��c�eA"1�8	e1�D#�  ��?    � ���l;AS��`�>Y|, _+�N'���y�X!@I�j×�T0 k� �c��g�eA"1�8	e1�D#�  ��?    � ���l;AS��`�>Y|, _+�N'���x�T!<I�j×�T0 k� �g��k�eA"1�8	e1�D#�  ��?    � ���l;AS��`�>Y|, _'�N#� �x�T!<J�j×�T0 k� �g��k�eA"1�8	e1�D#�  ��?    � ���l;AS��`�?Y|, _'�N#� �x�T!8J�j×�T0 k� �k��o�eA"1�8	e1�D#�  ��?    � ���l;AS��`�?Y|, _'�N#� �x�P!4J�i×�T0 k� �o��s�eA"1�8	e1�D#�  ��?    � ���l;AS��`�?Y|, _'�N#� �x�P!0J�i×�T0 k� �s��w�eA"1�8	e1�D#�  ��?    � ���l;AS��`�?Y|, _'�N#� �x�P!,J�i×�T0 k� �s��w�eA"1�8	e1�D#�  ��?    � ���l;AS��`�?Y|, _'�N�޸w�L!,J�i×�T0 k� �w��{�eA"1�8	e1�D#�  ��?    � ���l;AS��`�@Y|, _#�N�޸w�L!(J!|i×�T0 k� �{���eA"1�8	e1�D#�  ��?    � ���l;AS��`�@Y|, _#�N�޸wL!$J!xi×�T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AS��`�@Y|, _#���޼wH! K!pi×�T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AS��`�@Y|, _#���޼vH! K!li×�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��`�@Y|, _#���޼vH!K!di×�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��`�AY|, _#�����uH!K!`i×�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�AY|, _�����uD!K!Xi×�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�AY|, _�����uD!K!TiÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�AY|, _�����tDK!PiÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�AY|, _�����sDK!HiÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�AY|, _�����sM@L!DiÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�BY|, _�����rM@L!@iÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�BY|, _�����rM@L!8iÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�BY|, _���~�qM@L!4iÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�BY|, _���~�pM<� L!0iÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�BY|, _���~�oM<� L!(hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�BY|, _���~�oM<��L!$hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�CY|, _���~�nM<��L! hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�CY|, _�����mM8��L!hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�CY|, _�����l8��M!hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d�CY|, _�����k8��M!hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �CY|, _�����j8��M!hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �CY|, _�����j4��M!hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �CY|, _�����i4��M!hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �DY|, _�����h4��M! hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �DY|, _�����h�4��M �hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �DY|, _�����g�4��M �hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �DY|, _�����g�0��M �hÛ�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �DY|, _�����f�0��M �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �DY|, _�����f�0��N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �DY|, _�����f�0��N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �EY|, _�����e�0��N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �EY|, _�����e�0�N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �EY|, _�����e�,�N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��d �EY|, _�����e�,�N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��h �EY|, _�����e,�N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��h �EY|, _�����d,�N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��h �EY|, _�����d, �N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��h �EY|, _�����d( �N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��k��FY|, _�����d( �N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��k��FY|, _�����d( �N �hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��k��FY|, _�����d( �N�hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��k��FY|, _�����d( �O�hß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��k��FY|, _�����d( |O�gß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��k��FY|, _�����d�( tO�gß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��k��FY|, _�����d�$ lO�gß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��k��FY|, _�����d�$ hO�gß�T0 k� ������eA"1�8	e1�D#�  ��?    � ���l;AS��k��FY|, _�����d�$ `O�gß�T0 k� �����eA"1�8	e1�D#�  ��?    � ���l;AS��k��FY|, _�����d�$XO�gß�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _�����d�$TO�gß�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _������d�$LO�gß�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _������d�$DO�gß�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _������d� <O��gß�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _������d 8O��gß�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _������d 0O��gß�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _������d (O��gß�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _������d  O��gã�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _������d P��gã�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _������d P��gã�T0 k� ����eA"1�8	e1�D#�  ��?    � ���l;AS��k��GY|, _������d �P�|gã�T0 k� ���#�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _������d� P�xgã�T0 k� �#��'�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _������d��P�tgã�T0 k� �#��'�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _������d��P�lgã�T0 k� �'��+�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _�M����d��P�hgã�T0 k� �+��/�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _�M����d��P�dgã�T0 k� �+��/�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _�M����d��P�\gã�T0 k� �/��3�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _�M����d��P�Xg#��T0 k� �/��3�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _�M����d��P�Pg#��T0 k� �3��7�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _�M����d��P�Lg#��T0 k� �7��;�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _�=����d�P�Dg#��T0 k� �7��;�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _�=����d�P @g#��T0 k� �;��?�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _�=����d��P 8g#��T0 k� �?��C�eA"1�8	e1�D#�  ��?    � ���l;AS��k��HY|, _�=����d��P 0g#��T0 k� �?��C�eA"1�8	e1�D#�  ��?    � ���l;AS��k��IY|, _�=����d��P ,g#��T0 k� �C��G�eA"1�8	e1�D#�  ��?    � ��                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��� ]�1-1- � �� ;��   '	 � �"�     ;�� �"�                 	 	            [P     ���   0

 	 	         ����  +     � �j,    ���� �j�      ��   
                        ���   (	          ����            [��    ���� [��    ��            	   ��          |      ���   (
	           Lp�          �l��     Li��l��     k��                �$          ��      ��� @ P
B 	           �� ��	      .�X�      ���X�                              �K                ���   8		 1 	            ���     	    B����    ������z      ��   
        m �         �     ���   8
�          L�;  � �
	   V���@     LM���z�    ��           = Z��         �@�    ��`   8
	
          a  � �	   j����     a ���Ma    ����          ] 	 Z��         � �    ��`  0           ��  � �
	   ~�B�|     ���B�2      ��           s  Z��          ���    ��h   		�           Z��  � �
	   ����     Y�N���o    �             0	 Z��         	 ��    ��`   @4          j>y  � �
	   ���o�     j/�����     ��           g Z��         
 ���    ��`@ H
		         ���! ��     � �    ���! �s                            �� ;             �  ��@    0 )                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         ���K  ��        ���]    ���K��      �� "                x                j  �       �                         ��    ��       ���      ��  ��           "                                                 �                          � � [�l��������B���� �������      
    	       
  2    s Oz�G       ۤ  o� �� p  � `p  �� p� �� q  � q  �D s� �d s� ̄ 0m� �� n@ � 0n` �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À���� ����� � 
�| V ���� � 
� V� 
�| W ���� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �������� �� B  ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"   "D�j�
�� " �
� �  �  
� ��    ��     ���      ��    ��     ���           ��     ��B          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �U���      �� �  ���        � �T ��        �        ��        �        ��        �    ��    ������B�        ��                         T�) ,  ����                                     �                ����            �������%��   ����               25/47 (53%) rchuk  k   4:19                                                                        6  6      �C
� �Mc~ �O c� �]c� �l c� �V c� �N c� �*C(B	C"8 �
cjAcnA �cp) �cs! � cw9 cx( � � � � � � �cV& � c^& � c_6 �c`6 � cb. � cc+ �c�E � c�U � c�= � c�@ � c�F � c�H �c�5 � c�E �  c�- � !c�0 � "c�6 � #c�8 �$CB � � %CJ � �&"� � � '"� � �(� � �)
� � �*"� � � +"� � �,"� � �-*� �w."� �w /"� �g0� �g 
� � �2"�  � 3"�2 �4� � 
�' �6� � 
�' �8� � 
�' �:"P � ;*O� �  *H� � =*O� �  *H�@ *<t                                                                                                                                                                                                                         �� P         �     @ 
        �     a P E a  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    ���� ��������������������������������������������������������   �4, E� B ��� ��@��@&��@���)��t���Ђ�������� �                                                                                                                                                                                                                                                                                                        H�	A'��                                                                                                                                                                                                                                 
    y    1      �  L�J                                     ������������������������������������������������������                                                                                                                                      �    L�              X          ��                 	 	 ���������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ����           �                     /    � �  E�J      z�  	                           ������������������������������������������������������                                                                    
                                                                    �    � R       6      ��       �    �          
 	    � ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� ������������������           h                                                                                                                                                                                                                                                 
                                        	                    �             


           �   }�         wwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwww A C 6                                 � ��[ �\                                                                                                                                                                                                                                                                                     
)nE  "h        k      e      k                  m            `                                                                                                                                                                                                                                                                                                                                                                                                         @ $  � ��  � ��  � (��  � #��  J`$  ���������Y����������N�����B���������������H                      ��           �   & AG� �  y   
              �                                                                                                                                                                                                                                                                                                                                      p I H   �                       !��                                                                                                                                                                                                                            Y   �� �~ ���      �� 4      ���������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ����� ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� ������������������             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    <      8     ��                       4     �   �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$    `d     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@       �      �     ��     �D   	������2�������� �l� �l  �� � l         ��   @���� � ��� �� � ��� �$ ^$         ��f       @     1,�����2��������      �f  �&  yf  y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "! ""! " ""  "!  "! " ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "! ""! " ""  "!  "! " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "! " ""  "!  " ! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                          "  "  ""  ��  ��  �� ��  ��  �  �  �� ���T���T���ED��EUI���  /   /�  �   �   � ����ˊ}m��v��ɧk�̚���ɘ���̻̊����������    "  "  �/ ��/ ��� ��  ��        �  �  �  �  ��   ��                  ������� ��                       �   �   �   DUH�DUT�UT��T���H�� �O  ��� ��                        E �EUEUT��DC��33��������  E   �  �  �� �� "��"/�"/ �/ ��� �      "   " � "� ""  / �� ��                        ��  ��  ��� �   ��  ���   �                 ���������������������  ��  ��  ��  �   �    �          �         �                                                                                                "  "  ""  +  �" � ��            "" ""  "  �/ ��         ̴E��EU��DU���D���� ��UEU ��Tʌˈ����+�� ����               U@� UT��DE��CU��5T��UT��T���������  �                                           � �� ������̊��̚w�̚v�̚w�̚��̹�˻˙��̻���� ��� ��  ��  �                    "  ".� "" �/���      g�  ��� }�� ��� ��� ��� �        "  ""  ""/ �"� ��          �   �  � �� ��  �                        �   ��  �   ��  ��  �  �  �   �                                 �   ���                            �   �                      ��   ��                  �  �  �� � ���                                  �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��� ���� ��    �     �                                                                                                                                                                                                  �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �   �                                    ��                                ��                      �����                                  �  �˰ ��� �wp ���                                                                                                                                                                                �    � � U  T  �Z  J  �  �  �� �� ��� ��� +�� �� �"   ��     �           �  ̚ �ɪ�̹�̻٪�����ټ̭��ˌ����ɣDH� T����ɀ�ɀ�����̘뚌���.� ������ � �          ��� ��� ��� ��  ��  �݀ �ؘ�ݍ��3�݉C���D���������  ��  �   �   �   �   /�  ��������    ����                        �  �˰ ���      � ��� ��� ��  �                �   �     �   �                                          �   �           �   ̰  �˰     �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                                  �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                �����                         �     �                                                                                                                                                                                   "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��             �  �˰ ��� �wp ���      � �������������  �                                                                                                                                           �  ��� ݻ� g�� bm� ggz�'w���������������˛������ˊۼ�����˻������H�DH�@U�DPT�E X�T H�P H�@ Ȥ� ̻� ˘ "�� � ���/�"" �""/���               �   �                                                     �  �                      � �                       ���           �                      �  �  �          ����  �   �             ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                                                                                                                                                                    �� ݻ� ��� �ww�}}m�wgg��wp��� ٪�"ܙ�"�̛���˰ۼ̰ۋɀ������           �  
�  �  �   �   �������C�
�DLJ�UCJ�UCJ�TCUTUT EC DL �� 
�� �� +� ""�"""�""����� ��     �        �  �" ��"� �"  3"  3U  4E  4�  ;�  ��  ��  ��  ""  ""  "" �"����� �                �    �    �     ��   �      �          �   �   �   �  �    �  �                      �   �   �  �    �   /   "�  "�  "�  ��                          �   O   T     ��                                 � ���� ��   � � �                            ����                  �   �� �       �  �  ��  �   �   �   �                                         �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��        �  �  �  �                 ���� �                                                                                                                                                                                             �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��                     �    � �  ��                  ���                                                                                                                                                                               ̘����	�������͹���۸�����̌�+���(����ی��ی�N=��NC��U �� 	�� �� ��  ��  ��  ��  �� �� �� ��"� �    �            ��  ��  ̽� �݋ �ݨ�����)*������˚���ɛ���̽ݩ��ݚ���ɚ،̴X��E���E������������������������ ��� ��� �����������" � � �      �   �   �   �   �   �   �                   �   �   �   �   �   �   �   �   �  ��  �     ��     �   �  ��  ��  �   �            �   �   �   �    �                             �          �                                                                                                                                                                                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""������������������""""������������������������""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""���������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��������������D�����3333DDDDI����D��DI����3333DDDDADAIA����D������3333DDDD��������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
� �Mc~ �O c� �]c� �l c� �V c� �N c� �*C(B	C"8 �
cjAcnA �cp) �cs! � cw9 cx( � � � � � � �cV& � c^& � c_6 �c`6 � cb. � cc+ �c�E � c�U � c�= � c�@ � c�F � c�H �c�5 � c�E �  c�- � !c�0 � "c�6 � #c�8 �$CB � � %CJ � �&"� � � '"� � �(� � �)
� � �*"� � � +"� � �,"� � �-*� �w."� �w /"� �g0� �g 
� � �2"�  � 3"�2 �4� � 
�' �6� � 
�' �8� � 
�' �:"P � ;*O� �  *H� � =*O� �  *H�@ *<t3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������$���.�U�[�M��1�O�R�S�U�[�X� � � � � � � � �=��;�����������������������������������������$��1�R�K�T�T��+�T�J�K�X�Y�U�T� � � � � � �=��;�������������������������������������������.�G�R�K��2�G�]�K�X�I�N�[�Q� � � � � � �,�>�0�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������=��;� ��!�������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������,�>�0� �� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                