GST@�                                                           �t�                                                      �   B                 
      ����e j�	 J�����������`�������        i      #    ����                                d8<n    �  ?     R�����  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"    B�j�
�  B ��
  �                                                                              ����������������������������������      ��    bbo QQ g 11 44             		� 

                      ��                      nn� ))         888�����������������������������������������������������������������������������������������������������������������������������o=  0  o4   1  +      '           �                    	�  7�  V�  	�                    
          : �����������������������������������������������������������������������������                                (,  ,   �  ��   @  #   �   �                                                                                'w w  )n)n�  
    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E , �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��bD� �S�
M$3�{�Y|8B�� <i�����R��3��T0 k� �s��w�e1�t B�1	�"q  ��" 
   ��� G��cD߆ �W�2�w�a�8B�� 8hQ����R��3��T0 k� �w��{�e1�t B�1	�"q  ��" 
   ��� H��eDׇ �[�2�s�a�8B�� 4hQ����R��3��T0 k� �w��{�e1�t B�1	�"q  ��" 
   ��� I��fDχ �_�2�o�a�8B�� 4gQ����R��3��T0 k� �����e1�t B�1	�"q  ��" 
   ��� J��gDÇ �c�2�o�a�8B�� 0fQ����R��3��T0 k� ������e1�t B�1	�"q  ��" 
   ��� K��iD�� �c�1�k�a�8B�� 0fQ���{�R��3��T0 k� ������e1�t B�1	�"q  ��" 
   ��� L��jD�� �g� 1�g�a�8B�� 0eQ���s�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� M�kD�� �k��1�c�a�8B�� ,dA���o�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� N�lD�� �o���0�c�a�8B�#� ,cA���g�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� O�nD�� �s���0�_�a�8B�#��,bA���c�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� P�oD�� �w���0�_�a�8B�'��,bA���[�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� Q�pD�� �{���/�[�a�8B�'��,aA�W�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� RѨqC�� ����/�[�Y|8B�+��(`A�S�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� SѤrC�w� �����.�[�Y|8B�/��,_1�K�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� TќsC�o�����.�W�Y|8B�3��,_1�G�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� UєuC�g�����-�W�Y|8B�3��,^1�C�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� VьvC�_�����-�W�Y|8B�7��,]1�?�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� WфwC�S�����,�S�Y|8B�;��,]1�;�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� X�|xC�K�����,�S�Y|8B�?��0\1�7�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� Z�tyC�C�����+�S�Y|8B�C��0[!�3�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� \�pzC�;�����+�O�Y|8B�G��0[!�/�R��3��T0 k� ������e1�t B�1	�"q  ��" 	   ��� ^�h{EA3�����+�O�Y|8B�K��4Z!�+����3��T0 k� ����ãe1�t B�1	�"q  ��" 	   ��� `�`|EA+�����*�O�Y|8B�O��4Y!��+����3��T0 k� �Ǥ�ˤe1�t B�1	�"q  ��" 	   ��� b�X}EA#�����*�K�a�8B�S��8Y!��'����3��T0 k� �ˤ�Ϥe1�t B�1	�"q  ��" 	   ��� d�P}EA�����)�K�a�8B�[��8Y���#����3��T0 k� �Ӥ�פe1�t B�1	�"q  ��" 	   ��� f�H~EA�Ǭ��)�K�a�8B�_��<X���#����3��T0 k� �ۥ�ߥe1�t B�1	�"q  ��" 	   ��� h�@EA�Ϭ��)�K�a�8B�c��@X�������3��T0 k� �ߦ��e1�t B�1	�"q  ��" 	   ��� j�8�E@��ӭ��(�G�a�8B�g��@X�������3��T0 k� ����e1�t B�1	�"q  ��"    ��� l�0E@���ۮ��(�G�a�8B�o��DW�������3��T0 k� ����e1�t B�1	�"q  ��"    ��� n�(E@�����'�G�a�8B�s��HW�������3��T0 k� ������e1�t B�1	�"q  ��"    ��� p� E@�����'�G�a�8B�w��HW�������3��T0 k� ������e1�t B�1	�"q  ��"    ��� r�~E@ۏ����'�C�a�8I��LW�������3��T0 k� ����e1�t B�1	�"q  ��"    ��� t�~E0ӏ�����&�C�a�8I���PW�������3��T0 k� ����e1�t B�1	�"q  ��"    ��� v�}E0ˏ�����&�C�a�8I���TW������3��T0 k� ����e1�t B�1	�"q  ��"    ��� x��}E0Ð����&�C�Y|8I���XW������3��T0 k� ����e1�t B�1	�"q  ��"    ��� z��|E0������%�?�Y|8I���\W������3��T0 k� �#��'�e1�t B�1	�"q  ��"    ��� |��|E0������%�?�Y|8I���\W������3��T0 k� �'��+�e1�t B�1	�"q  ��"    ��� ~��{E0������%�?�Y|8I �� `W���2��3��T0 k� �/��3�e1�t B�1	�"q  ��"    ��� ���zE0���#���$�?�Y|8I �� dX���2��3��T0 k� �7��;�e1�t B�1	�"q  ��"    ��� ���zE0���+���$�;�Y|8I �� hX���2��3��T0 k� �?��C�e1�t B�1	�"q  ��"    ��� ���yE0���3���$�;�Y|8I �� pX�
B�2��3��T0 k� �K��O�e1�t B�1	�"q  ��"    ��� ���xE0���;���#�;�Y|8I �� tX�
B�2��3��T0 k� �S��W�e1�t B�1	�"q  ��"    ��� ���wE0��G���#�;�Y|8I��xX��
B�2��3��T0 k� �[��_�e1�t B�1	�"q  ��"    ��� ��vE w��O���#�;�Y|8I��|Y��
B�2��3��T0 k� �c��g�e1�t B�1	�"q  ��"    ��� ��uE o��W���"�7�Y|8I���Y��
B�2��3��T0 k� �k��o�e1�t B�1	�"q  ��"    ��� ��tE g��_���"�7�Y|8I���Y��"�2��3��T0 k� �w��{�e1�t B�1	�"q  ��"    ��� � �sE _��g���"�7�Y|8I���Y��"�2��3��T0 k� ������e1�t B�1	�"q  ��"    ��� � �rE W��o��!�7�Y|8B����Y�"�2��"s��T0 k� ������e1�t B�1	�"q  ��"    ��� � �pE O��{��!�7�Y|8B����Y�"�2��"s��T0 k� ������e1�t B�1	�"q  ��"    ��� � �nE ?����� �7�Y|8B�ǥ��Z"�2����"s��T0 k� ������e1�t B�1	�"q  ��"    ��� � �mE ;����� �7�Y|8B�˥��Z"�2����"s��T0 k� ������e1�t B�1	�"q  ��"    ��� � �lE 3�������7�Y|8B�ϥ��Z"�2����"s��T0 k� ������e1�t B�1	�"q  ��"    ��� � �jE /�������7�Y|8B�ӥ��Z"�2����"s��T0 k� ������e1�t B�1	�"q  ��"    ��� � |iE'�������7�Y|8B�ۥ��Z"�2����"s��T0 k� ������e1�t B�1	�"q  ��"    ��� � xhE#�������7�Y|8B�ߥ��["�B����"s��T0 k� ������e1�t B�1	�"q  ��"    ��� � tfE��ú���7�Y|8B����[�B����"s��T0 k� ������e1�t B�1	�"q  ��"    ��� � peE��˻���;�Y|8B����[#�B����"s��T0 k� ������e1�t B�1	�"q  ��"    ��� � lcE��Ӽ���;�Y|8B����['�B����3��T0 k� ������e1�t B�1	�"q  ��"    ��� ��lbE��߽���;�Y|8B����[+�B����3��T0 k� ������e1�t B�1	�"q  ��"    ��� ��d_E��߽���?�Y|8B�����\;�2����3��T0 k� ������e1�t B�1	�"q  ��"    ��� ��d^B��������C�Y|8B����\?�2����3��T0 k� ������e1�t B�1	�"q  ��"    ��� ��`]B��������C�Y|8B����\G�2����3��T0 k� ������e1�t B�1	�"q  ��"    ��� ��`[B���������G�Y|8B���\O�2����3��T0 k� ������e1�t B�1	�"q  ��"    ��� ��\ZB���������K�Y|8B���\S�2����3��T0 k� ������e1�t B�1	�"q  ��"    ��� ��\YB��������K�Y|8B���\[�"#����3��T0 k� ������e1�t B�1	�"q  ��"    ��� ��\XB�������O�Y|8B�'�� \�c�"#����3��T0 k� ������e1�t B�1	�"q  �"    ��� ��XVB�������S�Y|8B�/��(]�k�"'����3��T0 k� ������e1�t B�1	�"q  ��"    ��� ��XUB�������S�Y|8B�3��0]�s�"'����"���T0 k� ������e1�t B�1	�"q  ��"    ��� ��XTB�������W�Y|8B�;��8]�w�"+����"���T0 k� ������e1�t B�1	�"q  ��"    ��� ��XSB�������[�Y|8EC��@]��/����"���T0 k� ������e1�t B�1	�"q  ��"    ��� ��XRB�������_�Y|8EK��H]���3����"���T0 k� �����e1�t B�1	�"q  ��"    ��� ��\OB�������g�Y|8E[��\]���;����"���T0 k� ����e1�t B�1	�"q  ��"    ��� ��\NB�������k�Y|8Ec��d]���?����"���T0 k� �����e1�t B�1	�"q  ��"    ��� ��\MB�������o�Y|8Eg��l^���2C����"���T0 k� ����e1�t B�1	�"q  ��"    ��� ��`LB�������s�Y|8E�o��t^���2G����"���T0 k� ����e1�t B�1	�"q  ��"    ��� ��`KB�������w�Y|8E�w���^���2K����"���T0 k� ����e1�t B�1	�"q  ��"    ��� ��dJB�������{�Y|8E����^���2K����"���T0 k� �����e1�t B�1	�"q  ��"    ��� ��dIB��������Y|8E�����^���2O����3��T0 k� �����e1�t B�1	�"q  ��"    ��� ��hHB������܃�Y|8E�����^���2S����3��T0 k� ����e1�t B�1	�"q  ��"    ��� ��hGB������܇�Y|8E�����^r��BW����3��T0 k� ����e1�t B�1	�"q  ��"    ��� ��lFB������܏�Y|8E�����^r��B[����3��T0 k� ����e1�t B�1	�"q  ��"    ��� ��pEB������ܓ�Y|8E���Ѵ^r��B_�B��3��T0 k� ����e1�t B�1	�"q  ��"    ��� ��tCB������ܛ�Y|8E�����_r��Bg�B��3��T0 k� ����e1�t B�1	�"q  ��"    ��� ��xBB������ܣ�Y|8D�è��_���Bk�B��3��T0 k� �����e1�t B�1	�"q  ��"    ��� ��|AB�������ܧ�Y|8D�˨��_���Bo�B��3��T0 k� �����e1�t B�1	�"q  ��"    ��� ���@B������ܯ�Y|8D�ө	�_��Bs�B��3��T0 k� �����e1�t B�1	�"q  ��"    ��� ���@B������ܳ�Y|8D�۩	�_��Rw� ��3��T0 k� �����e1�t B�1	�"q  ��"    ��� ���?B�����ܷ�Y|8D��	�_��R{� ��3��T0 k� ������e1�t B�1	�"q  ��"    ��� ���>B��������Y|8E��	�_s�R� ��3��T0 k� ������e1�t B�1	�"q  ��"    ��� ���=B����� �ýY|8E��	�_s#�R�� ��3��T0 k� ������e1�t B�1	�"q  ��"    ��� ���<B�����$�˽Y|8E���	"_s'�R�� ��3��T0 k� ������e1�t B�1	�"q  ��"    ��� ���;B�����,�ϽY|8E��	"_s/�ҋ� b��3��T0 k� ������e1�t B�1	�"q  ��"    ��� ���:B�����4�׽Y|8E��	"_s7�ғ� b��3��T0 k� �����e1�t B�1	�"q  ��"    ��� ���9B�#����D��Y|8E��	"_sC�қ� b��3��T0 k� ����e1�t B�1	�"q  ��"    ��� �д8B�'����L��Y|8E�'�	 _sG�ң� b��3��T0 k� ����e1�t B�1	�"q  ��" 	   ��� �и7B�/����T��Y|8E�/�	(_sO�§� b��3��T0 k� ����e1�t B�1	�"q  ��" 	   ��� ���7B�3����\���Y|8D�7�	,_sS�«� b��3��T0 k� ����e1�t B�1	�"q  ��" 	   ��� ���6B�;����d���Y|8D�?�	0_c[�³� ���3��T0 k� ����e1�t B�1	�"q  ��" 	   ��� ���5B�?���l��Y|8D�G�	4_c_�·� ���3��T0 k� ����e1�t B�1	�"q  ��" 	   ��� ���4B�G���t��Y|8D�O�	"<_cc�¿� ���3��T0 k� ���#�e1�t B�1	�"q  ��" 	   ��� ���4B�O���|��Y|8D�W�	"@_cg�
��� ���3��T0 k� �#��'�e1�t B�1	�"q  ��" 	   ��� ���3B�W������Y|8E�c�	"D_co�
��� ���3��T0 k� �#��'�e1�t B�1	�"q  ��" 	   ��� ���2B�_������#�Y|8E�k�	"H_cs�
���B��3��T0 k� �'��+�e1�t B�1	�"q  ��" 	   ��� ���1B�o������/�Y|8E�{�	"L_c{�
���B��3��T0 k� �+��/�e1�t B�1	�"q  ��" 	   ��� ���0B�w�������7�Y|8E���	P_c�
���B��3��T0 k� �'��+�e1�t B�1	�"q  ��" 	   ��� ��0B��������?�Y|8E���	T_c��
���B��3��T0 k� �#��'�e1�t B�1	�"q  ��" 	   ��� ��/B���������G�Y|8E���	X_c��
���B��3��T0 k� ���#�e1�t B�1	�"q  ��" 	   ��� ��.B���������O�Y|8E���	\_S��
���B��3��T0 k� ����e1�t B�1	�"q  ��" 	   ��� ��.B��������W�Y|8E���	\_S��
���B��3��T0 k� ���#�e1�t B�1	�"q  ��" 	   ��� ��$-B��������_�Y|8E���	"`_S��
���R��3��T0 k� ���#�e1�t B�1	�"q  ��" 	   ��� ��,,B��������g�Y|8BB��	"`_S��
��R��3��T0 k� ���#�e1�t B�1	�"q  ��" 	   ��� ��8,E�������o�Y|8BB��	"d_S��
��R��3��T0 k� �#��'�e1�t B�1	�"q  ��" 	   ��� ��@+E�������s�Y|8BB��	"d_S��
��R��3��T0 k� �#��'�e1�t B�1	�"q  ��" 	   ��� ��H+EØ�����{�Y|8BBǾ	"h_S��
��R��3��T0 k� �'��+�e1�t B�1	�"q  ��" 	   ��� ��P*E˘ r���̓�Y|8BBϿ	h_S��
��R��3��T0 k� �'��+�e1�t B�1	�"q  ��" 
   ��� ��X*Eט r�� ͋�Y|8BB��	l_S��'�R��3��T0 k� �+��/�e1�t B�1	�"q  ��" 
   ��� ��`)Eߘ r��͓�Y|8BB��	l_��+�R��3��T0 k� �+��/�e1�t B�1	�"q  ��" 
   ��� ��h(E� r��͛�Y|8BB��	l_��/�R��3��T0 k� �/��3�e1�t B�1	�"q  ��" 
   ��� ��p(E� r��ͣ�Y|8BB��	l_��3�R��3��T0 k� �3��7�e1�t B�1	�"q  ��" 
   ��� ��x'E����$ͫ�Y|8BB��	"p_㛿;�R��3��T0 k� �3��7�e1�t B�1	�"q  ��" 
   ��� ���'E����,ݳ�Y|8BB��	"p_㛾?�2��3��T0 k� �3��7�e1�t B�1	�"q  ��" 
   ��� ���&E����4ݻ�Y|8BB��	"p_㛾C�2��3��T0 k� �3��7�e1�t B�1	�"q  ��" 
   ��� ���&E��#��<�ûY|8BB��	"p_㛽G�2��3��T0 k� �7��;�e1�t B�1	�"q  ��" 
   ��� ���%E��'��D�ǻY|8BC�	"p_S��K�2��3��T0 k� �;��?�e1�t B�1	�"q  ��" 
   ��� ���%E�#��+��L�ϻY|8BC�	p_S��O�2��3��T0 k� �?��C�e1�t B�1	�"q  ��" 
   ��� ���$E�3��3��\�߻Y|8BC�	p_S��W�"��3��T0 k� �G��K�e1�t B�1	�"q  ��" 
   ��� ���#E�?��7��d��Y|8BC�	p_S��[�"��3��T0 k� �K��O�e1�t B�1	�"q  ��" 
   ��� ���#E�G��;��l��Y|8E��	p_S��_�"��3��T0 k� �O��S�e1�t B�1	�"q  ��" 
   ��� ���#E�O��?��t���Y|8E��Bp_S��_�"��3��T0 k� �S��W�e1�t B�1	�"q  ��" 
   ��� ���"E�W��C��|���Y|8E��Bp_S��c�"� c��T0 k� �W��[�e1�t B�1	�"q  ��" 
   ��� ���"D�_��G�ބ��Y|8E�#�Bp_S��c��c��T0 k� �[��_�e1�t B�1	�"q  ��" 
   ��� ���!D�g�rK�ސ��Y|8E�#�Bp_S��g��c��T0 k� �_��c�e1�t B�1	�"q  ��" 
   ��� ���!D�s�rS�ޘ��Y|8Es'�Bp_ㇷk��c��T0 k� �c��g�e1�t B�1	�"q  ��" 
   ��� ��� D�{�rW�ޠ��Y|8Es+�Bp_ヶk��c��T0 k� �g��k�e1�t B�1	�"q  ��" 
   ��� ��  Dу�r[�ި�#�Y|8Es+�Bp_ヵo��c��T0 k� �k��o�e1�t B�1	�"q  ��" 
   ��� ��Dѓ�rc�޸�3�Y|8Es/�Bp_�{�s��c��T0 k� �s��w�e1�t B�1	�"q  ��" 
   ��� ��Dћ�rg����;�Y|8Es3�Bp_�w�s��	c��T0 k� �w��{�e1�t B�1	�"q  ��" 
   ��� �� Dѣ�rk����C�Y|8Es7�Bp_�s�w��
c��T0 k� �{���e1�t B�1	�"q  ��"    ��� ��(Dѯ�ro����K�Y|8Es;�Bp_�s�w��c��T0 k� �����e1�t B�1	�"q  ��"    ��� ��0Dѷ�rs����S�Y|8Ec;��p_�o�{���c��T0 k� ������e1�t B�1	�"q  ��"    ��� ��8Dѿ�rw����[�Y|8Ec?��p_�k�{���c��T0 k� ������e1�t B�1	�"q  ��"    ��� ��@D�Ǡr{����_�Y|8EcC��p_�g�{���c��T0 k� ������e1�t B�1	�"q  ��"    ��� ��HD�Ϡb����g�Y|8EcC��p_�c��� c��T0 k� �����e1�t B�1	�"q  ��"    ��� ��TD�סb�����o�Y|8EcG��p_�[���c��T0 k� �w��{�e1�t B�1	�"q  ��"    ��� ��\D��b����w�Y|8EcG��p_�W���c��T0 k� �s��w�e1�t B�1	�"q  ��"    ��� ��lE��b������Y|8EcK��p_�O���c��T0 k� �s��w�e1�t B�1	�"q  ��"    ��� ��tE����������Y|8EcO��p_�K���c��T0 k� �o��s�e1�t B�1	�"q  ��"    ��� ��|E������$���Y|8EcO��p_�C����c��T0 k� �o��s�e1�t B�1	�"q  ��"    ��� ���E������,���Y|8ESO��p_�?����c��T0 k� �k��o�e1�t B�1	�"q  ��"    ��� ���E������4���Y|8ESO��p_�;���� c��T0 k� �k��o�e1�t B�1	�"q  ��"    ��� ��E������<���Y|8ESS��p_�3�
����$c��T0 k� �k��o�e1�t B�1	�"q  ��"    ��� ��E�'�b���Dγ�Y|8ESS��p_�/�
����(c��T0 k� �k��o�e1�t B�1	�"q  ��"    ��� ��E�7�b���T�ùY|8ESS��p_�#�
����0c��T0 k� �k��o�e1�t B�1	�"q  ��"    ��� ��E�?�b���\�˹Y|8ESS��p_�
����4c��T0 k� �o��s�e1�t B�1	�"q  ��"    ��� ���E�G�b���h�ӹY|8ESO��p_�
����8c��T0 k� �o��s�e1�t B�1	�"q  ��"    ��� ���ErS�b���p�۹Y|8ESO��p_�
����@c��T0 k� �o��s�e1�t B�1	�"q  ��"    ��� ���Er[�b���x��Y|8ESO��p_�
Ӄ��Dc��T0 k� �o��s�e1�t B�1	�"q  ��"    ��� ��Er[�b����
��Y|8ECO��p_�
Ӄ��Hc��T0 k� �o��s�e1�t B�1	�"q  ��"    ��� ��Er_�R����
��Y|8ECK��p_��
Ӄ��Lc��T0 k� �s��w�e1�t B�1	�"q  �"    ��� ��Erc�R����
���Y|8ECK��p_��
Ӄ��Xc��T0 k� �{���e1�t B�1	�"q  ��/    ��� ��Erc�R��Ϡ
��Y|8ECG��p_��
Ӄ��\c��T0 k� ������e1�t B�1	�"q  ��/    ��� ��Erc�R��Ϩ
��Y|8ECG��p_��
Ӄ��`c��T0 k� ������e1�t B�1	�"q  ��/    ��� ��Ebc���ϰ
��Y|8ECC��p_R�
Ӄ�shc��T0 k� ������e1�t B�1	�"q  ��/    ��� ��Ebc���ϸ
��Y|8ECC��p_Rߧ
Ӄ�slc��T0 k� ������e1�t B�1	�"q  ��/    ��� �� Ebc�����
�'�Y|8E3?��p_Rߦ
Ӄ�spc��T0 k� ������e1�t B�1	�"q  ��/    ��� ��(Ebc�����
�/�Y|8E3?��p_Rۦ
Ӄ�stc��T0 k� ������e1�t B�1	�"q  ��/    ��� ��0Ebc�����
�7�Y|8E3;��p_Rצ
Ӄ�sxc��T0 k� ������e1�t B�1	�"q  ��/    ��� ��8D2c�"����
�?�Y|8E3;��p_Rץ��s�c��T0 k� ������e1�t B�1	�"q  ��/    ��� ��@D2c�"����
�G�Y|8E37��p_Rӥ��s�c��T0 k� ������e1�t B�1	�"q  ��/    ��� ��HD2c�"����
�O�Y|8E37��p_Rӥ��s�c��T0 k� ������e1�t B�1	�"q  ��/    ��� ��P D2c�"����
�S�Y|8E33��p_RϤ��s�c��T0 k� ������e1�t B�1	�"q  ��/    ��� ��`!D2c�"���
�c�Y|8E3/��p_Rˤ3�s�c��T0 k� ������e1�t B�1	�"q  ��/    ��� ��h"D2c�"���
�k�Y|8E3/��p_Rǣ3�c�c��T0 k� ������e1�t B�1	�"q  ��/    ��� ��p"D2c�2���	�s�Y|8CC+��p_Rǣ3�c�c��T0 k� ������e1�t B�1	�"q  ��/    ��� ��x#DBc�2���	�{�Y|8CC+��p_Rã3�c�c��T0 k� ����Àe1�t B�1	�"q  ��/    ��� ���$DBc�2���$	���Y|8CC'��p_Râ3�c�c��T0 k� ��~��~e1�t B�1	�"q  ��/    ��� ���%DBc�2���,	���Y|8CC'��p_R��3{�c�c��T0 k� ��}��}e1�t B�1	�"q  *�/    ��� ���&DBc�2���4	���Y|8CC'��p_R��3{�c�c��T0 k� ��}��}e1�t B�1	�"q  ��/    ��� ���'DBc�2���<	���Y|8@�#��p_R��3{�c�c��T0 k� ��~��~e1�t B�1	�"q  ��/    ��� �Ü(DBc�2���D	��Y|8@�#��p_R���w�c�c��T0 k� ��~��~e1�t B�1	�"q  ��/    ��� �ä)A�c�2���P	��Y|8@���p_R���w�c�c��T0 k� ��~��~e1�t B�1	�"q  ��/    ��� �è*A�c�2���X	��Y|8@���p_R���s�S�c��T0 k� ����e1�t B�1	�"q  ��/    ��� �ð,A�c�2���`	��Y|8@���p_R���s�S�c��T0 k� ����e1�t B�1	�"q  ��/    ��� �ô-A�c�2��h	��Y|8@���p_R���s�S�
c��T0 k� ����e1�t B�1	�"q  ��/    ��� �ü.A�c�2��p	�ǸY|8@���p_R���o�S�	c��T0 k� ����e1�t B�1	�"q  ��/    ��� ���/BBc�2��x	�ϸY|8@���p_R���o�S�c��T0 k� ����e1�t B�1	�"q  ��/    ��� ���0BBc�2{���	�׸Y|8@���p_R���o��c��T0 k� �����e1�t B�1	�"q  ��/    ��� ���2BBc�2{���	�߸Y|8@���p_R���k���c��T0 k� ������e1�t B�1	�"q  ��/    ��� ���3BBc�2{���	��Y|8@���p_R���k���c��T0 k� ������e1�t B�1	�"q  ��/    ��� ���4BBc�2w���	��Y|8@���p_B��ck���c��T0 k� �����e1�t B�1	�"q  ��/    ��� ���5@c�2w���	��Y|8@���p_B��cg���c��T0 k� ����e1�t B�1	�"q  ��/    ��� ���7@c�2w���	���Y|8@���p_B��cg���c��T0 k� ����e1�t B�1	�"q  ��/    ��� ���8@c�2s���	��Y|8@���p_B��cg���c��T0 k� ����e1�t B�1	�"q  ��/    ��� ���9@c�2s���	��Y|8@���p_B��cc���c��T0 k� ����e1�t B�1	�"q  ��/    ��� ���:@c�2s���	��Y|8@���p_���cc���c��T0 k� ����e1�t B�1	�"q  ��    ��� ��;B�c�2s���	��Y|8@���p_���c_���c��T0 k� ����e1�t B�1	�"q  ��    ��� ��=B�c�2o���	�#�Y|8@���p_���c[���c��T0 k� ����e1�t B�1	�"q  ��    ��� ��>B�g�2o����'�Y|8@���p_���c[��c��T0 k� ���#�e1�t B�1	�"q  ��    ��� ��?B�g�2o����/�Y|8@���p_���cW�� c��T0 k� ���#�e1�t B�1	�"q  ��    ��� ��@B�g�2o����7�Y|8@���p_����W�S�����T0 k� �#��'�e1�t B�1	�"q  ��    ��� ��AB�g�2k����?�Y|8E3��p_����S�S�����T0 k� �'��+�e1�t B�1	�"q  ��    ��� ��CB�g�2k��O�Y|8E3��p_����O�S�����T0 k� �/��3�e1�t B�1	�"q  ��    ��� ��DB�g�2g�	�W�a�8E3��p_����K�S�����T0 k� �3��7�e1�t B�1	�"q  ��    ��� ��ECg�2g�	�[�a�8E2���p_����K�C�����T0 k� �7��;�e1�t B�1	�"q  ��    ��� ��FCg�2g�	�c�a�8E"���p_����G�C�����T0 k� �;��?�e1�t B�1	�"q  ��    ��� ��GCk�2g�	$�k�a�8E"���p_����C�C�����T0 k� �?��C�e1�t B�1	�"q  ��    ��� ��HCk�2g�	(�s�a�8E"���p_����C�C�����T0 k� �C��G�e1�t B�1	�"q  ��    ��� ���ICk�2c�	0�{�a�8E"���p_���?�C�����T0 k� �K��O�e1�t B�1	�"q  ��    ��� ���KCo�2c�	!<���a�8E"���p_�{��;�������T0 k� �G��K�e1�t B�1	�"q  ��    ��� ���LCo�2c�	!D���a�8E����p_�{��;�������T0 k� �G��K�e1�t B�1	�"q  ��    ��� ���MCo�2_�	!H���a�8E����p_�w�7�������T0 k� �K��O�e1�t B�1	�"q  ��    ��� ���NCs�2_�	!P���a�8E����p_�w�7�������T0 k� �S��W�e1�t B�1	�"q  ��    ��� ���OCs�2_�	!T���Y|8E����p_�w�3�������T0 k� �S��W�e1�t B�1	�"q  ��    ��� ���PCs�2_�	X���Y|8E����p_�w�3�ӓ����T0 k� �W��[�e1�t B�1	�"q  ��    ��� ���PCs�2_�	`���Y|8E����p_�w�3�ӏ����T0 k� �[��_�e1�t B�1	�"q  ��    ��� ���QCs�2[�	d���Y|8E����p_�w�/�Ӌ����T0 k� �[��_�e1�t B�1	�"q  ��    ��� ���SCs�2[�	l�ǨY|8E����p_�w�/�Ӄ����T0 k� �[��_�e1�t B�1	�"q  ��    ��� ���TCs�2[�	!p�ϧY|8E����p_�s�/������T0 k� �[��_�e1�t B�1	�"q  ��    ��� ���UCw�2[�	!t�צY|8E����p_�o�/��{����T0 k� �[��_�e1�t B�1	�"q  ��    ��� ���UCw�2W�	!xpߦY|8E����p_Bk�/��w����T0 k� �[~�_~e1�t B�1	�"q  ��    ��� ���VC{�2W�	!|p�Y|8E����p_Bg��/��s����T0 k� �W��[�e1�t B�1	�"q  �    ��� �S�WC�2W�	!�p�Y|8EB���p_Bc��/��o����T0 k� �S��W�e1�t B�1	�"q  �    ��� �S�XC��2W� �p�a�8EB���p_B_��/��k����T0 k� �O��S�e1�t B�1	�"q  ��    ��� �S�YC"��2S� �p��a�8EB���p^2W��/�	sc����T0 k� �K��O�e1�t B�1	�"q  ��    ��� �S�ZC"��2S� �q�a�8EB���p^2S��3�	s_����T0 k� �K��O�e1�t B�1	�"q  ��    ��� �S�[C"��2S� �q�a�8EB���p^2O��3�	s[����T0 k� �O��S�e1�t B�1	�"q  ��    ��� �S�[C"��2S� �q�a�8EB���p^2O��3�	sW����T0 k� �O�Se1�t B�1	�"q  ��    ��� �S�\C"��2S� �q�a�8EB���p]2K��7�	sS����T0 k� �S~�W~e1�t B�1	�"q  ��    ��� �S�]C"��2S� ���a�8E2���p]2G��7�	�S����T0 k� �S�We1�t B�1	�"q  ��   ��� �S�]E���2O� ��#�a�8E2���p\"C��;�	�O����T0 k� �W�[e1�t B�1	�"q  ��    ��� �S�^E���2O� ��'�a�8E2���p\"?��;�	�K����T0 k� �W��[�e1�t B�1	�"q  ��    ��� �S�_E���2O� ��/�a�8E2���p["?��?�	�K����T0 k� �[��_�e1�t B�1	�"q  ��    ��� �S�_E���2O� ��3�Y|8E2���pZ";��?�	�G����T0 k� �[��_�e1�t B�1	�"q  ��    ��� �S�`E���2O� ��;�Y|8E2���pZ"7��C�	sG����T0 k� �_��c�e1�t B�1	�"q  ��    ��� �S�aE���2O� ��?�Y|8E2���pY"7��G�	sC����T0 k� �c��g�e1�t B�1	�"q  ��    ��� �S�aE���2K� ��C�Y|8E2���pX"3��G�	sC����T0 k� �c��g�e1�t B�1	�"q  ��    ��� �S�bE���2K� ��K�Y|8E2���pW3��K�	s?����T0 k� �g��k�e1�t B�1	�"q  ��    ��� �S�bE�ã2K� ��O�Y|8E2��pV/��O�	s?����T0 k� �_��c�e1�t B�1	�"q  ��    ��� �S�cE�ˢ2K� ��S�Y|8E2��pU/��S�	�?����T0 k� �[��_�e1�t B�1	�"q  ��    ��� �S|dB�ϡ2K� ��[�Y|8E"��pT/��S�	�?����T0 k� �S��W�e1�t B�1	�"q  ��   ��� �SxeB�۟2K� ��c�Y|8E"ǽpR+��[�	�;����T0 k� �W��[�e1�t B�1	�"q  ��    ��� �SteB�ߞ2K� ��g�Y|8E"û�tQ+��[�	�;����T0 k� �S��W�e1�t B�1	�"q  ��    ��� �StfB��2G� ��k�Y|8E"ú�tP+��_�	s;����T0 k� �S��W�e1�t B�1	�"q  ��   ��� �SpfB��2G� ��s�Y|8K����tO+��c�	s;����T0 k� �W��[�e1�t B�1	�"q  ��    ��� �SlgB��2G� ��w�Y|8K����xN�+��c�	s;����T0 k� �W��[�e1�t B�1	�"q  ��    ��� �SlhB���2G� ��{�Y|8K����xM�/��g�	s;����T0 k� �[��_�e1�t B�1	�"q  ��    ��� �ShhB��2G� ���Y|8K����|L�/��k�	s;����T0 k� �[��_�e1�t B�1	�"q  ��    ��� �SdiB��2G� ��Y|8K����|K�/��k�S7����T0 k� �W��[�e1�t B�1	�"q  ��    ��� �SdiB��2G� ��Y|8K����|I�/��o�S7����T0 k� �[��_�e1�t B�1	�"q  ��    ��� �S`jB�#�2G� ��Y|8K���ҀH�3��o�S7����T0 k� �[��_�e1�t B�1	�"q  ��    ��� �S\jB�+�2C� ��Y|8K���҄G�3��s�S7����T0 k� �_��c�e1�t B�1	�"q  ��    ��� �S\kB�7�2C� ��Y|8K���҄E�7��s�S7����T0 k� �_��c�e1�t B�1	�"q  ��    ��� �SXkB�?�2C� ��Y|8K���҈D�7��s��7����T0 k� �_��c�e1�t B�1	�"q  ��    ��� �STlB�G�2C� ��Y|8K����C�;��s��7����T0 k� �_��c�e1�t B�1	�"q  ��    ��� �STlB�O�2C� ��Y|8K����A�;��w��7����T0 k� �_��c�e1�t B�1	�"q  ��    ��� �SPlB�[�2C� ��Y|8K¯��@�?�w��7����T0 k� �W��[�e1�t B�1	�"q  ��    ��� �SPmB�c�2C� ��Y|8K¯��?�?�w��7����T0 k� �O��S�e1�t B�1	�"q  ��    ��� �SLmB�k�2C� ��Y|8K«��=�C�w��7����T0 k� �K��O�e1�t B�1	�"q  ��    ��� �SLnB�s�2C� ��Y|8K«��<�G�w��3����T0 k� �G��K�e1�t B�1	�"q  ��    ��� �SHnB�{�2?� ��Y|8K«��:�K�w��3����T0 k� �C��G�e1�t B�1	�"q  ��    ��� �SHoBデ2?� ��Y|8K§��9�O�w��3����T0 k� �?��C�e1�t B�1	�"q  ��    ��� �SDoB㋇2?� ��Y|8K§��7�S��w��3����T0 k� �G��K�e1�t B�1	�"q  ��    ��� �S@oB㓈2?� ��Y|8K§��6�W��w��3����T0 k� �K��O�e1�t B�1	�"q  ��    ��� �S@pB㛈2?� ��ËY|8K§��4�[��w��3����T0 k� �O��S�e1�t B�1	�"q  ��    ��� �S<pB㣈2?� ��ǋY|8K£��3�_��w��3����T0 k� �S��W�e1�t B�1	�"q  ��    ��� �S<qB㫉2?� ��ǋY|8K£��1�c��s��3����T0 k� �S��W�e1�t B�1	�"q  ��    ��� �S8qB㳉2?� ��ˊY|8K£��0�g��s��3����T0 k� �S��W�e1�t B�1	�"q  ��    ��� �S8qB㻊2?� ��ϊY|8K��.�k��s��3����T0 k� �S��W�e1�t B�1	�"q  ��    ��� �S8rB�Ê2?�  �ӊY|8K���,�o��s��3����T0 k� �S��W�e1�t B�1	�"q  ��    ��� �S4rB�ǊB?�  �׉Y|8K�r�+�s��o��3����T0 k� �O��S�e1�t B�1	�"q  ��    ��� �S4rB�ϋB;� �׉Y|8K�r�)�{��o��3����T0 k� �O��S�e1�t B�1	�"q  ��    ��� �S0sE#׋B;� �ۉY|8K�r�'���k��3����T0 k� �K��O�e1�t B�1	�"q  ��    ��� �S0sE#ߋB;� �߈Y|8K�r�%��k��3����T0 k� �K��O�e1�t B�1	�"q  ��    ��� �S,tE#�B;� ��Y|8K�r�#��g��3����T0 k� �G��K�e1�t B�1	�"q  ��    ��� �S,tE#�B;� ��Y|8K�r�"��g��3����T0 k� �G��K�e1�t B�1	�"q  ��   ��� �S(tE#�B;� ��Y|8K�r� �cc��3����T0 k� �7��;�e1�t B�1	�"q  ��    ��� �S(uE#��B;� ��Y|8K�r��c_�3����T0 k� �'��+�e1�t B�1	�"q  ��    ��� �S(uE$�B;� ��Y|8K����c_�3����T0 k� ���#�e1�t B�1	�"q  ��    ��� �S$uE$�R;� ��Y|8K���ҧ�c[�3����T0 k� ����e1�t B�1	�"q  ��    ��� �S vE$�R;� ���Y|8K���ҳ�cS�7����T0 k� ����e1�t B�1	�"q  ��    ��� �S vE�R;� ���Y|8K���һ�cO��7����T0 k� ����e1�t B�1	�"q  ��    ��� �S vE�R;� ���Y|8K��ҿ�cK��7����T0 k� ������e1�t B�1	�"q  ��    ��� �SwE'�R;� ���Y|8K��ǼsG��7����T0 k� ������e1�t B�1	�"q  ��    ��� �SwE+�R;� ���Y|8K� ϼsC��;����T0 k� ������e1�t B�1	�"q  ��    ��� �SwE3�R?� ���Y|8K�׽s?��;����T0 k� ������e1�t B�1	�"q  ��    ��� �SxE7�R?� ���Y|8K�
۽s;��?����T0 k� ������e1�t B�1	�"q  ��    ��� �SxE?�R?� ��Y|8K��s7��?����T0 k� ������e1�t B�1	�"q  ��    ��� �SxEC�RC� ��Y|8K��s3��C����T0 k� ������e1�t B�1	�"q  $�    ��� �SxEK�RC�  ��Y|8K��s+��C����T0 k� ������e1�t B�1	�"q  ��    ��� �SyEW�RG�  ��Y|8K�� ��s'��G����T0 k� ������e1�t B�1	�"q  ��    ��� �Sy@[�RG� $��Y|8K��#���s#��K����T0 k� ������e1�t B�1	�"q  ��    ��� �Sy@_�RG� $��Y|8K��'���s��K����T0 k� ������e1�t B�1	�"q  ��    ��� �Sz@_�RG� $��Y|8K��+������O����T0 k� ������e1�t B�1	�"q  ��    ��� �Sz@_�RK� (��Y|8K��/������S����T0 k� ������e1�t B�1	�"q  ��    ��� �Sz@_�RK� (��Y|8K���s3�������S����T0 k� ������e1�t B�1	�"q  ��    ��� �Sz@_�RK� (��Y|8K���s7�������W����T0 k� ������e1�t B�1	�"q  ��    ��� �S{@_�RK� (��Y|8K���s;�������[����T0 k� ������e1�t B�1	�"q  ��    ��� �S{@_�RO� ,��Y|8K���s?�������_����T0 k� ������e1�t B�1	�"q  ��    ��� �S{@c�RO� ,��Y|8K���sC��������_����T0 k� ������e1�t B�1	�"q  ��    ��� �S{@c�RO� ,��Y|8K���sG��������c����T0 k� ������e1�t B�1	�"q  ��    ��� �S|@c�RO� 0��Y|8@b���K��������g����T0 k� ������e1�t B�1	�"q  ��    ��� �S|@c�RS� 0��Y|8@b���K��������k����T0 k� ������e1�t B�1	�"q  ��    ��� �S|@c�RS� 0��Y|8@b���O����R���o�"���T0 k� ������e1�t B�1	�"q  ��    ��� �S |@c�RS� 0��Y|8@b���S����R���s�"���T0 k� ������e1�t B�1	�"q  ��   ��� �S }@_�RS� 4��Y|8@b���W����R���w�"���T0 k� ������e1�t B�1	�"q  ��    ��� �S }@_�RS� 4��Y|8B���[����R���{�"���T0 k� ������e1�t B�1	�"q  ��    ��� �S }@_�RW� 4��Y|8B���_����R���{�"���T0 k� ������e1�t B�1	�"q  ��    ��� �R�}@_�RW� 4��Y|8B���c����R����"���T0 k� ������e1�t B�1	�"q  ��    ��� �R�}@_�RW� 8��Y|8B���g����R����"���T0 k� ������e1�t B�1	�"q  ��    ��� �R�~@_�RW� 8��Y|8B���k����R����"���T0 k� �����e1�t B�1	�"q  ��   ��� �R�~@_�R[� 8��Y|8B���o���R����"���T0 k� �w��{�e1�t B�1	�"q  ��    ��� �R�~@[�R[� 8��Y|8B����s���R����"���T0 k� �s��w�e1�t B�1	�"q  ��    ��� �R�~@[�R[� 8��Y|8B����w���R����"���T0 k� �o��s�e1�t B�1	�"q  ��    ��� �R�~@[�R[� <��Y|8B����{���R�������T0 k� �k��o�e1�t B�1	�"q  ��    ��� �R�@[�R[� <��Y|8K�������R��s�����T0 k� �g��k�e1�t B�1	�"q  ��    ��� �R�@W�R[� <��Y|8K���Ӄ���R��s�����T0 k� �c��g�e1�t B�1	�"q  ��    ��� �R�@W�R_� <��Y|8K���s����R��s�����T0 k� �_��c�e1�t B�1	�"q  ��    ��� �R�@W�R_� @�#�Y|8K���s����R��s�����T0 k� �[��_�e1�t B�1	�"q  ��    ��� �R�@S�R_� @�#�Y|8K���s����R��s�����T0 k� �W��[�e1�t B�1	�"q  ��    ��� �R�@S�R_� @�#�Y|8K���s������s�����T0 k� �c��g�e1�t B�1	�"q  ��    ��� �R��@S�R_� @�#�Y|8K���s������s�����T0 k� �k��o�e1�t B�1	�"q  ��    ��� �R�@S�Rc� @�#�Y|8K���s������s�����T0 k� �s��w�e1�t B�1	�"q  ��    ��� �R�@S�Rc� @�'�Y|8K���s������s�����T0 k� �w��{�e1�t B�1	�"q  ��    ��� �R�@O�Rc� D�'�Y|8K����������s�����T0 k� �w��{�e1�t B�1	�"q  ��    ��� �R�@O�Rc� D�'�Y|8K����������së"���T0 k� �w��{�e1�t B�1	�"q  ��    ��� �R�~@O�Rc� D�'�Y|8K����������sǩ"���T0 k� �w��{�e1�t B�1	�"q  ��   ��� �R�~@O�Rc� D�'�Y|8K����������s˨"���T0 k� �w��{�e1�t B�1	�"q  ��    ��� �R�~@K�Rg� D�'�Y|8K���������sϦ"���T0 k� �s��w�e1�t B�1	�"q  ��    ��� �R�~@K�Rg� H�+�Y|8K���	ӫ���{��ӥ"���T0 k� �o��s�e1�t B�1	�"q  ��    ��� �R�}@K�Rg� H�+�Y|8K���	ӫ���{��פ"���T0 k� �o��s�e1�t B�1	�"q  ��    ��� �R�}@K�Rg� H�+�Y|8K���	ӯ���w��ۢ"���T0 k� �o��s�e1�t B�1	�"q  ��    ��� �R�}@K�Rg� H�+�Y|8K���	ӯ���s��ߡ"���T0 k� �k��o�e1�t B�1	�"q  ��    ��� �R�}@G�Rg� H�+�Y|8K���	ӯ���o��ߠ"���T0 k� �g��k�e1�t B�1	�"q  ��    ��� �R�}@G�Rg� H�+�Y|8K���	㳱��"k���"���T0 k� �c��g�e1�t B�1	�"q  ��    ��� �R�|@G�Rk� L�+�Y|8K���	㳰��"k���"���T0 k� �_��c�e1�t B�1	�"q  ��    ��� �R�|@G�Rk� L�/�Y|8K���	㳯��"g������T0 k� �_��c�e1�t B�1	�"q  ��    ��� �R�|@G�Rk� L�/�Y|8K���	㷮��"g������T0 k� �[��_�e1�t B�1	�"q  ��    ��� �R�|@C�Rk� L	�/�Y|8K���	㷭��"g������T0 k� �[��_�e1�t B�1	�"q  ��    ��� �R�|@C�Rk� L	�/�Y|8K���S����"c������T0 k� �[��_�e1�t B�1	�"q  ��    ��� �R�{@C�Rk� L
�/�Y|8K���S����"c�������T0 k� �W��[�e1�t B�1	�"q  ��    ��� �R�{@C�Rk� L
�/�Y|8K���S����"_�������T0 k� �W��[�e1�t B�1	�"q  ��    ��� �R�{@C�Rk� L
�/�Y|8K���S����"_�������T0 k� �S��W�e1�t B�1	�"q  ��    ��� �R�{@?�Ro� L�3�Y|8K���S����"[�������T0 k� �S��W�e1�t B�1	�"q  ��    ��� �R�{@?�Ro� L�3�Y|8K���S����"[������T0 k� �O��S�e1�t B�1	�"q  ��    ��� �R�z@?�Ro� L�3�Y|8K�ÊS����"W������T0 k� �O��S�e1�t B�1	�"q  ��    ��� �R�z@?�Ro� L�3�Y|8K�ÊS����"W������T0 k� �O��S�e1�t B�1	�"q  ��    ��� �R�z@?�Ro� L�3�Y|8K�ÊS����"S������T0 k� �K��O�e1�t B�1	�"q  ��    ��� �R�z@?�Ro� L�3�Y|8K�ǊSã��"S������T0 k� �K��O�e1�t B�1	�"q  ��    ��� �R�z@;�Ro� L�3�Y|8K�Ǌcâ��"S������T0 k� �G��K�e1�t B�1	�"q  ��    ��� �R�z@;�Ro� L�3�Y|8K�Ǌcá��"O������T0 k� �G��K�e1�t B�1	�"q  ��    ��� �R�y@;�Rs� L�7�Y|8K�ˊcáC�"O������T0 k� �C��G�e1�t B�1	�"q  ��    ��� �R�y@;�Rs� L�7�Y|8K�ˋcǠC�"K������T0 k� �C��G�e1�t B�1	�"q  ��    ��� �R�y@;�Rs� L�7�Y|8K�ˋcǟC�"K������T0 k� �C��G�e1�t B�1	�"q  ��    ��� �R�y@;�Rs� L�7�Y|8K�ˋcǞC�"K������T0 k� �?��C�e1�t B�1	�"q  ��    ��� �R�y@;�Rs� L�7�Y|8K�ϋcǝC�"G������T0 k� �?��C�e1�t B�1	�"q  ��   ��� �R�y@7�Rs� L�7�Y|8K�ϋcǝ��"G������T0 k� �?��C�e1�t B�1	�"q  ��    ��� �R�y@7�Rs� L�7�Y|8K�ϋc˜��"C������T0 k� �;��?�e1�t B�1	�"q  ��    ��� �R�x@7�Rs� L�7�Y|8K�Ӌc˛��"C������T0 k� �;��?�e1�t B�1	�"q  ��   ��� �R�x@7�Rs� L�7�Y|8K�Ӌc˚��"C������T0 k� �7��;�e1�t B�1	�"q  ��    ��� �R�x@7�Rs� L�;�Y|8K�ӌc˚��"?������T0 k� �7��;�e1�t B�1	�"q  ��    ��� �R�x@7�Rw� L�;�Y|8K�ӌcϙ�#�"?������T0 k� �7��;�e1�t B�1	�"q  ��    ��� �R�x@7�Rw� L�;�Y|8K�׌cϘ�#�"?������T0 k� �3��7�e1�t B�1	�"q  ��    ��� �R�x@3�Rw� L�;�Y|8K�׌cϗ�'�";������T0 k� �3��7�e1�t B�1	�"q  ��   ��� �R�x@3�Rw� L�;�Y|8K�׌cϖ�+�";������T0 k� �/��3�e1�t B�1	�"q  ��    ��� �R�w@3�Rw� L�;�Y|8K�یcӕ�/�"7������T0 k� �/��3�e1�t B�1	�"q  ��    ��� �R�w@3�Rw� L�;�Y|8K�یcӕ�/�"7������T0 k� �/��3�e1�t B�1	�"q  ��    ��� �R�w@3�Rw� L�;�Y|8K�یcӔ�3�"7������T0 k� �+��/�e1�t B�1	�"q  ��    ��� �R�w@3�Rw� L�;�Y|8K�یcӓ�7�"7������T0 k� �+��/�e1�t B�1	�"q  ��    ��� �R�w@3�Rw� L�?�Y|8K�ۍcӓ�7�"3�t����T0 k� �+��/�e1�t B�1	�"q  ��    ��� �R�w@3�R{� L�?�Y|8K�ߍcӒ�;�"3�t����T0 k� �+��/�e1�t B�1	�"q  ��    ��� �R�w@3�R{� L�?�Y|8K�ߍcג�?�"3�t����T0 k� �'��+�e1�t B�1	�"q  ��    ��� �R�w@3�R{� L�?�Y|8K�ߍcב�C�", t����T0 k� �'��+�e1�t B�1	�"q  ��    ��� �R�v@/�R{� L�?�Y|8K�ߍcא�G�", t����T0 k� �'��+�e1�t B�1	�"q  ��    ��� �R�v@/�R{� L�?�Y|8K��cא�K�, t����T0 k� �  �$ e1�t B�1	�"q  ��    ��� �R�v@/�R{� L�?�Y|8B��c׏�O�( t����T0 k� �  �$ e1�t B�1	�"q  ��    ��� �R�v@/�R{� L�?�Y|8B��c׏�O�( t����T0 k� �  �$ e1�t B�1	�"q  ��    ��� �R�v@/�R{� L�?�Y|8B��c׏�S�( t����T0 k� �  �$ e1�t B�1	�"q  ��   ��� �R�v@/�R{� L�?�Y|8B��c׏�W�( t����T0 k� � �  e1�t B�1	�"q  ��    ��� �R�v@/�R{� L�?�Y|8B��c׎�[�$t����T0 k� � �  e1�t B�1	�"q  ��    ��� �R�v@/�R{� L�?�Y|8B��c׎�_�R$t����T0 k� � � e1�t B�1	�"q  ��    ��� �R�v@/�R{� L�C�Y|8B��c׎�g�R$D����T0 k� �  � e1�t B�1	�"q  ��    ��� �R�v@/�R{� L�C�Y|8JB�c׎�k�R$D����T0 k� ����e1�t B�1	�"q  ��    ��� �R�u@/�R� L�C�Y|8JB�c׎�o�R D����T0 k� ����e1�t B�1	�"q  ��    ��� �R�u@/�R� L�C�Y|8JB�c׎�s�R D����T0 k� ����e1�t B�1	�"q  ��    ��� �R�u@+�R� L�C�Y|8JB��c׎�w�R D����T0 k� ����e1�t B�1	�"q  ��   ��� �R�u@+�R� L�C�Y|8JB��c׎{�R  ����T0 k� ����e1�t B�1	�"q  ��    ��� �R�u@+�R� L�C�Y|8E2��c׎�R  ����T0 k� ����e1�t B�1	�"q  ��    ��� �R�u@+�R� L�C�Y|8E2��c׎��R ����T0 k� ����e1�t B�1	�"q  ��    ��� �R�u@+�R� L�C�Y|8E2��S׎��R ����T0 k� ����e1�t B�1	�"q  ��    ��� �R�u@+�R� L�C�Y|8E2��S׎��R ����T0 k� ����e1�t B�1	�"q  ��   ��� �R�u@+�R� L�C�Y|8E3�S׎	�R ����T0 k� ����e1�t B�1	�"q  ��    ��� �R�u@+�R� L�C�Y|8EC�S׎	�R d����T0 k� ����e1�t B�1	�"q  ��    ��� �R�u@+�R� L�C�Y|8EC�S׎	� d����T0 k� ����e1�t B�1	�"q  ��    ��� �R�u@+�R� L�C�Y|8EC�S׍	� d����T0 k� ����e1�t B�1	�"q  ��    ��� �R�t@+�R� L�C�Y|8EC�S׍	� d����T0 k� ����e1�t B�1	�"q  ��    ��� �R�t@+�R� L�G�Y|8EC�S׍
�� d����T0 k� � �e1�t B�1	�"q  ��    ��� �R�t@+�R� L�G�Y|8ES�S׌
�� �����T0 k� ��e1�t B�1	�"q  ��    ��� �R�t@+�R� L�G�Y|8ES�S׌
�� �����T0 k� ��e1�t B�1	�"q  ��    ��� �R�t@+�R�� L�G�Y|8ES�S׌
�� �����T0 k� ��e1�t B�1	�"q  ��    ��� �R�t@'�R�� L�G�Y|8ES�S׌
�� �����T0 k� ��e1�t B�1	�"q  ��    ��� �R�t@'�R�� L�G�Y|8ES#�S׌	� �����T0 k� ��e1�t B�1	�"q  ��   ��� �R�t@'�R�� L�G�Y|8ES'�S׌	�����T0 k� ��e1�t B�1	�"q  ��    ��� �R�t@'�R�� L�G�Y|8J�+�S׌	�����T0 k� ��e1�t B�1	�"q  ��    ��� ����C����#
.�Y|8EQ3��v��ó�	R��3��T0 k� �˕�ϕe1�t B�1	�"q  ��"    ��� d���C�����$
.�Y|8EQ+��u��ó�	b��3��T0 k� �Ó�Ǔe1�t B�1	�"q  ��"    ��� b���C�{��ߧ�$
.�Y|8EQ'�ќu��÷�	b��3��T0 k� ����Óe1�t B�1	�"q  ��"    ��� `���C�w��ק�%
�Y|8EQ�єu��÷�	b��3��T0 k� ������e1�t B�1	�"q  ��"    ��� ^���Dk��˨
�&
��Y|8EQ�фu��÷�	b��3��T0 k� ������e1�t B�1	�"q  ��"    ��� [���Dg��ǩ
�'
��Y|8EQ��xt��û�	R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� Y���D_�࿩
�(
��Y|8EQ��pt��û�	R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� V��D[�෩
�(
��Y|8EP���ht���û�	R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� T��DS��
�)
��Y|8E@���`t���û�	R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� R��DO��
�*
��Y|8E@��Xt���û�	R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� P��DG��
�*
��Y|8E@��Lt���ӻ�B��3��T0 k� ������e1�t B�1	�"q  ��"    ��� N��
DC��
�+
��Y|8E@��Ds��ӻ�B��3��T0 k� ������e1�t B�1	�"q  ��"    ��� L��D3��
�,
��Y|8E@׶�4s��ӫ�B��3��T0 k� ������e1�t B�1	�"q  ��"    ��� J��D+����
�-
=��Y|8E@Ϸ�,s��ӣ�B��3��T0 k� ������e1�t B�1	�"q  ��"    ��� H��D'����
�-
=��Y|8E@˸�$s�#�ӟ�B��3��T0 k� ������e1�t B�1	�"q  ��"    ��� F��D���
.|.
=��Y|8E@ø�s�+�ӗ�B��3��T0 k� ������e1�t B�1	�"q  ��"    ��� D��D��{�
.t.
=��Y|8E@���s�3�ӏ�B��3��T0 k� ������e1�t B�1	�"q  ��"    ��� B��D��w�
.l/
=��Y|8E@��	�s�;�Ӌ�B��3��T0 k� ������e1�t B�1	�"q  ��"    ��� @��D� o�
.d/
=��Y|8E@��	�s�?�Ӄ�R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� ?��D� k�
.\0
={�Y|8E0��	��s�G��{�R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� >��D�� g�T1
=s�Y|8E0��	��s�O��w�R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� =!D�� c�L1
=k�Y|8E0��	��s�W��o�R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� <#D� _�D2
=c�Y|8E0��	��s�_��k�R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� ;%D� [�<2
=_�Y|8E0��	��sqg��c�R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� :'C�� W�43
W�Y|8E0��	��rqo��_�R��3��T0 k� ������e1�t B�1	�"q  ��"    ��� 9*C�۔ S�(3
O�Y|8E0{�	��rqs��W�R��3��T0 k� �����e1�t B�1	�"q  ��"    ��� 8,C�ӓ O� 4
G�Y|8E0s�	��rq{��S�R��3��T0 k� �{���e1�t B�1	�"q  ��"    ��� 7.C�ϒ K�4
?�Y|8E0o���rq���K�R��3��T0 k� �w��{�e1�t B�1	�"q  ��"    ��� 70C�ǐ�G�.4
7�Y|8E0g���rq���G�R��3��T0 k� �o��s�e1�t B�1	�"q  ��"    ��� 72C⿏�G�.5
/�Y|8E0c���rq���C�b��3��T0 k� �g��k�e1�t B�1	�"q  ��"    ��� 7�|4Cⷎ�C�. 5
'�Y|8E [��qq���;�b��3��T0 k� �_��c�e1�t B�1	�"q  ��"    ��� 7�x6CⳌ�C�-�5�Y|8E W��qq���7�b��3��T0 k� �_��c�e1�t B�1	�"q  ��"    ��� 7�x8C⫋�?�-�6�Y|8E S��qq���3�b��3��T0 k� �[��_�e1�t B�1	�"q  ��"    ��� 7�t:C⣊�?�
M�6�Y|8E K��pq���+�b��3��T0 k� �W��[�e1�t B�1	�"q  ��"    ��� 7�p<C⛈�?�
M�6�Y|8E G��pa���'� ���3��T0 k� �W��[�e1�t B�1	�"q  ��"    ��� 7�p>C◇�;�
M�6�Y|8E C��oa���#� ���3��T0 k� �W��[�e1�t B�1	�"q  ��"    ��� 7�hBC��;�
M�6��Y|8E ;���na���� ���3��T0 k� �S��W�e1�t B�1	�"q  ��"    ��� 7�dDC���;�
M�7��Y|8E 7���na���� ���3��T0 k� �S��W�e1�t B�1	�"q  ��" 
   ��� 7�`EC�{��;�
M�7��Y|8E 3�	Ѐna˿�� ���3��T0 k� �S��W�e1�t B�1	�"q  ��" 
   ��� 7�\GC�s� p;�
M�7��Y|8E /�	�|maӿ�� ���3��T0 k� �W��[�e1�t B�1	�"q  ��" 
   ��� 7�XIC�k� p;�
]�7,��Y|8E+�	�xma׾�� ���3��T0 k� �W��[�e1�t B�1	�"q  ��" 
   ��� 8�TKC�c� p;�
]�6,��Y|8E'�	�tma۽�����3��T0 k� �W��[�e1�t B�1	�"q  ��" 
   ��� 9�PLC�_� p;�
]�6,��Y|8E#�	�lma߼�����3��T0 k� �W��[�e1�t B�1	�"q  ��" 
   ��� :�HNC�W� p;�
]�6,��Y|8E#�	�hla������3��T0 k� �[��_�e1�t B�1	�"q  ��" 
   ��� ;�DPC�O� p?�
]�6,��Y|8E�	�dlQ������3��T0 k� �[��_�e1�t B�1	�"q  ��" 
   ��� <�@QC�G� p?�
]|6��Y|8E�	�`lQ������3��T0 k� �[��_�e1�t B�1	�"q  ��" 
   ��� =�8SD?� p?�
]t6��Y|8E�	�\lQ������3��T0 k� �[��_�e1�t B�1	�"q  ��" 
   ��� >�4UD3� pC�
]l5��Y|8E�	�XlQ������3��T0 k� �_��c�e1�t B�1	�"q  ��" 
   ��� ?�0VD+� �C�
]d5��Y|8B���TlQ������3��T0 k� �_��c�e1�t B�1	�"q  ��" 
   ��� @�(XD#� �C�
]\5��Y|8B���Pl�������3��T0 k� �c��g�e1�t B�1	�"q  ��" 
   ��� A�[D� �G�
]L4��Y|8B���Lk�������3��T0 k� �g��k�e1�t B�1	�"q  ��" 
   ��� B�\D� �K�
MD4��Y|8B���Hk�������3��T0 k� �g��k�e1�t B�1	�"q  ��" 
   ��� C�^D� �K�
M<4���Y|8B���Dj�����R��3��T0 k� �k��o�e1�t B�1	�"q  ��" 
   ��� D�_D�� �O�
M43���Y|8B�� @j�����R��3��T0 k� �k��o�e1�t B�1	�"q  ��" 
   ��� E�aD� �S�
M,3��Y|8B�� <i�����R��3��T0 k� �o��s�e1�t B�1	�"q  ��" 
   ��� F                                                                                                                                                                            � � �  �  �  c A�  �J����  �      � \���� ]�%'%& � �� tgH    >      � ���     tw� �ٕ    ��A                  9 �          �     ���   0		 
 
         ���        �	ɦ    ��*�	ט    ���.              � �          Ep     ���   (	 
          ���t           �=�    ���� �/�     � �              	    �         �      ���   8�          |u           �ug     T� �ug    S     	              ��                ���   (
          ��%           . �u�    ��� �gT     o �                ����          ��      ���   P
B           ݒ ��	     B���     ݒ���                           ���e              A  ���    81
           ���? � U     V �W    ��.� �Fn    ��               L �� �          �0
�   
  ��P  8	
           ��R%  � �	   j �hW    ��R% �hW                    @�� �          �   �  ��@   0	          ����  � �     ~ �    ���J �KP    ��H            	�� �          �`�    ��@  8
	           �R  � � 
	   � ��     ~6 �<    \�g              ' �� �         	 �     ��h  @

(         ���Z        ��2    ���t�    ��               L�� �         
 ��   
  ��@  H

 

         ��is ��       � �3�    ��is �3�                              ���I              o  ��@    8		'                ��      �                                                                           �                               ��        ���          ��                                                                 �                          V�  ��        � �u�     ?� ��|    \�g                   x                j  �    	   �                              ��        � �          �           "                                                 �                          �	 � � �� � � � � ��� � �       	  
        
  �   � ���L       � �t� �  u� �� @p� �d q  � �t� �  u� 6�  p� �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0� ���� ����� ����� � � 0i@ �d  i� פ i� � �r@ � s@ �d 0j� �� 0k  �$ k� �D  k� ��  k� $ @m@ � m� �  m�  n  � �t� �  u� � �c@ � d@���� � L�  a� H� �o� I�  p� J q  J$ q@ �� @m@ �d `m� �$ 0n� �� n� 
�< V� 
�� V� 
�| W  
�\ W� 
� W� 
�| W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� � �����  ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"    B�j
��  B �
� �  �  
�      ��     � �      ��    ��     �	           ��     � �          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �((      �� �T ���        �?T ��        �        ��        �        ��        �     ��    ��� �	        ��                         T�) , �� ��                                    �                ����            	  �	���%��  �� � ���2           20 Bob Sweeney ne      4:32                                                                        4  4     �C
�2Y �<X �;Fc�3> c�;:C. �O C6 �6CO-	C �M 
C �kV �k^ � � ~ � �	c � �c� � � c� � �cj � �cn � �cp � �cs � � cw � � cx � � c� �c� �c� � �c� � �J� �	�$ �	�; ��" ��Mh "�3h !"�EX"�/X#
�> �$"�
 � %"� �&"� �'*�h("�3h )"�EX*�/X+
�> �,!� | � -"G � �."( � � /"O � � 0"H � �1"6 � �2" � � 3"R � � 4"O � r5"$ � �6" � �7""D r8"T r9*$t � :"J � � ;"K � � <"B �="  | >"J �2 !� |                                                                                                                                                                                                                         �� P             @ 
      6 �     W P E a  ��        	            �������������������������������������� ���������	�
��������                                                                                          ��    �I�   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, 5� $ �� �� �@ɂ�A���                                                                                                                                                                                                                                                                                                                                        0@�                                                                                                                                                                                                                                          u    '    ��  L�J      	�  	                           �������������������������������������������������������                                                                      
                                                                  ]    " (            �          �   r             	 	 ���������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ����            x             
        *     �  9<�J      !                             ������������������������������������������������������                                                                                                                                        x  ��                  �     �   �                  ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� ������������������           �                                                                                                                                                                                                                                                
                                         	                   �             


           �   }�         ������������  '�  '|    ������������������������  N�����������������������������������������������������                                           +           N�  'v                     �ww�ww333wwwwwwww�ww�ww�ww�ww333wwww N @ 0 
                                � , � �t�                                                                                                                                                                                                                                                                                   )n)n�  
                        k      k                  k                                                                                                                                                                                                                                                                                                                                                                                                                            � � �  � ��  � (��  � (��  � @��  � ��  �����������P����������������������M����p�����p�                 w � :��	          �   & AG� �  �                 �                                                                                                                                                                                                                                                                                                                                      p I G   f                       !��                                                                                                                                                                                                                            Y    �� �� Ѱ�      �� X      ���������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ���� ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� ������������������             $�l�������l����������������������l��������������f���f���f��ff���f������ffffflffffffffffffffffffff����ff��lfflffffffffffffffffffffl��l��̼���l����l��lf���ll��������l�����ll������l�����������������l���������������l��������������fff�lff�ll��l���li��f���l���f��ffffffffffff��������������������fffffff�ffl��̻�����������������f�l���l�llll�l�̦ll̜f�̊�l̊���l����������������������������������������������������������������f���f���f���f���f���f��ɜ�����������������������̺��ƹ��li��fiy��������������˩�ff��fl��fk��fj���f̈�f̈�f̈�f̈�fl�{ʜ�����������l����������������̼��������������������������������������̼̼��������j���ˊ��̗��̸���ʈ���Ɉ��i���������������������������y��fj���k���̨��̹��l���̹��lɹ��ʘ�����ɬ��ȼ�������l���̘��̈���������̼����̼������̼�����̼��������������̼���������̼���̼̼���k�̼̈��̈��ˈ��˘̼����˘��̘�Ɉ����������������ˈ�����������k��ɫ��ɫ����ff��ɶ��ɻ�ll���������̉��ˈ��̈��̙��ˈ�̼���l�����������������̼����˼�̶���̻�������������˨̩��������������������ʈ����������|����i����Ʒi��i��������������������������j���f��������̹�̼���̘�fʘ��ɉ����̊�̼��ȸ�{�Ɉ��h�����l���j���h��fȹ����̈xx�������������f���l��l�������    (      8   �                        4     �   �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$ ^h  ��     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@       �      �    ������ ��  �� t� � �� t� � �$  �B  �� � B      �  ��  t���� e�����   g���        f ^�         �� ��     t      ���F���2�������J������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "" "  """ "! ""! " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  ""   "! " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """ "! ""! " ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         � 
��	�˽���w��{k��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            �  �  �  ��  �           K�  ��� ڬ� ۻ� +�" """ """ �"" ��"/����� ��   ��  ��  ��                        �          �   � � �  ��� ��  �                       �   �                      �������  ���    ��   �   ��� ������ �   �      �       �                        �   ��  ���  � �    �                                ����                  �   �� �       �  �  ��  �   �   �   �                                     �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �   �   �   ˰  ˙  ɪ  ��� ټ� �̰ �̰ ��� ��  ��                              ��                  �                        ���� ��� ����                            ��  ��  ���  �  �  �   �   ��  �                            �   ���                            �   �                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��               �   �   �  �  �  �  �   �   �                                       �  ���   �                          �   �   ��� ������ �   �      �       �                        �   ��  ���  � �    �                                                                                                                                        �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �            �  �� �  �  �   �     "  "  "                       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����            ����  �  �  �  �  ��  �                      � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        ɪ  ��� ټ� �̰ �̰ ��� ��  ��              �   ������  ��                   �                        ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                        �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �    � � �     �   �                   �  �� Ș ��  ��  �      �  �   �  �  ��  �  ��  �                                                                                                                    �  �  ��  �                                                                                        �  ɪ� ɪ� ̚� �ȍ ͷ  "�  "� .( 3># �4�
�T��T�"�UN"�UN(�Dɜ� ʨ����, � /�������� � ��                                ��  ��  ��  g}  �א vz� gz� ̊� �ɩ 8̜ D<� T� @��  �� ɀ ��  ��  "   .          �  ��� �������  ��                           "  "  "  "                  �   �   ��  �   �   �   �               �   �    �   �       �   �   �                .                      ��� ���� ��             �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                      �  ��� ݻ� g�� bm� ggz�'w���������������˛������ˊۼ�����˻������H�DH�@U�DPT�E X�T H�P H�@ Ȥ� ̻� ˘ "�� � ���/�"" �""/���               �   �                                                     �  �                      � �                       ���           �                      �  �  �          ����  �   �             ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                       �   ���                            �   �                                                                                                                1    1   "    �   �   �� �����  �    �   �   ,   "   "                   ���ۼ����� 9��C��UTDD�D33��0��  "��
/� � �, �"  �"   �   ˻ڛ��Ȱ��  ��  ��  TJ  EJ  DT  4E  �P  ��  �   /   ��  ��� �                                     � 	�� �� �˙	���
������                Ͱ  ˻  ˻  ۻ  ݻ  ��  ��� ��� ��˰��˰̼˚̽��                               �   �                .          � ��                    ���� �                                                                                                                                                                                          �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw         � ��                    ���� �                                              ����     �   �  �  �  ��  �   �                           ��   ��                  �  �  �� � ���                                                �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �                �                             ���                         �  ��                    �����                      �  �  �   �   ��  �                            �   ���                            �   �                                                                                                                     �� �����ݼڜ��ک��ک��z�	��� 
�� 
�� 	�� ̘ ɪ  ��  �  �� �� ������������ ���  � � � �� �� ������ ��                      �   ��  ��  �̰ ��� ��˰�̻��̻���������ˉ�U��EP�ET �I� ٕ  �D� �L� ��� ��" ����/�"�"�""�����                         ��  ��� ��  �                                        �� ��                  �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""������������������""""������������������������""""������������������������""""������ADAIA�A""""�������I�A�A�A""""�����DD�I""""�������DAADAI""""������IDA��""""��������DD��I�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD������������������������3333DDDD�A�AM�M�DM��M334CDDDD�A�AM�M�DDM����3333DDDDDM����DD�����3333DDDDMAM��D�DDM�����3333DDDDDD����M��DM�����3333DDDD������������DD������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��           	 
          
        ((((((( 
	(((( ����������������             ! " # $ % & '   ( $ % ) ! " # * ('(&(%($(#("(! (((���������������� + , -   . / 0 1  	 2         3       4 (((((((2	10/(.(-(,(+���������������� 5 6   7   8 9 1 :   $ % ) ! " #   ; ) ! " # $ % ) (#("(!()(%($ :198(((7(6(5����������������    <     = 8 0 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>108(=((( (<���������������� L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L����������������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7����������������  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
�2Y �<X �;Ec�3= c�;:C. �O C6 �6CO-	C �M 
C �kV �k^ � � ~ � �	c � �c� � � c� � �cj � �cn � �cp � �cs � � cw � � cx � � c� �c� �c� � �c� � �J� �	�$ �	�; ��" ��Mh "�3h !"�EX"�/X#
�> �$"�
 � %"� �&"� �'*�h("�3h )"�EX*�/X+
�> �,!� | � -"G � �."( � � /"O � � 0"H � �1"6 � �2" � � 3"R � � 4"O � r5"$ � �6" � �7""D r8"T r9*$t � :"J � � ;"K � � <"B �="  | >"J �2 !� |3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������ �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������$��7�O�Q�K��;�O�I�I�O� � � � � � � � � � �:�>�/�����������������������������������������$��4�U�K��<�G�Q�O�I� � � � � � � � � � � �:�>�/�������������������������������������������,�U�H��<�]�K�K�T�K�_� � � � � � � � � �,�>�0�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������:�>�/� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������,�>�0� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $������������������������     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %������������������������ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                