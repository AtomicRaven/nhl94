GST@�                                                           `m�                                                      r                          ���2���� 
 J�����������H���z���        �h      #    z���                                d8<n    �  ?     h����  �
fD�
�L���"����D"��   " `  J  jF��    "�j "����
��
��     �j�� 
   ��
  7�                                                                              ����������������������������������      ��    =b 0Qb 4 114  4c  c  c        	 
      	   
       ��G �� � ( �(                 Enn )1         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                �          �   @  &   �   �                                                                                 '      E)n1n  �    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������     ��@c�A���l@A�,-Y|,��}"�B�`�p��p3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�,.Y|,��}"�D�`	�o��p3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�,.Y|,��}"�F�_	�o��o3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�,/Y|,��}"�H�_	�o��o3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�,/Y|,��~"�J�^	�os�o3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�00Y|,��~�L�^	�ns�n3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�00Y|,��~�N�^Sns�n3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�00Y|,��~�P�^Sns�m3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�01Y|,��~�R�]Sms�m3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�01Y|,��~�R�]Smc�l3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�02Y|,��~�R�]Smc�k3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�02Y|,���S�]Smc�k3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�42Y|,���T�]Smc�j3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�43Y|,���U� ]Smc�i3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�43Y|,���V� ]Slc�i3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�43Y|,���W�$]S lS�h3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�44Y|,����X�$]S lS�g3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�44a�,����Y�(]S lS�g3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�44a�,����Z�(]S lS�f3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�45a�,�Ԁ��[�(]c lS�e3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�85a�,����\�,]c l��e3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�85a�,����\�,]c l��d3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�86a�,����\�,]c l��c3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�86a�,����\�,]c m��c3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�86a�,��~��\�,]cm��b3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A��l@A�87a�,��~��\�,]cm��a3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�|�l@A�87a�,��~��\�0]cn��a3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�|�l@A�87a�,��~��\�0]cn��`3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�|�l@A�88Y|,��}��\�0]cn��`3��T0 k� �����&5AC"3Q �2	4#Q  ��K   �  � ��@c�A�|�l@A�<8Y|,��}��]�0]cn��_3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�|�l@A�<8Y|,��}r�]�0]co��^3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�|�l@A�<8Y|,��}r�]�0]co��^3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�|�l@A�<9Y|,��}r�]�0]co��]3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�x�l@A�<9Y|,��}r�]�0]co��]3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�x�l@A�<9Y|,��}r�]�0]co��\3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�x�l@A�<:Y|,��}r�]�0]cp��\3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�x�l@A�<:Y|,��}r�]�0]cp��[3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�x�l@A�<:Y|,��}r�]�0]cp�[3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�x�l@A�@:Y|,��}r�]�0]cp�Z3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�x�l@A�@;a�,��}r�]�0]cp�Z3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�t�l@A�@;a�,r�}r�]�0]cp�Y3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�t�l@A�@;a�,r�}��]�0]cp�Y3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A�t�l@A�@;a�,r�}��]�0]cp�X3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  ��TE�E����fE�8Y|,����������@63�	T0 k� ��Z��Z&5AC"3Q �2	4#Q  ��    � 2 f�TE�+�E���gE�@Y|,��������#��P63�	T0 k� ��Z��Z&5AC"3Q �2	4#Q  ��    � 2 e�TE�3�E��� gE�HY|,��������+��\63�	T0 k� ��Z��Z&5AC"3Q �2	4#Q  ��    � 2 d�TE�?�E���$hE�PY|,�ǂ�����3��h63�	T0 k� ��Z��Z&5AC"3Q �2	4#Q  �� 	   � 2 cTE�G�E�߾,iB�Xa�,�ς.�����;��p63�	T0 k� �Z��Z&5AC"3Q �2	4#Q  �� 	   � 2 b�TE�O�E�߽4jB�`a�,�ׂ.��ј�C��|63�	T0 k� �Z��Z&5AC"3Q �2	4#Q  �� 	   � 2 a�TE�[�E�߻<jB�ha�,�߃.��ќ�K���63�	T0 k� �Z��Z&5AC"3Q �2	4#Q  �� 	   � 2 `� TE�c�E�߹DkB�pa�,��.��ќ�O���63�	T0 k� �Z��Z&5AC"3Q �2	4#Q  �� 	   � 2 _�(TE�o�E�߷LlB�xa�,��.��ќ�W���63�	T0 k� �Z��Z&5AC"3Q �2	4#Q  �� 	   � 2 ^�8TE���E�ߴ\mB��a�,��/�Ѡ�g���63�	T0 k� �Z��Z&5AC"3Q �2	4#Q  �� 	   � 2 ]�@TE���E�߲�dmB��a�,��/�� �o���63�	T0 k� �Z��Z&5AC"3Q �2	4#Q  �� 	   � 3 _�LTE���E�߰�lnB��a�,��/��"�s���73�	T0 k� �Y��Y&5AC"3Q �2	4#Q  ��3 	   � 4 `�TTEp��C�߯�tnB��a�,��/'��#�{���73�	T0 k� �X��X&5AC"3Q �2	4#Q  ��3 	   � 5 a�\TEp��C�߭�|oB��a�,�#�//��%���	�73�	T0 k� �Y��Y&5AC"3Q �2	4#Q  ��3 	   � 6 b�dUEp��C�۫��oB��Y|,�+��7��&���	�73�	T0 k� �Y��Y&5AC"3Q �2	4#Q  ��3 	   � 7 c�lUEp��C�۪	��oC�Y|,�3��?��'���	�73�	T0 k� �\��\&5AC"3Q �2	4#Q  ��3 	   � 8 d�tUEp��C�ר	�pC�Y|,�?��G��)���	�73�	T0 k� �Y��Y&5AC"3Q �2	4#Q  �3 	   � 8 ]�|VEp��C�צ	�pC�Y|,�G��O��*���	73�	T0 k� �V��V&5AC"3Q �2	4#Q  ��? 	   � 8 W��WEp��C�ӣ	�qC�Y|,�W��_��-���	73�	T0 k� �xQ�|Q&5AC"3Q �2	4#Q ��? 	   � 8 Q��WEp��C�Ϣ�qC�Y|,�_��k��.���	"73�	T0 k� �lO�pO&5AC"3Q �2	4#Q ��? 	   � 8 K��XEp��C�ˠ�qC�Y|,�g��s��/���	"$73�	T0 k� �`L�dL&5AC"3Q �2	4#Q ��? 	   � 8 E��XEp��C�˟�rC�Y|,�o��{��0�ǰ	",73�	T0 k� �PI�TI&5AC"3Q �2	4#Q ��? 	   � 8 ?��YEp��C�Ǟ�rC�Y|,�w�����1�ϯ	"473�	T0 k� �DG�HG&5AC"3Q �2	4#Q ��? 	   � 8 9��ZEq�C�Ü��rC�Y|,������3�ׯ	"<73�	T0 k� �8D�<D&5AC"3Q �2	4#Q ��? 	   � 8 4��[Ea�C���rCY|,�������4�ۮ	@73�T0 k� �,B�0B&5AC"3Q �2	4#Q ��? 	   � 8 /��\Ea�C���sCY|,�������5��	H73�T0 k� � ?�$?&5AC"3Q �2	4#Q ��? 	   � 8 *��\Ea�C���sCY|,�������6��	P73�T0 k� �<�<&5AC"3Q �2	4#Q ��? 
   � 8 %��]Ea#�C���sCY|,�������7��	T73�T0 k� �:�:&5AC"3Q �2	4#Q ��? 
   � 8  ��^Ea+�C���tC$Y|,�������|8���	\73�T0 k� ��7��7&5AC"3Q �2	4#Q ��? 
   � 8 ��_D1/�C���tC,Y|,�������x9��	"`73�T0 k� ��5��5&5AC"3Q �2	4#Q ��? 
   � 8 ��`D17�C���tC4Y|,�������t;��	"d73�T0 k� ��2��2&5AC"3Q �2	4#Q ��? 
   � 8 ��aD1;�D����tC<Y|,�������p<��	"l73�T0 k� ��0��0&5AC"3Q �2	4#Q ��? 
   � 8 ��bD1C�D����uCDY|,�Ð����l=��	"p73�T0 k� ��-��-&5AC"3Q �2	4#Q ��? 
   � 8 	��cD1G�D����uCLY|,�ˑ����d>�#�	"x73�T0 k� ��*��*&5AC"3Q �2	4#Q ��? 
   � 8 ��eEaK�D��� uCTY|,�ϒ����`?�+��|73�T0 k� ��(��(&5AC"3Q �2	4#Q ��? 
   � 8 � fEaO�D���uC\Y|,�ד����\@�/���73�T0 k� ��%��%&5AC"3Q �2	4#Q ��? 
   � 8���gEaS�D���vC.dY|,�ߔ����XA�7���73�T0 k� ��#��#&5AC"3Q �2	4#Q  ��? 
   � 8���hEaW�D��vC.hY|,������PB�?���73�T0 k� �� �� &5AC"3Q �2	4#Q  ��? 
   � 8���iEa[�E�w��vC.pY|,�����LC�G���73�T0 k� �x�|&5AC"3Q �2	4#Q  ��? 
   � 8���jE�_�E�o��vC.xY|,�����DD�O���73�T0 k� �l�p&5AC"3Q �2	4#Q  ��? 
   � 8���kE�c�E�k��vC.�Y|,�����@D�W���73�T0 k� �`�d&5AC"3Q �2	4#Q  /�? 
   � 8���mE�g�E�c�� wC.�Y|,������8E�_���73�T0 k� �T�X&5AC"3Q �2	4#Q  ��? 
   � 8���oE�o�E�W��,wC.�Y|,���#��,G�o���73�T0 k� �<�@&5AC"3Q �2	4#Q  ��? 
   � 8��� pE�o�E�O��0wC.�Y|,���+��(G�w�"�73�T0 k� �,�0&5AC"3Q �2	4#Q  ��? 
   � 7��� qE�s�E�G��4xC.�Y|,���/�� H��"�73�T0 k� � �$&5AC"3Q �2	4#Q  ��? 
   � 6���$rE�w�E�?��8xC.�Y|,���3��I���"�73�T0 k� �	�	&5AC"3Q �2	4#Q  ��? 
   � 5���$sE�w�E�7��<xE��Y|,���;��I���"�63�T0 k� ��&5AC"3Q �2	4#Q  ��?    � 5���$tE�{�E�/��@xE��Y|,���?��I���"�63�T0 k� ����&5AC"3Q �2	4#Q  ��D    � 5���(uE�{�C�'��DxE��Y|,���C��J���"�63�T0 k� ����&5AC"3Q �2	4#Q  ��D    � 5���(wE��C���PxE��Y|,���K���K���"�53�T0 k� ����&5AC"3Q �2	4#Q  ��D    � 5���(xE��C���TxE��Y|,���O���K���2�53�T0 k� ����&5AC"3Q �2	4#Q  ��D    � 4���(yEa��C���XxE��Y|,���S���K ��2�43�T0 k� ����&5AC"3Q �2	4#Q  ��D    � 4���(zEa��C����\xE��Y|,�#��W���K ä2�43�T0 k� ����&5AC"3Q �2	4#Q  ��D    � 4���({Ea��C����`xE��Y|,�#��[���K ˣ2�33�T0 k� ����&5AC"3Q �2	4#Q  ��D    � 3���(|Ea��C���lxE� 
Y|,�'��_���K ۣ2�23�T0 k� �'��+�&5AC"3Q �2	4#Q  ��D    � 2���$}Ea�C�߃�px@
Y|,�'��c���K0ߣ2�23�T0 k� �/��3�&5AC"3Q �2	4#Q  ��D    � 2���$~Ea�C�׃qxw@	Y|,�'��c���K0�2�13�T0 k� �7��;�&5AC"3Q �2	4#Q  ��D    � 1���$Ea�C�˃q|w@	Y|,�'��g��J0�2�03�T0 k� �?��C�&5AC"3Q �2	4#Q  ��D    � 1��� �Ea�I�Ãq�w@ Y|,�'��g��J0��B�/3�T0 k� �G��K�&5AC"3Q �2	4#Q  ��D    � 0��� �D1�I���q�v@(Y|,�'��g��J0��C .3�T0 k� �O��S�&5AC"3Q �2	4#Q  ��D    � 0���D1�I���q�u@8Y|,�#��k��IA�C-3�T0 k� �_��c�&5AC"3Q �2	4#Q  ��D    � / �D1�I���q�u@@Y|,�#��k� �HA�C,3�T0 k� �g��k�&5AC"3Q �2	4#Q  ��D    � . �D1�I���q�t@HY|,�#��k� �HA��+3�T0 k� �o��s�&5AC"3Q �2	4#Q  ��D    � - ~D1�I���q�t@LY|,�#��k� �GA��+3�T0 k� �w��{�&5AC"3Q �2	4#Q  ��D    � - ~D1�I���q�s@TY|,���o� �FA#��*3�T0 k� �����&5AC"3Q �2	4#Q  ��D    � , 
~D1�I���q�r@\Y|,���o� �FA'��)3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � , ~D1|I���a�q@�dY|,���o� �EA/��)3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � + ~D1|I��a�q@�lY|,���o�ЀDA3��(3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � *  }D1xI�w�a�p@�tY|,���o��|DA;�� (3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � * �}D1tI�o�a�n@�� Y|,���o��xBAG��$'3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � ) �}Eat!I�g�a�m@�� Y|,��o��tAAK��$&3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � ( �|Eap$I�c�a�l@���Y|,��o��p@QO��$&3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � ' �|Eap&I�_�a�k@���Y|,��o��l?QW��$%3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � & �|Eal(I�[�a�j@���Y|,��o��l>Q[��$%3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � % �|Eah*I�W�a�i@���Y|, ���o��h=Q_��($3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � % �|Eah,I�S�a�h@���Y|, ���o��h<Qg��(#3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � $  �{Ead.I�O�Q�g@���Y|, ���s��d;Qk��(#3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � # "�{Ea`0I�K�Q�f@���Y|, ���s��d:Qo��("3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � " $�{Ea\2I�G�Q�e@���Y|, ���s��d9Qs��("3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � " &�{EaX5I�C�Q�d@���Y|, ���s��`8Q{��(!3�T0 k� ������&5AC"3Q �2	4#Q  ��D    � ! (�{EQT7I�C�Q�c@���Y|, �� s��`7Q��$ 3�T0 k� ������&5AC"3Q �2	4#Q  ��D    �   *�{EQP9I�?�Q�b@���Y|,�� s��`5Q���$3�T0 k� �����&5AC"3Q �2	4#Q  ��D    �  ,�zEQH=I�;�Q�`@���Y|,�� s��\3a���$3�T0 k� ����&5AC"3Q �2	4#Q  ��D    �  .�zEQD?I�7�Q�`@���Y|,�� w��\2a���$3�T0 k� ����&5AC"3Q �2	4#Q  ��D    �  0�zEQ@AI�3�Q�_@���Y|,�� w��\0a���$3�T0 k� ����&5AC"3Q �2	4#Q  ��D    �  2�zEQ<CI�3�Q�^@���Y|,��� w��\/a��$3�T0 k� �#��'�&5AC"3Q �2	4#Q  ��D    �  4�zEQ8EI�/�Q�]@��Y|,��� {��\-a��$3�T0 k� �#��'�&5AC"3Q �2	4#Q  ��D    �  6�yEQ0GI�/�Q�\@��Y|,л��{��`,a��$3�T0 k� �'��+�&5AC"3Q �2	4#Q  ��D    �  8�yEQ,II�/�Q�[@��Y|,з����`+a��$3�T0 k� �'��+�&5AC"3Q �2	4#Q  ��D    �  :�xyEQ(JI�+�Q�Z@��Y|,Я����`)a��(3�T0 k� �+��/�&5AC"3Q �2	4#Q  ��D    �  <�lyEQNI�+�Q�Y@�+�Y|,У�����`&a���(3�T0 k� �;��?�&5AC"3Q �2	4#Q  ��D    �  >�dyEAPI�+�Q�X@�/�Y|,Л�����d%q���(3�T0 k� �?��C�&5AC"3Q �2	4#Q  ��D    �  @�\xEAQI�'�Q�W@�7�Y|,�������d#q���(3�T0 k� �G��K�&5AC"3Q �2	4#Q  ��D    �  B�TxEASI�'�Q�V@�?�Y|,�������h"q���,3�T0 k� �O��S�&5AC"3Q �2	4#Q  ��D    �  D�LxEATI�'�Q�V@�G�Y|,�������h qô�,3�T0 k� �W��[�&5AC"3Q �2	4#Q  ��D    �  F�8xE@�WI�'�Q�TE S�Y|,�{�����lq˷03�T0 k� �c��g�&5AC"3Q �2	4#Q  ��D    �  H�0xE@�YI�'�Q�SE [�Y|,�s�����pqϹ03�T0 k� �k��o�&5AC"3Q �2	4#Q  ��D    �  J�(xE@�ZI�'�Q�SE _�Y|,�k���� pqӺ4
3� T0 k� �s��w�&5AC"3Q �2	4#Q  ��D    �  L� wE@�[I�'�Q�RE g�Y|,�c���� tq׼4	3� T0 k� �w��{�&5AC"3Q �2	4#Q  ��D    �  N�wE@�]I�'�Q�QEw�Y|,�S���� xqۿ83� T0 k� ������&5AC"3Q �2	4#Q  ��D    �  P�wE@�^A�'�Q�PE{�Y|,�O���� |A��<3� T0 k� ������&5AC"3Q �2	4#Q  ��D    �  R� wE@�_A�'�Q�OE��Y|,�G���� �A��@3� T0 k� �����&5AC"3Q �2	4#Q  ��D    �  T��wE0�`A�'�Q�OE��Y|,�?���� �A��@3� T0 k� �����&5AC"3Q �2	4#Q  ��D    � 
 V�wE0�aA�'�Q�NE��Y|,�7���� �A��D 3� T0 k� �����&5AC"3Q �2	4#Q  ��D    � 	 X�vE0�bA�'�Q�ME��Y|,�'���� �	1���K�3��T0 k� �����&5AC"3Q �2	4#Q  ��D    �  Z�vE0�cB@'�Q�LE��Y|,�����	�1���O�"s��T0 k� �����&5AC"3Q �2	4#Q  ��D    �  \�vE0�dB@'�Q�KE��Y|,��@��	�1���S�"s��T0 k� �����&5AC"3Q �2	4#Q  ��D    �  ^�vE0�dB@'�Q�KE��Y|,��@��	�1���W�"s��T0 k� ������&5AC"3Q �2	4#Q  ��D    �  `�vE0�eB@'�Q�JE��Y|,��@��	�1���_�"s��T0 k� ������&5AC"3Q �2	4#Q  ��D    �  c�vE0�eB@'�Q�IE���Y|,���@��	��"��c�"s��T0 k� ������&5AC"3Q �2	4#Q  ��D    �  f�vE0�e@'�Q�HE���Y|,���@��
 ��"��g�"s��T0 k� ������&5AC"3Q �2	4#Q  ��D    �  h�vE0xe@'�Q�HE���Y|,���@��
 ��"��k�"s��T0 k� ������&5AC"3Q �2	4#Q  ��D    �  k�uE0te@'�Q�GE���Y|,���@��
 ��"��o�"s��T0 k� ������&5AC"3Q �2	4#Q  ��D    �   m|uE he@'�Q�FBP��Y|,���@��
 ��"��{�"s��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� ptuE deB�+�Q�FBP��Y|,���P��	��"���3��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� sluE `eB�+�Q�EBQ�Y|,��P��	��"����3��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� uduE XeB�/�Q�DBQ�Y|,��P��	��"����3��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� wTuB�PeB�3�R CBQ�Y|,��P��	��"'����3��T0 k� �+��/�&5AC"3Q �2	4#Q  ��D    ��� z	�LuB�LdB�3�R CBQ�Y|,�� ��
 ��"'����3��T0 k� �3��7�&5AC"3Q �2	4#Q  ��D    ��� }	�DuB�HdB�7�R BBQ'�Y|,��!�
 ��"+����3��T0 k� �;��?�&5AC"3Q �2	4#Q  ��D    ��� 	�<uB�DdB�;�R BBQ/�Y|,��!�
 ��"/����3��T0 k� �C��G�&5AC"3Q �2	4#Q  ��D    ��� �	�4uB�@cB�;�R ABQ7�Y|,��!�
 ��"/����3��T0 k� �K��O�&5AC"3Q �2	4#Q  ��D    ��� �	�,uB�@cB�?�R ABQ?�Y|,��!�
 ��"3����3��T0 k� �S��W�&5AC"3Q �2	4#Q  ��D    ��� �	� uB�8bB�G�R@BQO�Y|,��!�	��"7����3��T0 k� �c��g�&5AC"3Q �2	4#Q  ��D    ��� �	�uC 8aB�K�R?BaW�Y|,��!�	��";����"���T0 k� �k��o�&5AC"3Q �2	4#Q  ��D    ��� �	�uC 4aB�O�R?Ba_�Y|,����	��2;����"���T0 k� �s��w�&5AC"3Q �2	4#Q  ��D    ��� �	�uC 4`B�S�R?Bag�Y|,���#�	��2?����"���T0 k� �{���&5AC"3Q �2	4#Q  ��D    ��� �	�uC 0`B�W�R>Bao�Y|,���+�	��2?����"���T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� �	� uC 0_B�[�R>Baw�Y|,���/�
 ��2C����"���T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ���uC ,]B�g��=E���Y|,���7�
 ��2G����"���T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ���uC ,]E�k��<E���Y|,���?�
 ��2G����"���T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ���uC (\E�o��<E���Y|,���@ 
 ��2K����"���T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ���uE ([E�w��<E���Y|,���H	��2K����"���T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ���uE (ZE�{��;E���Y|,���L	��BK����"���T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ���uE (YE���;E���Y|,���T	��BO����3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ���uE (WE����:E���Y|,���`	��BS���3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ���uE (VE���� :E���Y|,����d@��BW���3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� �иuE (UE���� 9E���Y|,����l@��BW���3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ��uE(TE�����9E���Y|,����t@��
�[���3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ��uE,SDУ���8E���Y|,����x@��
�_���3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ���tE,QDЯ���8E���Y|,��������
�c��#�3��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� ���tE,PDз���7E���Y|,���ь���
�g��#�3��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� ���tE�0ODп���7E���Y|,���є���
�k��'�3��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� ���tE�0NE�Ǌ��7E��Y|,���Ѡ���
�k��+�3��T0 k� ���#�&5AC"3Q �2	4#Q  ��D    ��� ��|sE�4ME�ˊ��6@r�Y|,���Ѭ���
�o��+�3��T0 k� �'��+�&5AC"3Q �2	4#Q  ��D    ��� ��tsE�4LE�Ӌ��6@r�Y|,���Ѹ���
�s��/�3��T0 k� �/��3�&5AC"3Q �2	4#Q  ��D    ��� ��drE�<JE����5@r#�Y|,��������
�{��/�3��T0 k� �?��C�&5AC"3Q �2	4#Q  ��D    ��� ��\rE�<HE����5@r+�Y|,ϛ������
���3�3��T0 k� �G��K�&5AC"3Q �2	4#Q  ��D    ��� ��TqE�@GE����5E3�Y|,ϛ������
����3�3��T0 k� �K��O�&5AC"3Q �2	4#Q  ��D    ��� ��LqE�DFE����4E;�Y|,ϟ��� ���
����3�3��T0 k� �O��S�&5AC"3Q �2	4#Q  ��D    ��� ��DpE�DEB���4EC�Y|,ϣ��� ���
����3�3��T0 k� �W��[�&5AC"3Q �2	4#Q  ��D    ��� ��<oB�HCB���4EK�Y|,ϧ������
����3�3��T0 k� �_��c�&5AC"3Q �2	4#Q  ��D    ��� ��4oB�LBB���4ES�Y|,ϫ������
����3�3��T0 k� �g��k�&5AC"3Q �2	4#Q  ��D    ��� ��$mB�T?B�#��4Ec�Y|,ϳ��#����
����3�3��T0 k� �w��{�&5AC"3Q �2	4#Q  ��D    ��� �� lB�X>B�+��3Ek�Y|,Ϸ��+����
���43�3��T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ��kE\=B�3��3Es�Y|,ϻ��3����
���43�3��T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ��jE`<B�?��3E{�Y|,Ͽ��?����
���43�3��T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ��iEd:B�G��3E���Y|,�á�G����
���43�3��T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� �� hEh9B�O��3E���Y|,�ˠ�O���R��43�c��T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ���gEl8B�W��3E���Y|,�Ϡ�[���R��4/�c��T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ��fEt7B�_��3E���Y|,�ӟ�c���R��4/�c��T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ��eEx6B�g��3E���Y|,�מ�k���R��4/�c��T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ��cE�4B�w��3E���Y|,���{��#����4+�3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ��bB��2B���3E���Y|,����+����T+�3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ��`B��1B����3E���Y|,����3����T'�3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ��_B��0B����3E���Y|,�����;����T'�3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ��^B��/B����3E���Y|,�������?����T#�3��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ��\B��.B����3E���Y|,������G�R��T�c��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ��ZB��,B����3Er��Y|,������W�R��T�c��T0 k� ������&5AC"3Q �2	4#Q  ��D    ��� ��XB��+B����3Er��Y|,������_�R��T�c��T0 k� �����&5AC"3Q �2	4#Q  ��D    ��� ���WB��*B�×Q�3Er��Y|,������g�R��T�c��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� ���VB��)B�˗Q�3Er��Y|,�#�����o�B��T�c��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� ���TB��(B�ӗQ�3Es�Y|,�+�����w�B����c��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� ���SB��'B�ߘQ�3Es�Y|,�3������B����c��T0 k� ����&5AC"3Q �2	4#Q  ��D    ��� ���RB��&B��Q�3Es�Y|,�;�������B����c��T0 k� �#��'�&5AC"3Q �2	4#Q  ��D    ��� ���OB��$B����3Es#�Y|,�K�r�����B�����c��T0 k� �/��3�&5AC"3Q �2	4#Q  ��D    ��� ���NB��$B����4Es'�Y|,�S�r�����3�S��c��T0 k� �7��;�&5AC"3Q �2	4#Q  ��D    ��� ���MB��#B���4Es/�Y|,�[�r�����3�S��c��T0 k� �?��C�&5AC"3Q �2	4#Q  ��D    ��� ���LB� "B���4Ec7�Y|,�c�r�����3�S��c��T0 k� �3��7�&5AC"3Q �2	4#Q  ��D    ��� ���JB�!B���4Ec;�Y|,�k�r�����3�S��c��T0 k� �/��3�&5AC"3Q �2	4#Q  ��D    ��� ���IB� B����4EcC�Y|,�s������3�S��c��T0 k� �#��'�&5AC"3Q �2	4#Q  �D    ��� ���GB�$B�3���5EcO�Y|,��������3�S��c��T0 k� ����&5AC"3Q �2	4#Q ��O 
   ��� ���FB�,B�;���5H#S�Y|,��������C�C��3��T0 k� �����&5AC"3Q �2	4#Q ��O 
   ��� ���EB�4B�C���5H#[�Y|,������C�C��3��T0 k� ������&5AC"3Q �2	4#Q ��O 
   ��� ���DB�@B�K�A�5H#_�Y|,�������C�C��3��T0 k� ������&5AC"3Q �2	4#Q ��O 
   ��� ���BB�HB�S�A�6H#g�Y|,������C�C��3��T0 k� ������&5AC"3Q �2	4#Q ��O 
   ��� ���@B�\B�g�A�6H#o�Y|,�����C#�C��3��T0 k� ������&5AC"3Q �2	4#Q ��? 
   ��� ���?B�dB�o�A�7H3w�Y|,�����C#�C��3��T0 k� �����&5AC"3Q �2	4#Q ��? 
   ��� ���>B�lB�w�a�7H3{�Y|,�Ô����C'�C��3��T0 k� ���&5AC"3Q �2	4#Q ��? 
   ��� ���=B�tB��a�7H3�Y|,�˔����C'�C��3��T0 k� ���&5AC"3Q �2	4#Q ��? 
   ��� ���<B��B���a�7H3��Y|,�ӕ���'�C'�C��3��T0 k� ���&5AC"3Q �2	4#Q ��? 
   ��� ���;B��B���a�8H3��Y|,�ߕ�#��/�C+����3��T0 k� ���&5AC"3Q �2	4#Q ��? 
   ��� ���:B��B���a�8HC��Y|,���+��7�C+����3��T0 k� �|
��
&5AC"3Q �2	4#Q ��? 
   ��� ���8BѤE���a�8HC��Y|, ���3�BG�S( ���3��T0 k� �d�h&5AC"3Q �2	4#Q ��? 
   ��� �ϸ7BѬE���a�9HC��Y|, ��C7�BO�S( ���3��T0 k� �X�\&5AC"3Q �2	4#Q ��? 
   ��� �ϼ7BѸE���a�9HC��Y|,�C;�BW�S, ��3��T0 k� �L�P&5AC"3Q �2	4#Q ��? 
   ��� ���6B��E�ßa�9HC��Y|,�C?�B_�S, Cw�3��T0 k� �@�D&5AC"3Q �2	4#Q ��? 
   ��� ���5B��E�ˠa�9HC��Y|,�CC�Bg�S, Cs�3��T0 k� �4�8&5AC"3Q �2	4#Q ��? 
   ��� ���4E��E�Ӡa�:HC��Y|,�CG��k�
�, Ck�3� T0 k� �(�,&5AC"3Q �2	4#Q ��? 
   ��� ���2E��E��a�:HC��Y|,3�	�O��{�
�0 C_�3�T0 k� ��&5AC"3Q �2	4#Q ��? 
   ��� ���1E��E��a�:HC��Y|,;�	�S���
�4 CW�3�T0 k� �!�!&5AC"3Q �2	4#Q ��? 
   ��� ���0E��E���a�;HC��Y|,C�	�W����
�4 CO�3�T0 k� ��$� $&5AC"3Q �2	4#Q ��? 
   ��� ���0E� D���a�;HC��Y|,K�	�W����S8 CK�3�T0 k� ��&��&&5AC"3Q �2	4#Q  ��? 
   ��� ���/B�D��a�;HC��Y|,S�	�[��S8 CC�3�T0 k� ��(��(&5AC"3Q �2	4#Q  ��? 	   ��� ���.B�
D��a�;HC��Y|,[�
_��S< C;�3�T0 k� ��*��*&5AC"3Q �2	4#Q  ��? 	   ��� ���,B�$D��a�<HC��Y|,�o�
c�§�S@ C/�3�T0 k� ��/��/&5AC"3Q �2	4#Q  .�? 	   ��� ���,B�,D�'�a�<HC��Y|,�w�
g�«�SD 3'�3�T0 k� �1��1&5AC"3Q �2	4#Q  ��? 	   ��� ���+B�8D�/�a�<HC��Y|,��
g�¯�SD 3�3�T0 k� �4��4&5AC"3Q �2	4#Q  ��? 	   ��� |� *B�@D�7�a�=HC��Y|,���sk�%r��SH 3�3�T0 k� �6��6&5AC"3Q �2	4#Q  ��? 	   �   x�)B�HD�?�a�=HC��Y|,���so�%r��SH 3�3�T0 k� �8��8&5AC"3Q �2	4#Q  ��? 	   �  u�)B�PD�G�a�=Ec��Y|,���so�%r��SH 3�3�T0 k� �:��:&5AC"3Q �2	4#Q  ��? 	   �  r�'B�dD�W�a�>Ec��Y|,���sw�%r��SL 2��3�T0 k� �p?�t?&5AC"3Q �2	4#Q  ��? 	   �  n� 'B�lD�c�a�>Ec��Y|,���sw�%r��SP 2��3�T0 k� �dA�hA&5AC"3Q �2	4#Q  ��? 	   �  k�(&Ct D�k�a|>Ec��Y|,���c{�%r��SP 2��3�T0 k� �XD�\D&5AC"3Q �2	4#Q  �? 	   �  t�0%C�D�s�a|>Ec��Y|,�Þc{�%r��SP B��3�T0 k� �lA�pA&5AC"3Q �2	4#Q ��? 	   �  |�4%C��D�{�a|>Ec��Y|,�˟c�%r��SP B��3�T0 k� �?��?&5AC"3Q �2	4#Q ��? 	   �  ��<$C��Dレa|?Ec��Y|,�ӟc�%r��SP B��3�T0 k� �<��<&5AC"3Q �2	4#Q ��? 	   �  ��D#C��E���Qx?ET�Y|,�۟c��%r��ST B��3�T0 k� �:��:&5AC"3Q �2	4#Q ��? 	   � 	 ��T"I2��E���Qx?ET�Y|,��c��%r��ST 2��3�T0 k� ��5��5&5AC"3Q �2	4#Q ��? 	   � 
 ��\!I2��E���Qx@ET�Y|,��S��%r��ST 2��3�T0 k� ��3��3&5AC"3Q �2	4#Q ��? 	   �  ��d!I2��E���Qt@ET�Y|,	��S��%r��ST 2��3�T0 k� ��0� 0&5AC"3Q �2	4#Q ��? 	   �  ��l I2��E���At@C��Y|,	�S��%r��
�T 2��3�T0 k� �.�.&5AC"3Q �2	4#Q ��?    �  ��tI2��E���At@C��Y|,	�S��%s�
�T 2��3�T0 k� �$,�(,&5AC"3Q �2	4#Q ��?    �  ��|B��EsòAt@C��Y|,	�S��%s�
�T 2��3�T0 k� �8)�<)&5AC"3Q �2	4#Q ��?    �  ���B��Es˳ApAC��Y|,	���%s�
�T 2��3�T0 k� �L'�P'&5AC"3Q �2	4#Q ��?    �  ���B���EsϴApAC��a�,	"���%s�
�T 2��3�T0 k� �`$�d$&5AC"3Q �2	4#Q ��?    �  ���B���Es׵ApAC���a�,	"#���%s�
�T 2��3�T0 k� �t"�x"&5AC"3Q �2	4#Q ��?    �  ���B���Es߶ApAC���a�,	"'���%s�
�T "��3�T0 k� � �� &5AC"3Q �2	4#Q ��?    �  ���B���Es�ApAC���a�,	"/���%s�
�X "��3�T0 k� ���&5AC"3Q �2	4#Q ��?    �  ���B���Es�AlBC���a�,	"3���%��
�X "��3�T0 k� ���&5AC"3Q �2	4#Q ��?    �  ���B���Es�AlBC���a�,	7���%��
�X "��3�T0 k� ����&5AC"3Q �2	4#Q �?    �  � �B���Es��lBAS��a�,	;��{�%��
�\ "��3�T0 k� ����&5AC"3Q �2	4#Q �?    �  � �B���A��lBAS��a�,	C��{�%��3\ "��3�T0 k� ����&5AC"3Q �2	4#Q ��?    �  � �B���A��lBAS��a�,	G��w�%��3` "��3�T0 k� ��&5AC"3Q �2	4#Q ��?    �  � �B���A��lBAS��a�,	K�Sw�%�#�3`"��3�T0 k� ��&5AC"3Q �2	4#Q ��?    �  � �B���A��lBAS��a�,�W�Ss�%�#�3d"�3�T0 k� �@
�D
&5AC"3Q �2	4#Q ��?    �  � �B���A�#�lBAS��Y|,�[�So�%�#�3h��3�T0 k� �T�X&5AC"3Q �2	4#Q ��?    �  � �B���A�+�QlBAS��Y|,�c�So�%�'�3h�{�3� T0 k� �h�l&5AC"3Q �2	4#Q ��?    �  � �B���A�/�QlBAS��Y|,�g�Sk�%s+�3l�w�3� T0 k� �|��&5AC"3Q �2	4#Q $�?    �  �  B���A�7�QlBAS��Y|,�o�Sk�%s+�3l�w�3� T0 k� #|��&5AC"3Q �2	4#Q ��?    �  � B���A�;�QlBAS��Y|,�s�Sg�%s/�Cp�s�3��T0 k� #���&5AC"3Q �2	4#Q ��?    �  � B���A�C�QlBAS��Y|,�{�Sg�%s/�Cp�s�3��T0 k� #���&5AC"3Q �2	4#Q ��?    �  � B���A�G��lBAS��Y|,��Sc�%s3�Cp�s�3��T0 k� #���&5AC"3Q �2	4#Q ��?    �  � B���A�O��lBAS��Y|,���Sc�%s3�Ct�o�3��T0 k� #���&5AC"3Q �2	4#Q ��?    �  � $B���A�S��lBAS��Y|,���S_�%s7�Ct�l 3��T0 k� #���&5AC"3Q �2	4#Q ��?    �  � (B���A�W��lBAS��Y|,���S_�%s7�Cx�l3��T0 k� ����&5AC"3Q �2	4#Q ��?    �  � 0B���A�_��lBAS��Y|,���S[�%s;�Cx�h3��T0 k� ����&5AC"3Q �2	4#Q ��;    �  � 8B���A�c��lBAS��a�,���S[�%s;�C|	�h3��T0 k� �� �� &5AC"3Q �2	4#Q ��;    �  � <B���A�g��lBAS��a�,���SW�%�?�C|
h3��T0 k� ������&5AC"3Q �2	4#Q ��;    �  � DB���A�o��lBAS��a�,���SW�%�?�C|h	3��T0 k� ������&5AC"3Q �2	4#Q ��K    �  � HB���A�s��lBES��a�,B��SS�%�C�C�h3��T0 k� 3�����&5AC"3Q �2	4#Q ��K    �  � TB�  A�{��lBES��a�,B��SO�%�C�C�h3��T0 k� 3�����&5AC"3Q �2	4#Q ��K    �  � \B�  A���lBES��a�,B��SK�%�G�S�h3��T0 k� 3�����&5AC"3Q �2	4#Q ��K    �  � `B� A���lBES��a�,B��CG�%�G�S�h3��T0 k� 3�����&5AC"3Q �2	4#Q ��K    �  � hB� A���lBES��a�,BîCC�%�K�S�h3��T0 k� ������&5AC"3Q �2	4#Q ��K    �  � lB� A���lBEC��a�,BǯC?�%�K�S�h3��T0 k� ������&5AC"3Q �2	4#Q ��K    �  � pB� A����lBEC��a�,B˱C;�%�O�S�l3��T0 k� ������&5AC"3Q �2	4#Q ��K    �  � xB� A����lBEC��Y|,BϲC7�3O�Èl3��T0 k� ������&5AC"3Q �2	4#Q ��K    �  � |B� A����lBEC��Y|,BӳC3�3O�Èl3��T0 k� ������&5AC"3Q �2	4#Q  ��K    �  � �@c A����lBEC��Y|,B۵C/�3S�Èl3��T0 k� #�����&5AC"3Q �2	4#Q  -�K    �  � �@cA����lBE���Y|,B�3+�3W�Èp!3��T0 k� #�����&5AC"3Q �2	4#Q  ��K    �  � �@cA����lBEӿ�Y|,R�3'�3W�Èp#3��T0 k� #�����&5AC"3Q �2	4#Q  ��K    �  � �@cA����lBEӻ�Y|,R�3'�3W���t%3��T0 k� #�����&5AC"3Q �2	4#Q  ��K    �  � �@cA����lBEӷ�Y|,R�3'�3[���t'3��T0 k� �����&5AC"3Q �2	4#Q ��K    �  � �@cA���lBEӳ�Y|,R�3'�3X �� x)3��T0 k� �����&5AC"3Q �2	4#Q ��K    �  � �@cA���lBEӯ�Y|,R�C'�3\ ��!x+3��T0 k� �����&5AC"3Q �2	4#Q ��K    �  � �@cA���lAEӫ�Y|,R�C'�C\��#|-3��T0 k� �����&5AC"3Q �2	4#Q ��K    �  � �@cA���lAEӣ�Y|,R��C+�C`��%�13��T0 k� �����&5AC"3Q �2	4#Q ��K    �  � �@cA���lAEӟ�Y|,R��C+�C`��'"�33��T0 k� C�����&5AC"3Q �2	4#Q ��K    �  � �
@cA���lAEӗ�Y|,R��C+�C`��("�63��T0 k� C�����&5AC"3Q �2	4#Q ��K    �  � �
@cA���lAEӓ�Y|,R��C+�Cd��*"�83��T0 k� C�����&5AC"3Q �2	4#Q ��K    �  � �
@c A���lAEӋ�Y|,b��C/�Cd�|,"�:3��T0 k� C�����&5AC"3Q �2	4#Q ��K    �  � �
@c A���lAE��Y|,b��C/�Cd�|-"�<3��T0 k� C�����&5AC"3Q �2	4#Q ��K    �  � �	@c A���lAE��Y|,b��C/�Ch�|/"�>3��T0 k� �����&5AC"3Q �2	4#Q ��K    �  � �	@c A���lAE�{�Y|,b��C/�Ch	�x0"�@3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � �	@c$A���lAE�w�Y|,b��C/�Ch
�t2"�B3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � �	@c$A���lAE�o�Y|,b��S3�Cl�t3"�D3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � �@c$A���lAA�k�Y|,b��S3�Sl�p5"�F3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � �@c(A���lAA�_�Y|,b��S3�Sp�l8"�J3��T0 k� #�����&5AC"3Q �2	4#Q  /�K    �  � �@c(A���lAA�[�Y|,b��S3�Sp�h:"�L3��T0 k� #�����&5AC"3Q �2	4#Q  ��K    �  � �@c,A���lAA�S�Y|,b��S3�Sp�h<"�N3��T0 k� #�����&5AC"3Q �2	4#Q  ��K    �  � �@c,A���lAA�O�Y|,r��S3�St�d="�P3��T0 k� #�����&5AC"3Q �2	4#Q  ��K    �  � �@c,A���lAA�K�Y|,r��S/�St�`?"�R3��T0 k� #�����&5AC"3Q �2	4#Q  ��K    �  � �@c,A���lAA�G�Y|,r��S/�St�\A"�T3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � �@c0A���lAA�C�Y|,r��S/�Sx�XC�V3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @c0A�{��lAA�;�Y|,r��S+�Sx�TF�Y3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @c0A�{��lAA�;�Y|,r���+�cx�PH�[3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @c4A�{��lAA�7�Y|,r���'�c|	sLJ�]3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @c4A�{��lAA�3�Y|,r���'�c|!	sHK�_3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @c4A�{��lAA�3�Y|,r���'�c|#	sHM��a3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @c4A�w��lAA�3�Y|,r���#�c|$	sDN��b3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @c8A�w��lAA�3�Y|,B���#�À&	sDO��d3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @c8A�w��lAA�/�Y|,B���#�À(	�@Q��f3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @c8A�w��lAA�/�Y|,B����À*	�@R��h3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  �  @c8A�w��lAA�/�Y|,B����À,	�<S��i3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � $@c<A�w��lAA�/�Y|,B����À.	�<T��k3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � $@c<A�s��l@A�/�Y|,B����À0	�8U��l3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � (@c<A�s��l@A�/�Y|,B����À2	s8V��n3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ,@c<A�s��l@A�+�Y|,B����À4	s8W��p3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � 0@c<A�s��l@A�+�Y|,B�����|6	s8X��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � 0@c@A�s��l@A�+�Y|,�����|8	s8Y��s3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � 8@c@A�s��l@A�'�Y|,�����|<	s4[�v3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � 8@cDA�o��l@A�'�Y|,�����x>	�4\�w3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � <@cDA�o��l@A�'�Y|,��
���x@	�4\�x3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @@cDA�o��l@A�'�Y|,�����tB	�4]�z3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � @@cDA�o��l@A�'�Y|,�����tD	�4^�{3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � D@cHA�o��l@A�#�Y|,�����tG	�4^�}3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � H@cHA�o��l@A�#�Y|,�����pI	s4_�~3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � H@cHA�o��l@A�#�Y|,�����pK	s4_�3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � L@cH	A�o��l@A�#�Y|,�����lM	s4`� �3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � L@cL	A�k��l@A��Y|,�����hO	s4`�$�3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � P@cL	A�o��l@A��Y|,�����hQ	s4`�$�3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � T@cL
A�o��l@A��Y|,�����dS	�4a�(�3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � T@cL
A�o��l@A��Y|,�����`U	�4a�,3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � X@cP
A�o��l@A��Y|,�����`U	�4b�03��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � X@cP
A�o��l@A��Y|,�����`U	�0b�03��T0 k� �����&5AC"3Q �2	4#Q  ��K   �  � \@cPA�s��l@A��Y|,�!���`V	�0c�43��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � \ @cPA�s��l@A��Y|,�#���`W	s,d�8~3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ` @cTA�s��l@A��Y|,�$���`X	s,d�<~3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ` @cTA�s��l@A��Y|,�&���\Y	s(e�<~3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � d @cTA�s��l@A��Y|,�'���\Z	s(f�@}3��T0 k� �����&5AC"3Q �2	4#Q  ��K   �  � d @cTA�w��l@A��Y|,�)���\[	s$f�D}3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � h @cTA�w��l@A� Y|,�*���X\�$g�D}3��T0 k� �����&5AC"3Q �2	4#Q  ��K   �  � h @cXA�w��l@A� Y|,�,���X]�$g�H}3��T0 k� �����&5AC"3Q �2	4#Q  ��K   �  � l @cXA�w��l@A� Y|,�-���X]� h�L|3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � o�@cXA�w��l@A�Y|,�/���X^� h�L|3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � s�@cXA�w��l@A�Y|,�0���T_�i�P|3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � s�@cXA�{��l@A�Y|,�1����T_�j�P|3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � w�@c\A�{��l@A�Y|,�3����P_�j�T{3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � w�@c\A�{��l@A�Y|,�4����P`�k�X{3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � {�@c\A�{��l@A�Y|,�5����L`�k�X{3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � {�@c\A�{��l@A�Y|,�7����L`�l�\{3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � {�@c\A�{��l@A�Y|,�8����H`�l�\z3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � �@c`A�{��l@A�Y|,�9����H`m�`z3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � �@c`A���l@A�Y|,�:����D`m�`z3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c`A���l@A�Y|,�<����D`n�dz3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c`A���l@A�Y|,�=����@`n�dz3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c`A���l@A�Y|,�>����@`o�hy3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c`A���l@A�Y|,�?����@`o�hy3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cdA���l@A�Y|,�@����@`p�ly3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cdA���l@A�Y|,�A���S<`p�ly3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cdA���l@A�Y|,�B���S<`q�py3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cdA���l@A�Y|,�C���S<`q�px3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cdA���l@A�Y|,�E���S8`r�tx3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cdA���l@A�Y|,�F���S8` r�tx3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@chA���l@A�Y|,�G���S8` s�xx3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@chA���l@A�Y|,�HB��S8` s�xx3��T0 k� �����&5AC"3Q �2	4#Q  ��K   �  � ��@chA���l@A�Y|,�IB��S8`�s�|w3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@chA���l@A�Y|,�JB��S4`�t�|w3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@chA���l@A�Y|,�KB��S4`�t��w3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@chA���l@A�Y|,�LB��S4`�u��w3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@chA���l@A�Y|,�LB��S4`�u��w3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@chA���l@A�	Y|,�MB��S0`�u��w3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@clA���l@A�	Y|,�NB��S0`�v��v3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@clA���l@A�
Y|,ҘOB��c0`�v��v"���T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@clA���l@A�
Y|,ҘPB��c0`�w��v"���T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@clA���l@A�
Y|,ҔQB��c0`�w��v"���T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@clA���l@A�Y|,ҔRB��c,`�w��v"���T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@clA���l@A�Y|,ҔSR��c,`�x��v"���T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@clA���l@A�Y|,ҔTR��c,`�x��v"���T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@clA���l@A�Y|,B�TR��c,`�x��u"���T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cpA���l@A�Y|,B�UR��c,`�y��u"���T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cpA� �l@A�Y|,B�VR��c(`�y��u"���T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cpA� �l@A�Y|,B�WR��c(`�y��u"���T0 k� �����&5AC"3Q �2	4#Q  ��K   �  � ��@cpA� �l@A�Y|,B�XR��c(`�z��u"���T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cpA� �l@A�Y|,B�YR��c(`�z��u3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cpA� �l@A�Y|,B�[R��c(`�z��u3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cpA� �l@A�Y|,B�\R� c(`�{��t3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cpA� �l@A�Y|,B�]R�c$`�{��t3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@ctA��l@A�Y|,"�_b�c$`�|��t3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@ctA��l@A�Y|,"�ab�c$`�|��t3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@ctA��l@A�Y|,"�bb�c$`�|��t3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@ctA��l@A�Y|,"�cb�c$`�|��t3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@ctA��l@A�Y|,"�eb�c `��}��t3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@ctA��l@A�Y|,"�fb�c `��}��t3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@ctA��l@A�Y|,"�gb�c `��}��s"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@ctA��l@A�Y|,"�ib�c `��~��s"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@ctA��l@A�Y|,"�jb�	c `��~��s"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@ctA��l@A�Y|,"�lb�	c `��~��s"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,�mr�
c `��~��s"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,�or�c`��~��s"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,�pr�c`����s"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,�qr�c`����s"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,�sr�c`����s"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,�tr�c`����r"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,�ur�c`����r"s��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,�vr�c`R���r3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,�vr�c`R���r3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,�vr�c`R���r3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A�Y|,��vr�c`R����r3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@cxA���l@A� Y|,��wB�c`R���r3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A� Y|,��xB�c`����r3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A�!Y|,��xB�c`����r3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A�"Y|,��yB�c`����r3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A�"Y|,��yB�S`��~��r3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A�#Y|,��yB�S`��~��r3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A�#Y|,��yB�S`��~��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A�$Y|,��zB� S`��}��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A� %Y|,��z2�"S`��}��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A� %Y|,Ҭz2�#S`��|��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A� &Y|,Ҭz2�%S`��|��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K   �  � ��@c|A���l@A� &Y|,Ұz2�'S`��{��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A� 'Y|,Ұ{2�)S`��{��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A�$'Y|,Ұ{2�+�`��z��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c|A���l@A�$(Y|,r�{2�,�`��y��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�$)Y|,r�{2�.�`��x��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�$)Y|,r�{2�0�`��x��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�$*Y|,r�|"�2�`��w��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�$*Y|,r�|"�4�`��v��q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�(+Y|,r�|"�6�`��u �q3��T0 k� �����&5AC"3Q �2	4#Q  ��K   �  � ��@c�A���l@A�(+Y|,r�|"�8�`��t �q3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�(,Y|,r�|"�:�`� s �p3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�(,Y|,r�|"�<�`� r �p3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�(,Y|,r�}"�>�`� q �p3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  � ��@c�A���l@A�,-Y|,��}"�@�`�p��p3��T0 k� �����&5AC"3Q �2	4#Q  ��K    �  �                                                                                                                                                                            � � �  �  �  d A�  �K����   �      6 \�� ]�'�'� � �
����          � ��-    ���� ��|    �� �              `           �0     ���   0
&


          "Z        � �fL     � �^     � |               	�� �         �@     ���   0	
           ��         �j     �z�~     ��,                � �         ��     ���   (
 
           @B�          [%1     @B� [%1           
           !   J           ��     ���   H	$
          ;��    	    / �^�     ;� �G�    �Z                
   �j          �0     ���   03 
           � �	      C���     ����                            ���d                ���   P		 5              }�P  � �    W ��4     }�� ��    �� �           ? Z �         ���    ��`  8	 

          ]�:  � �
	   k �rj     ]�� �a�     � �           s Z �         ���  &  ��`  8
)           ]��    	    ���     ]�� ���                    4		 Z �         �     ��@   (
	           p��  � �	    � Ö�     p�+ �h�    9�             S	 Z �         	 ��    ��`  0
3
          Xˣ  @ @     � ��n     YC^ ���    ���            > Z �         
 ��    ��@  H


         ���� ��     � �{    ���� �{                            �� �              l  ��H    		 5 	                 ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��ye  ��        � �ZP    ��ye �ZP         "                 x                j  �       �                         ��    ��       � �      ��   �           "                                                 �                          � � [ �� � � � � � ��� � �  	              
 
  ;    � �� �H�O       �$ �m` �$ n` �D n� �d n� Є n� Ф n� &� u����X � B� v  ̄ 0p� �� p� � 0q  ��  w` �$ �w� �d  x� <�  u� �d  x� פ y  �� `w� τ x@ D� `[� E�  \� E�  \� 
�\ X  �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ���� ����� ����� � � b  � �j� �  k� �� 0[� �D  \@ ̄ 0\� �� \� � 0]  �d �o� �d p� � �c` � d` � �w` � 0x` �d  x� פ y   � �r` � s` (� `^` )D  _   � �t� � u� �$  }� �d  }����� � 
�\ W  
�\ W� 
�< W� 
�\ X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���� �  ���7  ������  
�fD
��L���"����D"� �  " `   J jF��    "�j "���
��
���     �j��  
  �
� �  �  
� ��   ��     � �       ;    ��     � �      ��   ��     � �          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �K 53 5      ��7T ���        � � �  ���        �        ��        �        ��        �   >�     
���/��        ��                         T�) , ����� �                                      �                 ����           �� ����&��    � 2  �            9 Pelle Eklund e                                                                                   5  4     �GC,\ C#$ �B� � �cWi �c_a � cbY �ccQ �ckH � 	csP � 
ct@ � cu@ � cvK � cwF �c�a �c�b �c�Z � c�i �c�X �cI � c�A �K/% � K75 �J� �J� � � � � � � � �c� � �c� � �c� � � c� � �c�H �  c�X � !c�P �	"� � �	#� � �$� � �%� �&K � � 'K �("� � � )"� � �*� � �+
� � �,"�$ � -"�6 �."�  �/*�/ �0"� � � 1"� � �2� � �3
� � q  *R} � 
� � q  *R} �7� � �8
� � q  *R}; :"J �K ;"Q �S <"P �[  "I �@  *Gz(  *Kr                                                                                                                                                                                                                         �� P         �     ` 
             \ P E _  ��                    ������������������������������������� ���������	�
���������                                                                                          ��    ��e�� ��������������������������������������������������������   �4, H� 0 8�� }�� �A A ���&��.����U�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   3    "    �� ��J       �  	                           ������������������������������������������������������                                                                      	                                                                    ����  ��                                             �������������������� � ������ ���� ��� �������������������������� ���������������� ������������������� ���������� ��������������� �������������������������������������������   ������ ����� ���������������� ������������ ���������                           	        K    '     �� 
ĳJ      �}                             ������������������������������������������������������                                                                                                                                      �3R���  �                                           ����� ���� �� ����������� �� ����� ������������������� ���� ��������������������������� � ��������������� ���������� ��� � ������� ������������������������ �������������������������������� ���� ���� �������������������������                                                                                                                                                                                                                                                               	                                                           �              


            �   }�         ����  6�  6�  0�����  �  V����������������������������������������������������������������������������      Z          HF  Z     8�                                                      ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � �� �m`                                                                                                                                                                                                                                                                                          E)n1n  �                                      m      b                                                                                                                                                                                                                                                                                                                                                                                                              
 �  
>�  J�  (�  (�  J`�  ��H�L�˶��̎����� ���d�2���������������̿                 x � : ���       $   �   &  QW  �   �                    �                                                                                                                                                                                                                                                                                                                                        K K   �               "         !��                                                                                                                                                                                                                        Z   �� �~ ��      �� m      �������������������� � ������ ���� ��� �������������������������� ���������������� ������������������� ���������� ��������������� �������������������������������������������   ������ ����� ���������������� ������������ �������������� ���� �� ����������� �� ����� ������������������� ���� ��������������������������� � ��������������� ���������� ��� � ������� ������������������������ �������������������������������� ���� ���� �������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     2      2   � ��                       B     �   �����J���J'      ��     p      �      �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��    �� � �� �� �z � � �N ^$     �(        �� ��  � ��     � ��   	 ��   p �� �� �z   p���� �$    ��s �������s  ��   0 ����  �� �� �  ��   ��     ��   � �� ��      � �N ��   ' �� K �� ��   	 ��  �� �� m` �� �� �z m` �$ �$ r  ��r       �      �������2����  g���        f ^�         ��b             ��v���2�������J��~T���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                                                  U  T   T   T     T UDUDDUDDDDDDDDDDDDDDDP   E�  DU� DDU�DDDUDDDDDDDDDDDD                UP  E�  E   E                                           ���U�UTD�DDDDDDTDD TDD   �   U_ DEU�DDDUDDDDD��DZT�DDDDDDDDDDDDTDDDDDDDDUTU�����DDDDDDDDDDDEDDDEDDDDTUTU�Ԫ���Z_   P   � �U�UTDUDDDDUTD�DT��D        U_��DEU_DDD_DDDPDDE�DDE  �DD DD DD �DD �UD  �U       DZTDEDDDDE�DDE�DDE�TDDT�DE�TE���DDTU�ZD���������DDTDD��ZT�T���ZTDDE��D��T�T��DUTTT��Z��TQTDDUTD�DDDTDDD�DDDDDDE�DD_TDE�DD_ DDP DDP DD_ DU_ U�  �                                       TE�DDD�UUU                    ���DDDUUUTD  D  D  D  D  U��D�TDDDDEUUDP  DP  DP  DP  UP  TDE�DDDPUUU_                                                    wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwtwwwCwwt1wwCwt1wC�t1��C1����������""""���������������!���""!����,���ww��7����������������wwwwwwwwwwwwwwwwwwww7wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwws��w1wt1�wC�t1��s��s��s������"$��Gw�!������������L���q��"r��������!�����!ww�r�w�ww!�wwrwwwwwwqwwwrwwww�7ww�ww�ww��7w��w���G��'!wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  " ! " "" """ "!   " ""                                                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  " ! " ""  "!  " ! " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  " ! " "" """ "!   " ""                                                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �              "      �              "   "   "�  �                            �   ��  �ڛ�}ک�"   "   "  �� ��                   �".��".���                                ".  ".  ���                                                                                                                                                                                                                        	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           "� /���  �       �   �   �                                                   ��                     �   �                      �".��".  ���    �    �   �   �   D   E�  U�  UO                         "  "  "                                                                                                                                                                �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���        T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ��"� �"� ����                        �   ��  "   "   �   "  "  "   �                                 �   ���                            �   "                                                                                                  �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���                            .   .   �             �  "� "  "  "  �                         �                 ��"� �"� ����                            ".  ".  ���   ���� �                                                                                                                                                                                        �� ��� ��� ww� &'� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                               " "/ �/� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   �".��".���                                        � ��       "   "   "�  �                            �   ���                            �   "                                                                                                         �  �  �  �  w  �  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �   ؛  �(� !"� "/ !/� "� �    ��   �   �   �          �        �!� �                                                                                                                                         �  �  "   "                                                                     �� ̽ ̽��۽ }�  wz  � ��������ɜ���̚��̸ ��  ��  �  �  T�  T�  H� �E �E �D�[ ˻  ˸  ��  
� ,"�"" �"  �"              "   *�  ��� ��� �ة��ڋ�̽� ��  ��  ̻� ̻� ��� ��@ ��@ DD0 T30 B3� ��  ��  ��  
� +� �"" �"� �" ��� ����  ��          ���    �                       
 "� ""� ""� "                       �                             ���                         �"  �"                    ���.�                                            "  "  "                            ���                          ����                  �   �� �       �  �  "�  "   "                                                  �  �  �  �� ݚ� }�Ȫ��˙������˼� ��  ��  ��  ��  ��  I� H� �E X�T X�S T�D �[ ˻  ˸  ��  
� �,"��"" "  �" �  ""� �� ˻ �˻ ��ݪ��کɨ��ˀ�̽ ��� ��  ̽  ̻  ̻  ˉ  ��  �D  DC  C3  #;  ;�� �� ��  �� "�  "  �"/ / ����� ��  �      �   �          �  �  "     "  "  "   "�  �  �   �   
                            �          �   �          �                    �   �".� .�    ���.�                                  �  �˰ ��� �wp �&                                                                                                                                                                 �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���                              "  "             ��.�  .                 ����                         � "            � "�",�"+� ",                       "  .���"    �     �                         � ".��".��/����  �                                �   "                                                                                                   ۻ� ۽� ��� H�DH�D�DP�E X�T H�P H�@ Ȥ� ̻� ˘ �� "*� �/�""/""/���                       ��  ۼ� ݻ� w�� b}ذgvz�w������ɨ�ͨ���ڋ��٭���ۻݻ� �   �          �   �   .   ."  ""  ""  ,   �   
            "  "  ""  "�   �           �   ��  �      �                                     .  .     "   "  "                     �   �   �             � � "            � "�",�"+� ",                       "  .���"    �     �                           ""  "".  . �    �                                                                                                                                       	�� ��� ��� ��� ��r ��g �۶ �� ��  -�  �8 
3� D> 	D3 �C0˳ "+  ""  "   ��  �  ��  �  ��   ��  ��  wڐ bک g���w����ə�ͼ���܈��;��33̽�B��N�+0 ""@ B�  B$� K� ȋ  ʠ  +   "  �"" "�             �  "� "  �   �   �� ��� ��       �                     �  "� "     �   �     "  "  "                       �  ��  ��  ww  &'  vv  w                �                        ��"� �"� ����                         " "" "�  ��                        ����                               ���                          ����                  �   �� �       �  �  "�  "   "                                                                    �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ���������""��""��""�����        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                   �       �   �   �                                                                                                                                                                                      2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ DD D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD l � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������  � �!�aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� X � �!�aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w � �!�aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww���������������� � � �!�aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� L  . M + , N    O P Q R S S S T S S S T S S 0 Z S ST S S ST S S SRQPO(( (N(,(+(M(.L����������������  7  N 5 U V W X Y S S [ S S S _ S S S _ S S \ ] S S_ S S S_ S S S[ S SY(X(W(V(U(5(N((7����������������  `  V    a b c S S f g h i j i i i j i i ^ d i ij i i ij ihgf S Scb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � �� � � � � � ���	����� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � �� ��������� � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � � �������� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � � ���� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � ��	� � � ��� � � � � � � � � � � ��	� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w � � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� � � � i i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� W � � u u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� a � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(�����������������  � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������LDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDDGC,\ C#$ �B� � �cWi �c_a � cbY �ccQ �ckH � 	csP � 
ct@ � cu@ � cvK � cwF �c�a �c�b �c�Z � c�i �c�X �cI � c�A �K/% � K75 �J� �J� � � � � � � � �c� � �c� � �c� � � c� � �c�H �  c�X � !c�P �	"� � �	#� � �$� � �%� �&K � � 'K �("� � � )"� � �*� � �+
� � �,"�$ � -"�6 �."�  �/*�/ �0"� � � 1"� � �2� � �3
� � q  *R} � 
� � q  *R} �7� � �8
� � q  *R}; :"J �K ;"Q �S <"P �[  "I �@  *Gz(  *Kr3333DDDDAqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD��������������������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ��������������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ��������������������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE��������������������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD��������������������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD��������������������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD��������������������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� ����7�\�J��<�V�I�P�[�H�P�S�S�L�������8�>�7���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� ��!��-�V�I��0�Z�Z�L�U�Z�H����������8�>�7���""""������A�D��I��""""�������D����� ��%��:�L�S�S�L��0�R�S�\�U�K���������8�>�7���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �8�>�7���!���A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �>��<�����""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,�����������DDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �����<�L�Z�\�T�L��2�H�T�L����������������� ����4�U�Z�[�H�U�[��<�L�W�S�H�`��������������� ����.�O�H�U�N�L��2�V�H�S�P�L���������������� ������0�K�P�[��7�P�U�L�Z��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 