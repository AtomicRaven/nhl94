GST@�                                                            \     �                                               9    ��              
      ����e �	 J�����������`���z���        �h     #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"��   " `  J  jF��     �j  
 ���
��
��    "�j��" " ��
   �                                                                              ����������������������������������      ��    bb? QQ0 5 118 44               		 


     
               ��� 4    �                 nnY ))         88:�����������������������������������������������������������������������������������������������������������������������������=  0b  4  11                                         �  �  �  �                  �  
          = �����������������������������������������������������������������������������                                (  ;   �  ��   @  #   �   �                                                                                '      )n)nY  
�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    dR@��3�d�,K���|,�#�B�0eE/��	�$E�Z3�T0 k� �"��"	E1 4#Q&�1D"3Q  $�    � < �dQ@r�1�l�4K���|,�+�B�8eE/��	�#E�Z3�T0 k� � �� 	E1 4#Q&�1D"3Q  ��    � < ��dO@r�0�t�<K��|,�3�B�@eE/��	�#E�Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��    � < ��dM@r�/�|�@K��|,�;�B�LeE��	�"E�Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��    � < ��hL@r�.���HK��|,�C�B�TdE��!A��Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��    � < ��hH@r�,���XK�#�|,�W�B�ddE�� A��Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��    � < ��lG@r�+���\K�+�|,�_�ClcE�� A��Z3�T0 k� ����	E1 4#Q&�1D"3Q  ��    � < ��lE@r�)���dK�3�|,�g�CtcE��$A��Z3�T0 k� � �	E1 4#Q&�1D"3Q  ��    � < ��pC@r�(���lK�;�|,�o�C|cE��(E� Z3�T0 k� ��	E1 4#Q&�1D"3Q  ��    � < ��pB@r�(���tK�C�|,�w�C�bB����0E� Z3�T0 k� ��	E1 4#Q&�1D"3Q  ��    � < ��t@@r�'���|K�K�|,��C�bB����4E� Z3�T0 k� ��	E1 4#Q&�1D"3Q  ��    � < ��x?E�&����K�S�|,߇�E��aB����<E�!Z3�T0 k� ��	E1 4#Q&�1D"3Q  ��    � < ��|<E%����K�c�|,ߗ�E��`B����DE�"Z3�T0 k� � �$	E1 4#Q&�1D"3Q  ��    � < ���:E$����K�k�|,ߟ�E��`E���LE�#Z3�T0 k� �$�(	E1 4#Q&�1D"3Q  ��    � < ���9E#����K�s�|,߫�E��`E��PF�#Zc�T0 k� �(�,	E1 4#Q&�1D"3Q  ��    � < ���7E"����K�{�|,߳�E��_E��TF�$Zc�T0 k� �,�0	E1 4#Q&�1D"3Q  ��    � < ���6E !�� ��K���|,߻�E��^E��\F�%Zc�T0 k� �4!�8!	E1 4#Q&�1D"3Q  ��    � < ���4E(!� ��K���|,�ìE��^E��`F�%Zc�T0 k� �<!�@!	E1 4#Q&�1D"3Q  ��    � < ���3FC0 � ��K���|,�ˬE��]E��dF�&Zc�T0 k� �H!�L!	E1 4#Q&�1D"3Q  ��    � < ���0FC0 � ��K���|,�۫E��\E��pF�(Zc�T0 k� �X!�\!	E1 4#Q&�1D"3Q  ��    � < ���/FC4 �( ��K���|,��E��[E��tE��)Zc�T0 k� �`!�d!	E1 4#Q&�1D"3Q  ��    � < ���.FC<�3���K���|,��E��ZE��|E��)Zc�T0 k� �d!�h!	E1 4#Q&�1D"3Q  ��    � < ���-FC@�;���K���|,���E� YE���E��*Zc�T0 k� �l!�p!	E1 4#Q&�1D"3Q  ��    � < ���+FCH�C���K���|,���E�XE�˾�E��+Zc�T0 k� �p!�t!	E1 4#Q&�1D"3Q  ��    � < ���*FCL�K���K���|,��E�WE�Ͻ�E��,Zc�T0 k� �x �| 	E1 4#Q&�1D"3Q  ��    � < ���)FCT�S��K���|,��CBVE�ӻ�E��-Zc�T0 k� �| �� 	E1 4#Q&�1D"3Q  ��    � < ���(FCX�[��K���|,��CBUE�׺�E��-Zc�T0 k� ���	E1 4#Q&�1D"3Q  ��    � < ���%FCd�o��K���|,�'�CB,SE�۸	�E��/Zc�T0 k� ���	E1 4#Q&�1D"3Q �    � < ���$FSh�w�� K���|,�/�CB0QE�߷	�E��0Zc�T0 k� ���	E1 4#Q&�1D"3Q ��    � < ���#FSp���(K��|,�;�CB8PE��	�E��1Zc�T0 k� ���	E1 4#Q&�1D"3Q ��    � < ���"FSt����0K��|,�C�CB@OE��	�
E��2Zc�T0 k� ����	E1 4#Q&�1D"3Q ��    � < ���!FSx����8K��|,�K�CBDMD��	�
E��3Zc�	T0 k� ����	E1 4#Q&�1D"3Q ��    � < �� FSx����@K��|,�S�CBLLD��	�
Er�4Zc�	T0 k� ����	E1 4#Q&�1D"3Q $�    � < ��Fcx����HK�'�|,�[�CBTJD���
�	Er�5Zc�
T0 k� #���	E1 4#Q&�1D"3Q ��    � < �Fcx����XK�;�|,�k�CB`GD���
�Er�7^�
T0 k� #���	E1 4#Q&�1D"3Q ��    � < �Fcx����`K�C�|,�s�CRdFD��
�Er�9^�
T0 k� #���	E1 4#Q&�1D"3Q ��    � < �Fc|����hK�K�|,��CRlED��
�Er�:^�
T0 k� #���	E1 4#Q&�1D"3Q ��    � < � Fc�����pK�S�|,���CRlED���Er�:^�
T0 k� #���	E1 4#Q&�1D"3Q ��    � < �(Fc�����xK�[�|,���CRpDD���Er�;^�T0 k� ����	E1 4#Q&�1D"3Q ��    � < �0Fc����ހK�c�|,���CRpCD���Er�<^�T0 k� ����	E1 4#Q&�1D"3Q ��    � < �8Fc����ވK�o�|,���CRtBD���Er�=^�T0 k� ����	E1 4#Q&�1D"3Q ��    � < �@Fc��� ސK�w�|,���CRtAD�#��Er�=^�T0 k� ����	E1 4#Q&�1D"3Q ��    � < �PFc��� ޠK��|,���CRx?D�/���Er�?^�T0 k� ����	E1 4#Q&�1D"3Q ��    � ; �XFc�� ިK��|,�åCRx>D�3���Eb�@^�T0 k� 3���	E1 4#Q&�1D"3Q ��    � : �`Fc��ްK��|,�ˤCR|=D�;���Eb�A^�T0 k� 3���	E1 4#Q&�1D"3Q ��    � 9 �hFc��޸K��|,�ӤCb|<D�?���Eb�B^�T0 k� 3���	E1 4#Q&�1D"3Q ��    � 8 �pFc�� ��K��|,�ۤCb�;D�G���Eb�C^�T0 k� 3���	E1 4#Q&�1D"3Q ��    � 7 �xFc��(��K	��|,��Cb�9E�K���Eb�D^�T0 k� 3���	E1 4#Q&�1D"3Q ��    � 6 ҀFc�0��K	��|,��Cb�8E�S���I��D^�T0 k� ����	E1 4#Q&�1D"3Q ��    � 5 ҈Fc�8��K	��|,��Cb�7E�W���I��E^�T0 k� ����	E1 4#Q&�1D"3Q ��    � 4 ��Fc�@��K	��|,���Cb�5E�_���I��F^�T0 k� ����	E1 4#Q&�1D"3Q ��    � 4 ��Fc�P��J	��|,	�E��3E�k���I��G^�T0 k� ����	E1 4#Q&�1D"3Q ��    � 4 ��
E��X��J	/��|,	�E��1E�o���I��G^�T0 k� #���	E1 4#Q&�1D"3Q  ��    � 4 ��	E��`��J	/��|,	�E��0E�w�C�I��H^�T0 k� #���	E1 4#Q&�1D"3Q  -�    � 4 ��	E��h�J	/��|,	#�E��.E��C�I��H^�T0 k� #���	E1 4#Q&�1D"3Q  ��    � 4 ��E��h�I	/��|,	+�E��,E���C�I� I^�T0 k� #���	E1 4#Q&�1D"3Q  ��    � 3 ��E��l�I	/��|,	/�E��+E���C�I� I^�T0 k� #���	E1 4#Q&�1D"3Q  ��    � 3 ��O��p�I	��|,	!7�E��)Ep��C�I�I^�T0 k� ����	E1 4#Q&�1D"3Q ��    � 3 ��O��x	�,H	��|,	!C�E��%Ep����I�J^�T0 k� ����	E1 4#Q&�1D"3Q ��    � 3 ��O��|
	�4H	�|,	!K�E��$Ep����I�J^�T0 k� ����	E1 4#Q&�1D"3Q ��    � 3 ��O��|	�8H	�|,	!O�E"Ep����I�J^�T0 k� ����	E1 4#Q&�1D"3Q ��    � 3 ��O���	�@H	 �|,	S�E Ep���� A�J^�T0 k� C���	E1 4#Q&�1D"3Q ��    � 3 � O� ��	�DH	 �|,	[�EEp���� A�K^�T0 k� C���	E1 4#Q&�1D"3Q �    � 3 �O�#���TH	 �|,	c�EEpós��A�K^�
T0 k� C���	E1 4#Q&�1D"3Q �    � 3 � O�$���XH	 �|,	k�EA�˴s��A�K_t 
T0 k� C���	E1 4#Q&�1D"3Q ��    � 3 �  O %���`H�#�|,	!o�EA�ϵs��FL_t 
T0 k� ����	E1 4#Q&�1D"3Q ��    � 3 �3�O'���lH�/�|,	!w�EA�۶s��FL_t 
T0 k� ����	E1 4#Q&�1D"3Q ��    � 3 �;�O)C��tG�3�|,	!{�EA�����FL_t 
T0 k� ����	E1 4#Q&�1D"3Q ��    � 3 �C�O*C��|G�;�|,	!��A�A�����FL_t 
T0 k� ����	E1 4#Q&�1D"3Q ��    � 3 �K�O+C���G�?�|, ��A�A�����FM_t 
T0 k� #�
��
	E1 4#Q&�1D"3Q  ��    � 3 �W�O ,C���G�C�|, ��A�A�����BCM_t 
T0 k� #�	��		E1 4#Q&�1D"3Q  ��    � 3 �_�O$-C���G�K�|, ��A�A������BC M_t 	T0 k� #���	E1 4#Q&�1D"3Q  ��    � 3 �g�O(.C���G�O�|, ��A�	A������BC M_t 	T0 k� #���	E1 4#Q&�1D"3Q  ��    � 3 �o�O0/C���G�W�|, ��A�A�����BC$M_t 	T0 k� #���	E1 4#Q&�1D"3Q  /�    � 3 ��O81C�!��G�c�|, ��A�A�����BC$N_s�	T0 k� ����	E1 4#Q&�1D"3Q  ��    � 3 ���O<2C�"��G�k�|, ��A�A�����BC(N_��	T0 k� ����	E1 4#Q&�1D"3Q  ��    � 3 ���O@3C�$��G�o�|, ��A�A�����BC(N_��	T0 k� ����	E1 4#Q&�1D"3Q  ��    � 3 ���OH4C�&��G�w�|, ��A� A�����BC(N_��	T0 k� ��
��
	E1 4#Q&�1D"3Q  �    � 3 ���FL5S�(��G��|, ��A��A�����BC,N_��	T0 k� ����	E1 4#Q&�1D"3Q  ��    � 3 ���FP6S�)��G���|, ��A��A�#����Es,O_��	T0 k� ����	E1 4#Q&�1D"3Q ��    � 3 ���FT7S�+��G���|, ��A��A�+����Es,O[s�	T0 k� ����	E1 4#Q&�1D"3Q ��    � 3 C��F`9S�/��G���|, ãA��A�3���Es0P[s�	T0 k� ���	E1 4#Q&�1D"3Q ��    � 3 C��E�d:S�1��G���|, ãA��A�7���Es0P[s�	T0 k� ���	E1 4#Q&�1D"3Q ��    � 3 C��E�l;S�3� G���|, ǣA��A�;���Es4Q[s�
T0 k� � �� 	E1 4#Q&�1D"3Q ��    � 3 C��E�p;S�5�F���|, ˣA��A�?���Es4Q[��
T0 k� �#��#	E1 4#Q&�1D"3Q ��    � 3 C��E�t<S�7�F���|, ϣA��A�C���Ec4R[��
T0 k� �&��&	E1 4#Q&�1D"3Q ��    � 3 ���E�x=S�9�F���|, ӣA��A�G���Ec4R[��T0 k� �)��)	E1 4#Q&�1D"3Q ��    � 3 ���@|>S�;� F���|, ףA��A�K���Ec8S[��T0 k� �,��,	E1 4#Q&�1D"3Q ��    � 3 ���@|?c�=�(F���|, ۣA��A�O���Ec8T[��T0 k� �0��0	E1 4#Q&�1D"3Q ��    � 3 ���@|@c�?�0F���|, ߣA��A�S���Ec8T[��T0 k� �3��3	E1 4#Q&�1D"3Q ��    � 3 ���@|Ac�A�8F���|, �A��A�W���Ec8U[� T0 k� �6��6	E1 4#Q&�1D"3Q ��    � 3 ���@xAc�C�@F���|, �A��A�[���ES8V[� T0 k� �9��9	E1 4#Q&�1D"3Q ��    � 3 ���@xBc�E�HF���|, �A��A�_���ES8W[� T0 k� �<��<	E1 4#Q&�1D"3Q ��    � 3 �� @xCc�G�PF���|, �A��A�c���ES8W[tT0 k� �?��?	E1 4#Q&�1D"3Q ��    � 3 �� @tDc�I�XF���|, �A��A�g���ES4X[tT0 k� �B��B	E1 4#Q&�1D"3Q ��    � 3 ��@tE	S�K�`F��|, �A��A�k���ES4Y[tT0 k� �E��E	E1 4#Q&�1D"3Q  ��    � 3 3�@tE	S�M�hF��|, �A��A�o���ES4Y[tT0 k� �I��I	E1 4#Q&�1D"3Q  ��    � 3 3�@tF	S�O�pF��|, ��A��A�s���ES0Z[tT0 k� �L��L	E1 4#Q&�1D"3Q  ��   � 3 3�@pG	S�Q�xF�#�|, ��A��A�w���C�0[[tT0 k� �|O��O	E1 4#Q&�1D"3Q  /�   � 3 3�@pG	S�S��F�+�|, ��A��A�{���C�0[[tT0 k� �xR�|R	E1 4#Q&�1D"3Q  ��    � 3 3�@pH	S�U��F�3�|, ��A��A�{���C�,\[tT0 k� �tU�xU	E1 4#Q&�1D"3Q  ��    � 3 3�@pI	c�V��F�;�|, �A��A����C�,][tT0 k� �pX�tX	E1 4#Q&�1D"3Q  ��    � 3 3�@lJ	c�Y��F�K�|, �A��A����C�$^[tT0 k� �h^�l^	E1 4#Q&�1D"3Q  ��    � 3 3�@lK	c�[ШF�S�|, �A��A����C�$^[tT0 k� �ha�la	E1 4#Q&�1D"3Q  ��    � 3 C�@hL	c�\аF[�|, �A��A����C� _[tT0 k� �de�he	E1 4#Q&�1D"3Q  ��    � 3 C�@hL	S�^иFc�|, �A��A����C�`[tT0 k� �`h�dh	E1 4#Q&�1D"3Q  ��    � 3 C�@hM	S�_��Fk�|, �A��A����C�`[tT0 k� �\k�`k	E1 4#Q&�1D"3Q  ��    � 3 C�	@dN	S�`��Fs�|, �A��A���#�C�a[tT0 k� �Xn�\n	E1 4#Q&�1D"3Q  ��    � 3 C�
@dN	S�a��F{�|, �A��A���#�C�a[tT0 k� �Tq�Xq	E1 4#Q&�1D"3Q  ��    � 3 C�
@`O	S�c��F��|, �A��A���#�C�bZ4T0 k� �Pt�Tt	E1 4#Q&�1D"3Q  ��    � 3 C�@`P	c�d��F��|, �A��A���#�C�bZ4T0 k� �Lw�Pw	E1 4#Q&�1D"3Q  ��    � 3 C�@`P	c�e��E��|, �A��A���#�C�cZ4 T0 k� �Hz�Lz	E1 4#Q&�1D"3Q  ��    � 3 C�L�\Q	c�f��E��|, #�A��A���'�C� dZ4 T0 k� �H}�L}	E1 4#Q&�1D"3Q  ��    � 3 C�L�\R	c�g��E��|, #�A��A���'�C��dZ4 T0 k� �D��H�	E1 4#Q&�1D"3Q  ��    � 3 C�L�XS	c�h� E�|, +�A��A���'�C��eZ4$T0 k� �<��@�	E1 4#Q&�1D"3Q  )�    � 3 S�L�XS	S�i�E�|, +�A��A���'�C��fZ4(T0 k� �8��<�	E1 4#Q&�1D"3Q  /�    � 3 S�L�TT	S�j�E�|, /�A��A���+�ER�fZ4(T0 k� �4��8�	E1 4#Q&�1D"3Q  ��    � 3 S�L�TU	S�k�E�|, /�A��A���+�ER�gZ4(T0 k� �0��4�	E1 4#Q&�1D"3Q  ��    � 3 S�L�TU	S�k�E�!�, 3�A��A���+�ER�gZ4,T0 k� �0��4�	E1 4#Q&�1D"3Q  ��    � 3 S�L�PV	S�l� E�!�, 3�A��A���+�ER�hZ4,T0 k� �,��0�	E1 4#Q&�1D"3Q  ��    � 3 S�L�PV	c�m�$E�!�, 7�A��A���+�ER�hZ40T0 k� �(��,�	E1 4#Q&�1D"3Q  ��    � 3 S�L�PW	c�m�,E�!�, 7�A��A���+�I��hZ40T0 k� �$��(�	E1 4#Q&�1D"3Q  ��    � 3 S�L�LW	c�n�0E�!�, ;�A��A����/�I��iZ40T0 k� � ��$�	E1 4#Q&�1D"3Q  ��    � 3 S�L�LX	c�n�8E�!�, ;�A��A����/�I��iZ44T0 k� �� 	E1 4#Q&�1D"3Q  ��    � 3 S�L�LX	c�n�<E� 	!�, ?�A��A����/�I��iZ44T0 k� ��	E1 4#Q&�1D"3Q  ��    � 3 S�!L�LY	S�o�DE�
!�, ?�A��A����/�I��jZ48T0 k� �~�~	E1 4#Q&�1D"3Q  ��    � 3 c�"L�HY	S�o�HE�!�, C�A��A����/�EҰjZ48 T0 k� �}�}	E1 4#Q&�1D"3Q  ��    � 3 c�$L�HZ	S�o�LE�!�, C�A��A����/�EҬjZ48 T0 k� �|�|	E1 4#Q&�1D"3Q  ��    � 3 c�&L�HZ	S�p�TE� !�, G�A��A����3�EҤjZ4< T0 k� �|�|	E1 4#Q&�1D"3Q  ��    � 3 c�(L�D[	S�p�XE�$|, G�A��A����3�EҠkZ4<!T0 k� �{�{	E1 4#Q&�1D"3Q  ��    � 3 c�)L�D[	c�p�\E�,|, K�A��A����3�EҜkZ4<!T0 k� �z�z	E1 4#Q&�1D"3Q  ��    � 3 ��+L�D\	c�p�dE�4|, K�A��A����3�E�kZ4@"T0 k� �y�y	E1 4#Q&�1D"3Q  ��    � 3 ��-L�D\	c�p�hE�<|, O�A��A����3�E�kZ4@"T0 k� � y�y	E1 4#Q&�1D"3Q  ��    � 3 ��.L�@]	c�p�lE�@|, O�A��A����3�E�lZ4@"T0 k� ��x� x	E1 4#Q&�1D"3Q  ��    � 3 ��0L�@]	c�p�tE�H|, O�A��A����7�E�lZ4@#T0 k� ��w��w	E1 4#Q&�1D"3Q  ��    � 3 ��2L�@^�p�xE�L|, S�A��A����7�E�|mZ4D#T0 k� ��w��w	E1 4#Q&�1D"3Q  ��    � 3 ��3L�@^�p�|E�T|, S�A��A����7�E�xmZ4D$T0 k� ��v��v	E1 4#Q&�1D"3Q  ��    � 3 ��5L�<^�p��E�\|, W�A��A����7�E�pnZ4D$T0 k� ��u��u	E1 4#Q&�1D"3Q  ��    � 3 ��7L�<_�p��E�`|, W�A��A����7�E�lnZ4H$T0 k� ��t��t	E1 4#Q&�1D"3Q  ��    � 3 ��8@<_�p��E�h|, W�A��A����7�E�doZ4H%T0 k� ��t��t	E1 4#Q&�1D"3Q  ��    � 3 ��:@<`S�p��E�l!�, [�A��A����7�E�`oZ4H%T0 k� ��s��s	E1 4#Q&�1D"3Q  ��    � 3 ��;@8`S�p��E�t!�, [�A��A����7�E�XpZ4L%T0 k� ��r��r	E1 4#Q&�1D"3Q  ��    � 3 ��=@8`S�p��E�x!�, _�A��A����;�E�TpZ4L&T0 k� ��r��r	E1 4#Q&�1D"3Q  ��    � 3 ��>@4aS�p��E!�, _�A��A����;�E�LqZ4L&T0 k� ��q��q	E1 4#Q&�1D"3Q  ��    � 3 ��@@4aS�p��E!�, _�A��A����;�E�DqZ4L&T0 k� ��p��p	E1 4#Q&�1D"3Q  ��    � 3 ��A@0a��p��E!�, c�A��A����;�E�@qZ4P'T0 k� ��o��o	E1 4#Q&�1D"3Q  ��    � 3 ��B@0b��p��E!�, c�A��A����;�E�8pZ4P'T0 k� ��o��o	E1 4#Q&�1D"3Q  ��    � 3 ��D@0b��p��E!�, c�A��A����;�E�4pZ4P'T0 k� ��n��n	E1 4#Q&�1D"3Q  ��    � 3 ��E@,b��p��E!�, g�A��A����;�E�0pZ4P(T0 k� ��m��m	E1 4#Q&�1D"3Q  ��    � 3 ��F@,b��p��E !�, g�A��A����;�E�(pZ4T(T0 k� ��m��m	E1 4#Q&�1D"3Q  ��    � 3 ��H@(c��p��E¤!�, g�A��A����?�E�$pZ4T(T0 k� ��l��l	E1 4#Q&�1D"3Q  ��    � 3 ��I@(c��p��E¨|, k�A��A����?�E�pZ4T)T0 k� ��k��k	E1 4#Q&�1D"3Q  ��    � 3 ��J@(c��p��E¬|, k�A��A����?�E�pZ4T)T0 k� ��j��j	E1 4#Q&�1D"3Q  ��    � 3 ��K@$c��o��E´|, k�A��A����?�FpZ4X)T0 k� �j��j	E1 4#Q&�1D"3Q  ��    � 3 ��M@$d��o��E¸|, o�AûA����?�FpZ4X*T0 k� �i��i	E1 4#Q&�1D"3Q  ��    � 3 ��N@$d��o��E¼|, o�AúA����?�FpZ4X*T0 k� �h��h	E1 4#Q&�1D"3Q  ��    � 3 ��O@ d��n��E��|, o�AúA���?�FpZ4X*T0 k� �h��h	E1 4#Q&�1D"3Q  ��    � 3 ��P@ dS�n��E��|, s�AúA���?�F qZ4X*T0 k� �g��g	E1 4#Q&�1D"3Q  ��    � 3 ��Q@ dS�n��E��|, s�AùA���?�F�qZ4\+T0 k� �f��f	E1 4#Q&�1D"3Q  ��    � 3 ��S@ dS�n��E��|, s�AùA���C�F�qZ4\+T0 k� �f��f	E1 4#Q&�1D"3Q  ��    � 3 ��T@ dS�n��E�� |, s�AøA���C�F�rZ4\+T0 k� �e��e	E1 4#Q&�1D"3Q  ��    � 3 ��U@ dS�n��E�� |, w�AøA���C�E��rZ4\,T0 k� �d��d	E1 4#Q&�1D"3Q  ��    � 3 ��V@ dS�n��E��!|, w�AøA���C�E��rZ4`,T0 k� �d��d	E1 4#Q&�1D"3Q  ��    � 3 ��W@ dS�m��E��!|, w�A÷A���C�E��sZ4`,T0 k� �c��c	E1 4#Q&�1D"3Q  ��    � 3 ��W@$dS�m��E��"|, {�A÷A���C�E��sZ4`,T0 k� �b��b	E1 4#Q&�1D"3Q  ��    � 3 ��X@$dS�m��E��"|, {�AöA���C�E��sZ4`-T0 k� �b��b	E1 4#Q&�1D"3Q  ��    � 3 ��X@$eS�m��E��#|, {�AöA���C�E��tZ4`-T0 k� �a��a	E1 4#Q&�1D"3Q  ��    � 3 ��Y@$eS�l��E��#|, {�AöA���C�E��tZ4d-T0 k� �`��`	E1 4#Q&�1D"3Q  ��    � 3 ��Z@$eS�l��E��#|, �AõA���C�E��tZ4d-T0 k� �`��`	E1 4#Q&�1D"3Q  ��    � 3 ��Z@(fS�l��E��$|, �AõA���C�E��uZ4d-T0 k� �_��_	E1 4#Q&�1D"3Q  ��   � 3 ��[@(fS�l��E��$|, �AõA���G�E��uZ4d.T0 k� �^��^	E1 4#Q&�1D"3Q  ��    � 3 ��[@(fc�l�E� %|, �AôA���G�E��uZ4d.T0 k� �^��^	E1 4#Q&�1D"3Q  ��    � 3 ��\@(fc�l�E�%|, ��AôA���G�E��vZ4d.T0 k� �]��]	E1 4#Q&�1D"3Q  ��    � 3 ��\@(gc�m�E�%|, ��AôA���G�E��vZ4h.T0 k� �|\��\	E1 4#Q&�1D"3Q  ��    � 3 ��]@(gc�m�E�&|, ��AóA���G�E��vZ4h/T0 k� �|\��\	E1 4#Q&�1D"3Q  ��    � 3 ��]@(gc�m�E�&|, ��AóA���G�E��wZ4h/T0 k� �x[�|[	E1 4#Q&�1D"3Q  ��    � 3 ��]@(gc�m�E�'|, ��AóA���G�@�wZ4h/T0 k� �tZ�xZ	E1 4#Q&�1D"3Q  ��    � 3 ��]@$gc�m� E�'|, ��AǲA���G�@�wZ4h/T0 k� �pZ�tZ	E1 4#Q&�1D"3Q  ��    � 3 ��^@$fc�n�$E�'|, ��AǲA���G�@�wZ4h/T0 k� �pY�tY	E1 4#Q&�1D"3Q  ��    � 3 ��^@$fc�n�(E�(|, ��AǲA���G�@�xZ4l0T0 k� �lX�pX	E1 4#Q&�1D"3Q  ��    � 3 ��^@$fc�n�0E�(|, ��AǲA���G�@�xZ4l0T0 k� �hX�lX	E1 4#Q&�1D"3Q  ��    � 3 ��^@ fc�n�4E� (|, ��AǱA���G�@�xZ4l0T0 k� �dW�hW	E1 4#Q&�1D"3Q  ��    � 3 ��^L� fc�n�<E�$)|, ��AǱA���G�@�xZ4l0T0 k� �dV�hV	E1 4#Q&�1D"3Q  ��    � 3 ��^L� fc�o�@E�()|, ��AǱA���K�@�yZ4l0T0 k� �`V�dV	E1 4#Q&�1D"3Q  ��    � 3 ��^L� fc�o�HE�()|, ��AǱA�#��K�@�yZ4l1T0 k� �\U�`U	E1 4#Q&�1D"3Q  ��    � 3 ��^L� fc�o�LE�,*|, ��AǰA�#��K�@�yZ4l1T0 k� �XT�\T	E1 4#Q&�1D"3Q  ��    � 3 ��^L� fc�o�TE�0*|, ��AǰA�#��K�@�yZ4p1T0 k� �XT�\T	E1 4#Q&�1D"3Q  ��    � 3 ��^L� fc�o�XE�4*|, ��AǰA�#��K�@�zZ4p1T0 k� �TS�XS	E1 4#Q&�1D"3Q  ��    � 3 ��^L�fc�o�`E�8+|, ��AǯA�'��K�@�zZ4p1T0 k� �PR�TR	E1 4#Q&�1D"3Q  ��    � 3 ��^L�fc�p�dE�<+|, ��AǯA�'��K�@�zZ4p1T0 k� �PN�TN	E1 4#Q&�1D"3Q  ��3    � 3 ��^L�fc�p�hE�<,|, ��AǯA�'��K�@�zZ4p2T0 k� �\K�`K	E1 4#Q&�1D"3Q  ��3    � 3 C�^L�fc�p�pE�@,|, ��AǯA�'��K�@�{Z4p2T0 k� �dI�hI	E1 4#Q&�1D"3Q  ��3    � 3 C�^L�fc�p�tE�D-|, ��AǯA�'��K�@�{Z4p2T0 k� �lH�pH	E1 4#Q&�1D"3Q  ��3    � 3 C�^L�gc�p�xE�H.|, ��AǮA�+��K�@�{Z4t2T0 k� �pG�tG	E1 4#Q&�1D"3Q  ��3    � 3 C�_L�gc�p��E�L.|, ��AǮA�+��K�@�{Z4t2T0 k� �tF�xF	E1 4#Q&�1D"3Q  ��3    � 3 C�_L�gc�q��E�P/|, ��AǮA�+��K�@�{Z4t2T0 k� �|E��E	E1 4#Q&�1D"3Q  ��3    � 3 C�`L�gc�q��E�T0|, ��AǮA�+��K�@�|Z4t3T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 C�`L�gc�q��E�X0|, ��AǭA�+��K�@�|Z4t3T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 C�aL�gc�q��E�\1|, ��AǭA�/��K�@�|Z4t3T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 C�aL�gc�q��E�`1|, ��AǭA�/��O�@�|Z4t3T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 C�aL�gc�q��E�d2|, ��AǭA�/��O�@�}Z4t3T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 C�aL�gc�q��E�h3|, ��A˭A�/��O�@�}Z4x3T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 3�aL�gc�r��E�p4|, ��A˭A�3��O�@�}Z4x4T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 3�aL�gc�s��E�p4|, ��AˬA�3��O�@�}Z4x4T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 3�aL�gc�s��E�t5|, ��AˬA�3��O�@�}Z4x4T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 3�aL�gc�t��E�x5|, ��AˬA�3��O�@�~Z4x4T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 3�aL�gc�t��E�|6|, ��AˬA�3��O�@�~Z4x4T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 #�aL�gc�t��E��6|, ��AˬA�3��O�@�~Z4x4T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 #�bL�gc�u��EÄ7|, ��AˬA�7��O�@�~Z4x4T0 k� �E��E	E1 4#Q&�1D"3Q  ��3    � 3 #�b@gc�u��EÄ7|, ��AϬA�7��O�@�~Z4x5T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 #�c@gc�v��EÈ8|, ��AϬA�7��O�@�Z4|5T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 #�d@gS�v��EÌ8|, ��AϫA�7��O�@�Z4|5T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 #�e@gS�v��EÐ9|, ��AϫA�7��O�@�Z4|5T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 �e@gS�w��EÐ9|, ��AϫA�7��O�@�Z4|5T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 �f@dhS�w��EÔ:|, ��AϫA�7��O�@�Z4|5T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 �g@dhS�x��EØ:|, ��AϫA�;��O�@�Z4|5T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 �g@dhS�x��EÜ;|, ��AϫA�;��O�@�Z4|5T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 �g@d h��x��EÜ;|, ��AϫA�;��O�@��Z4|5T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 �h@d h��x��Eà<|, ��AϫA�;��S�@�Z4|6T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 ��iE� h��y��Eä<|, ��AϫA�;��S�@�Z4|6T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 ��iE�$g��y��Eä<|, ��AӫA�;��S�@�Z4�6T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 ��jE�$g��y��Eè=|, ��AӪA�;��S�@�Z4�6T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 ��jE�$g��y��Eì=|, ��AӪA�?��S�@�~Z4�6T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 ��jE�(f��y� Eì>|, ��AӪA�?��S�@�~Z4�6T0 k� ��E��E	E1 4#Q&�1D"3Q  ��3    � 3 ��kE�(f��y�Eð>|, ��AӪA�?��S�@�~Z4�6T0 k� ��E� E	E1 4#Q&�1D"3Q  ��3    � 3 s�kE�(f�x�Eô>|, ��AӪA�?��S�@�~Z4�6T0 k� ��E� E	E1 4#Q&�1D"3Q  ��3   � 3 s�kE�(e�x�Eô?|, ��AӪA�?��S�@�}Z4�6T0 k� � E�E	E1 4#Q&�1D"3Q  ��3    � 3 s�kE�(e�x�Eø?|, ��AӪA�?��S�@�}Z4�7T0 k� �E�E	E1 4#Q&�1D"3Q  ��3    � 3 s�kE�(d�x�Eø@|, ��AӪA�?��S�@�}Z4�7T0 k� �E�E	E1 4#Q&�1D"3Q  ��3    � 3 s�kC�(c�w�Eü@|, ��AӪA�?��S�@�}Z4�7T0 k� �E�E	E1 4#Q&�1D"3Q  ��3    � 3 s�kC�(c�w�Eü@|, ��AӪA�C��S�@�}Z4�7T0 k� �E�E	E1 4#Q&�1D"3Q  ��3    � 3 s�kC�(b�v�E��A|, ��AӪA�C��S�@�|Z4�7T0 k� �E�E	E1 4#Q&�1D"3Q  ��3    � 3 ��kC�(a�v�E��A|, ��AӪA�C��S�@�|Z4�7T0 k� �E�E	E1 4#Q&�1D"3Q  ��3    � 3 ��kC�(`�u� E��A|, ��AשA�C��S�@�|Z4�7T0 k� �E�E	E1 4#Q&�1D"3Q  ��3    � 3 ��jC�(`�u� E��B|, ��AשA�C��S�@�|Z4�7T0 k� �E�E	E1 4#Q&�1D"3Q  ��3    � 3 ��jC�(_�t�$E��B|, ��AשA�C��S�@�|Z4�7T0 k� �E� E	E1 4#Q&�1D"3Q  ��3    � 3 ��iC�(_�t�(E��B|, ��AשA�C��S�@�{Z4�7T0 k� � E�$E	E1 4#Q&�1D"3Q  ��3    � 3 ��iC�(^�s�(E��C|, ��AשA�C��S�@�{Z4�7T0 k� �$E�(E	E1 4#Q&�1D"3Q  ��3    � 3 ��iC�(^Ӵr�,E��C|, ��AשA�C��S�@�{Z4�8T0 k� �$E�(E	E1 4#Q&�1D"3Q  ��3    � 3 ��hC�(]Ӵr�0E��C|, ��AשA�G��S�@�{Z4�8T0 k� �(E�,E	E1 4#Q&�1D"3Q  ��3    � 3 ��hC�(]Ӵq�0E��D|, ��AשA�G��S�@�{Z4�8T0 k� �,E�0E	E1 4#Q&�1D"3Q  ��3    � 3 ��hC�(\Ӵp�4E��D|, ��AשA�G��S�@�{Z4�8T0 k� �,E�0E	E1 4#Q&�1D"3Q  ��3    � 3 ��hC�(\Ӹo�8E��D|, ��AשA�G��S�@�zZ4�8T0 k� �0E�4E	E1 4#Q&�1D"3Q  ��3    � 3 ��hC�(\Ӹn�8E��E|, ��AשA�G��S�@�zZ4�8T0 k� �0E�4E	E1 4#Q&�1D"3Q  ��3    � 3 ��hC�([Ӹn�<E��E|, ��AשA�G��W�@�zZ4�8T0 k� �4E�8E	E1 4#Q&�1D"3Q  ��3    � 3 ��gC�([Ӹm�<E��E|, ��AשA�G��W�@�zZ4�8T0 k� �8E�<E	E1 4#Q&�1D"3Q  ��3    � 3 ��gC�([Ӹl @E��E|, ��AשA�G��W�@�zZ4�8T0 k� �LD�PD	E1 4#Q&�1D"3Q  ��3    � 3 ��xE}3���>��<���'��G�A��6E����EˣZ3�T0 k� �;��?�	E1 4#Q&�1D"3Q  ��    �������wE}7���>��<���'��?�A��4E����EˣZ3�T0 k� �?��C�	E1 4#Q&�1D"3Q  ��    ������vE}7���=��<���'��;�A��3E����EϤZ3�T0 k� �C��G�	E1 4#Q&�1D"3Q  ��    ������uE};���=��<���'��3�E��2E����EϤZ3�T0 k� �G��K�	E1 4#Q&�1D"3Q  ��    ������tE}?���=���l���'��/�E��1E����EӤZ3�T0 k� �K��O�	E1 4#Q&�1D"3Q  ��    ������sEmC���=�� l���'��'�E��0E����EӤZ3�T0 k� �?��C�	E1 4#Q&�1D"3Q  ��    ������qEmC���=�� l���'��#�E��/E����EפZ3�T0 k� �3��7�	E1 4#Q&�1D"3Q  ��    �������pEmG���=��l���'���E��/E�����E�ۤZ3�T0 k� �/��3�	E1 4#Q&�1D"3Q  ��    �������oEmK���=��l���'���E��.E�����E�ۤZ3�T0 k� �+��/�	E1 4#Q&�1D"3Q  ��    �������mEmO���=��l���'���E��-E����E�ߤZ3�T0 k� �+��/�	E1 4#Q&�1D"3Q  ��    �������kEmO���=��l���'�	}�E��,E���E��Z3�T0 k� �'��+�	E1 4#Q&�1D"3Q  ��    �������jEmO���=��l��|'�	|��E��,E��w�E��Z3�T0 k� �#��'�	E1 4#Q&�1D"3Q  ��    �������iEmS���=��l��|+�	|��E}�+E��s�E��Z3�T0 k� �'��+�	E1 4#Q&�1D"3Q  ��    �������gEmS���=��l��|+�	|��E}�+E��o�E��Z3�T0 k� �'��+�	E1 4#Q&�1D"3Q  ��    �������fEmS���=��l��|+�	|��E}�+E��k�E��Z3�T0 k� �'��+�	E1 4#Q&�1D"3Q  ��    �������eI�S���=��
��|+�	|��E}�+E��g�D��Z3�T0 k� �+��/�	E1 4#Q&�1D"3Q  ��    ������cI�W���=��
��|+�	���E}�*E��_�D���Z3�T0 k� �/��3�	E1 4#Q&�1D"3Q  ��    ������bI�W���=��
��|+�	���BM�*E��[�D���Z3�T0 k� �3��7�	E1 4#Q&�1D"3Q  ��    ������`I�W���=��	
��|+�	���BM�*E��W�D���Z3�T0 k� �3��7�	E1 4#Q&�1D"3Q  ��    ������_I�W���=��

��|+�	���BM�*E��O�D��Z3�T0 k� �3��7�	E1 4#Q&�1D"3Q  ��    ������]E�W���=��

��|/�	���BM�*E��K�D��Z3�T0 k� �3��7�	E1 4#Q&�1D"3Q  ��    ������\E�S���=��
��|/�L��BM�*E��G�D��Z3�T0 k� �3��7�	E1 4#Q&�1D"3Q  ��    ������YE�S���=��
��|/�L��@m�*E��;�D��Z3�T0 k� �3��7�	E1 4#Q&�1D"3Q  ��    ������WE�S���=��
��|/�L��@m�*E��3�D��Z3�T0 k� �3��7�	E1 4#Q&�1D"3Q  ��    ������UE�S���=��
��|/�L��@m�*E��+�D��Z3�T0 k� �/��3�	E1 4#Q&�1D"3Q  ��    �������TE�O���=��
��|/�L��@m�*E��'�D��Z3�T0 k� �,�0	E1 4#Q&�1D"3Q  ��    �������RE�O���=��
L��|/�L��@m�)E���D�#�Z3�T0 k� �,�0	E1 4#Q&�1D"3Q  ��    �������QE�O���=��
L��|/�L��B��)E���D�+�Z3�T0 k� �4�8	E1 4#Q&�1D"3Q  ��    �������OE�K���=��
L��|/�L��B��)E���D�/�Z3�T0 k� �<�@	E1 4#Q&�1D"3Q  ��    �������ME�K���=��
L��|/�	|��B��)E���D�3�Z3�T0 k� �D	�H		E1 4#Q&�1D"3Q  ��    �������ME�G���=��
L��|/�	|��B��(E���D�7�Z3�T0 k� �D�H	E1 4#Q&�1D"3Q  ��    �������ME�G���<��
L��|/�	|��B��(E�����F?�Z3�T0 k� �H�L	E1 4#Q&�1D"3Q  ��    �������KE�C���;��
L��|/�	|��E��'E�����FG�Z3�T0 k� �H�L	E1 4#Q&�1D"3Q  ��    �������KE�@ ��;��
L��|/�	|��E��'E�����FO�Z3�T0 k� �L�P	E1 4#Q&�1D"3Q  ��    �������JE�@��;��
L��|/�	���E��&E�����FS�Z3�T0 k� �L�P	E1 4#Q&�1D"3Q  ��    �������IE�<��:��
L��|/�	�� E��&D��A��E�[�Z3�T0 k� �H�L	E1 4#Q&�1D"3Q  ��    �������HE�<��:��
L��|/�	�� E��%D��A��E�_�Z3�T0 k� �H�L	E1 4#Q&�1D"3Q  ��    �������GF<	��:�� ���|, 	��E��$D��A��E�g�Z3�T0 k� �P�T	E1 4#Q&�1D"3Q  ��    �������GF<��:��"���|,	��E��$D���A��E�k�Z3�T0 k� �T�X	E1 4#Q&�1D"3Q  ��    �������FF8��:��#���|,	|�E��#D���A��E�s�Z3�T0 k� �X�\	E1 4#Q&�1D"3Q  ��    ������EF8��9��&���|,	|�E��!D���A��B��Z3�T0 k� �\!�`!	E1 4#Q&�1D"3Q  ��    ������EF8��9��(���|,	|�E��!D���A��B���Z3�T0 k� �`"�d"	E1 4#Q&�1D"3Q  ��    ������DF8��9��)���|,	|�E�� D���A��B���Z3�T0 k� �d$�h$	E1 4#Q&�1D"3Q  ��    ������DF8��9��+���|,	��E��D���A��B���Z3�T0 k� �d'�h'	E1 4#Q&�1D"3Q  ��    ������CF8��9��,���|,	��E��D���A��B���Z3�T0 k� �d)�h)	E1 4#Q&�1D"3Q  ��    ������ CF8��9��.���|,	��E��D���1�B���Z3�T0 k� �d+�h+	E1 4#Q&�1D"3Q  ��    ������(CF8 ��9��/���|,	��E��D��1w�B���Z3�T0 k� �d.�h.	E1 4#Q&�1D"3Q  ��    ������,CF8"��9��0���|,	��E��D��1o�B���Z3�T0 k� �d0�h0	E1 4#Q&�1D"3Q  ��    ������4CE�<$��9��2���|,�|E��D��1g�B���Z3�T0 k� �d.�h.	E1 4#Q&�1D"3Q  ��    ������8CE�<'��9��3���|,�|E��D��1_�B���Z3�T0 k� �`.�d.	E1 4#Q&�1D"3Q  ��    ������DCE�@+��9	��5���|,	�xE��D��1S�B���Z3�T0 k� �`0�d0	E1 4#Q&�1D"3Q  ��    ������LCE�@-^�9	��6���|,	�xE��D��1K�B���Z3�T0 k� �\0�`0	E1 4#Q&�1D"3Q  ��    ������PCE�D0^�9	��8���|,	�tE��D��1C�B���Z3�T0 k� �`1�d1	E1 4#Q&�1D"3Q  ��    ������TCE�D2^�9	��9���|,	�pA��D��1;�B���Z3�T0 k� �`3�d3	E1 4#Q&�1D"3Q  ��    ������\D@-H4^�9	��:����,	�pA��D��17�B���Z3�T0 k� �t5�x5	E1 4#Q&�1D"3Q  ��    ������`D@-L6^�9	��:����,	�lA��D��1/�B���Z3�T0 k� ��7��7	E1 4#Q&�1D"3Q  ��    ������dE@-P8^�9	��;����,
�lA��D��!'�B���Z3�T0 k� ��9��9	E1 4#Q&�1D"3Q  ��    ������lE@-P:^�9	��<L���(
�l	A��D��!#�B��Z3�T0 k� ��;��;	E1 4#Q&�1D"3Q  ��    ������tF@-X>^�9	��>L���$
�h
E��D��!�B��Z3�T0 k� ��?��?	E1 4#Q&�1D"3Q  ��    ������xG@-\@^�9��?L���$�hE��D��!�B��Z3�T0 k� ��A��A	E1 4#Q&�1D"3Q  ��    ������|H@-`B^�9��?L���$�hE��D��!�B��Z3�T0 k� ��C��C	E1 4#Q&�1D"3Q  ��    �����πH@-dC^�9��@,���$�dE��D��!�B�'�Z3�T0 k� ��D��D	E1 4#Q&�1D"3Q  ��    �����τI@-hE^�9��A,���$�dE��D�߫ ��B�/�Z3�T0 k� ��F��F	E1 4#Q&�1D"3Q  ��    �����ψJE�pG^�9��B,���$�dEm�D�߬ ��B�7�Z3�T0 k� ��F��F	E1 4#Q&�1D"3Q  ��    �����όKE�tI^�9�C,���$�dEm�D�߮ ��B�?�Z3�T0 k� ��H��H	E1 4#Q&�1D"3Q  ��    �  ��ϐLE��L^�9�D,���$�`Em�D�߰ ��B�O�Z3�T0 k� ��K��K	E1 4#Q&�1D"3Q  ��    � ��ϔME��N^�9�E,���$�`Em�D�۲ ��B�W�Z3�T0 k� ��M��M	E1 4#Q&�1D"3Q  ��    � ��ϘNE��P^�9�F,���$�`E��D�۳��B�[�Z3�T0 k� ��N��N	E1 4#Q&�1D"3Q  ��    � ��ߘOE��R^�9�G����$�`E��D�۵��B�c�Z3�T0 k� ��P��P	E1 4#Q&�1D"3Q  ��    � ��ߜPE��S^�9�G����$�`E��D�۶��B�k�Z3�T0 k� ��R��R	E1 4#Q&�1D"3Q  ��    � 
��ߜQE��U^�9�H����$�`E��D�׸��B�s�Z3�T0 k� ��S��S	E1 4#Q&�1D"3Q  ��    � ��ߠRE��V^�9�I����$�`E��D�׺��B�{�Z3�T0 k� ��U��U	E1 4#Q&�1D"3Q  ��    � ��ߠRE��X^�9�I����$�`F�D�׻���B߃�Z3�T0 k� ��W��W	E1 4#Q&�1D"3Q  ��    � ���SE��Z^�9��J����$�`F�D�׽���Bߋ�Z3�T0 k� ��T��T	E1 4#Q&�1D"3Q  ��    � ���TE��[^�9��J����$�`F�D�׿���Bߓ�Z3�T0 k� ��S��S	E1 4#Q&�1D"3Q  ��    � ���UE��^^�9��K����$�`F�!D������Bߣ�Z3�T0 k� ��S��S	E1 4#Q&�1D"3Q  �� 	   � ���UE��_^�9��K����$�`F�"D������Bߧ�Z3�T0 k� ��S��S	E1 4#Q&�1D"3Q  �� 	   � ����VE��`^�9��K����$�`F�#D������B߯�Z3�T0 k� ��S��S	E1 4#Q&�1D"3Q  �� 	   � ����VE��a^�9��KL���$�`F�$Eb�����B߷�Z3�T0 k� ��S��S	E1 4#Q&�1D"3Q  �� 	   � ����WE��b^�9��KL���$�`F�%Eb�����B߿�Z3�T0 k� ��S� S	E1 4#Q&�1D"3Q  �� 	   � ����WE��c^�9��KL���$�`E��&Eb�����B���Z3�T0 k� �T�T	E1 4#Q&�1D"3Q  �� 	   � ����W@}�d^�9��KL���$�`E��'Eb�����B���Z3�T0 k� �S�S	E1 4#Q&�1D"3Q  �� 	   � ��O�W@}�e^�9��KL���$�`E��(Eb�����B���Z3�T0 k� �R�R	E1 4#Q&�1D"3Q  �� 	   � ��O�W@~ f^�9��K	\���$�`E��)Eb�����B���Z3�T0 k� �R� R	E1 4#Q&�1D"3Q  �� 	   �  ��O�W@~g^�9��K	\���$�`E��*Eb�����B���Z3�T0 k� �$Q�(Q	E1 4#Q&�1D"3Q  �� 	   � !��O�W@~g^�9��K	\���$�`B��+Eb�����B���Z3�T0 k� �,Q�0Q	E1 4#Q&�1D"3Q  �� 	   � "��O�WEh^�9��K	\���$�`B��+D2�����B���Z3�T0 k� �0Y�4Y	E1 4#Q&�1D"3Q  �� 	   � #���WE i^�9��K	\���$�`B��,D2�����B���Z3�T0 k� �4_�8_	E1 4#Q&�1D"3Q  �� 	   � $���WE(i��9��K	l���$�`B��-D2�����B��Z3�T0 k� �<c�@c	E1 4#Q&�1D"3Q  �� 	   � %���VE0j��9��K	l���$�`B��.D2���� B��Z3�T0 k� �Dg�Hg	E1 4#Q&�1D"3Q  �� 	   � &���VE<k��9��K	l���$�`B��/D2����J@�Z3�T0 k� �Lj�Pj	E1 4#Q&�1D"3Q  �� 	   � '���VE�Dk��9��K	l���$�`B��0D2����J@�Z3�T0 k� �\f�`f	E1 4#Q&�1D"3Q  �� 	   � (����VE�Ll��9L�K	l���$�dB��1D2����J@#�Z3�T0 k� �dd�hd	E1 4#Q&�1D"3Q  �� 	   � )����VE�Tm��9L�K	\���$�dB��1D2����J@+�Z3�T0 k� �lb�pb	E1 4#Q&�1D"3Q  �� 	   � *����VE�\m��9L�K	\���$�dB��2D2����J@/�Z3�T0 k� �ta�xa	E1 4#Q&�1D"3Q  �� 	   � +����VE�hm��9L�K	\���$�dB��3D2����E 7�Z3�T0 k� ��`��`	E1 4#Q&�1D"3Q  �� 	   � ,����UE�pn��9L�K	\���$�dB��4D2����E ;�Z3�T0 k� ��`��`	E1 4#Q&�1D"3Q  �� 	   � -����UExn��9L�K	\���$�hB��5D2����E C�Z3�T0 k� ��e��e	E1 4#Q&�1D"3Q  �� 	   � .����UE�n��9L�K	l���$�hB� 5DB����	E G�Z3�T0 k� ��h��h	E1 4#Q&�1D"3Q  �� 	   � /����UE�oN�9L�K	l���$�hB�6DB����
E K�Z3�T0 k� ��l��l	E1 4#Q&�1D"3Q  �� 	   � 0����UE�oN�9L�K	l���$�lB�7DB����E S�Z3�T0 k� ��n��n	E1 4#Q&�1D"3Q  �� 
   � 1����UE�oN�9L�K	l���$�lB�7DB����E0W�Z3�T0 k� ��o��o	E1 4#Q&�1D"3Q  �� 
   � 2����UE�pN�9 �K	l���$�pB�$8DB����E0[�Z3�T0 k� ��q��q	E1 4#Q&�1D"3Q  �� 
   � 3����UE�pN�9 �K	\���$�pB�,9DB����E0_�Z3�T0 k� ��r��r	E1 4#Q&�1D"3Q  �� 
   � 4����UE��pN�9 �K	\���$�tB�4:DB����E0g�Z3�T0 k� ��m��m	E1 4#Q&�1D"3Q  �� 
   � 5����TE��pN�9 �K	\���$�tB�<:DB|  �E0k�Z3�T0 k� ��j��j	E1 4#Q&�1D"3Q  �� 
   � 6����TE��qN�9 �K	\���$�xB�D;DBx! E0o�Z3�T0 k� ��h��h	E1 4#Q&�1D"3Q  �� 
   � 7��� TE��qN�9 �K	\���$�xB�L<DBt!E0s�Z3�T0 k� ��f��f	E1 4#Q&�1D"3Q  �� 
   � 8���TE��qN�9 �K	l���$�|
B�T<DBp!E0w�Z3�T0 k� ��e��e	E1 4#Q&�1D"3Q  �� 
   � 9���TE��qN�9 �K	l���$�	B�\=DRl	!E0{�Z3�T0 k� � d�d	E1 4#Q&�1D"3Q  �� 
   � :���TE��qN�9 �K	l���$�	B�d=DRh!E0�Z3�T0 k� �c�c	E1 4#Q&�1D"3Q  �� 
   � ;���TE��q �9 �K	l���$�B�l>DR`!E0��Z3�T0 k� �b�b	E1 4#Q&�1D"3Q  �� 
   � < �TE�q �9 �K	l���$�B�t?DR\!E@��Z3�T0 k� �b� b	E1 4#Q&�1D"3Q  �� 
   � < �$TE�q �9 �K ����$�B�|?DRX�E@��Z3�T0 k� �(b�,b	E1 4#Q&�1D"3Q  �� 
   � < �,T@q �9 �K ����$��B��@EbT�E@��Z3�T0 k� �0`�4`	E1 4#Q&�1D"3Q  �� 
   � < �0T@ q �9 �K ����$��B��@EbP� E@��Z3�T0 k� �<^�@^	E1 4#Q&�1D"3Q  �� 
   � < 
�8S@(p��9 �K ����$��O��AEbL�$!E@��Z3�T0 k� �H\�L\	E1 4#Q&�1D"3Q  �� 
   � < �@S@0p��9 �K ����$��O��BEbD�("E@��Z3�T0 k� �P[�T[	E1 4#Q&�1D"3Q  �� 
   � < �HS@<p��9 �K l��|$��O��CEb@1,#E@��Z3�T0 k� �XZ�\Z	E1 4#Q&�1D"3Q  �� 
   � < �PS@Dp��9 �K l��|$��O��DEb<10$E@��Z3�T0 k� �dY�hY	E1 4#Q&�1D"3Q  �� 
   � < �XS@Lo��8 �K l��|$�� O��DEb8 14%E@��Z3�T0 k� �lX�pX	E1 4#Q&�1D"3Q  �� 
   � < �\S@Xo��8 �K l��|$���O��EER0"18&E@��Z3�T0 k� �tX�xX	E1 4#Q&�1D"3Q  ��    � < �dS@`o��8 �K l��|$���O��FER,$1<'EP��Z3�T0 k� ��X��X	E1 4#Q&�1D"3Q  ��    � < �lS@hn��8 �K l��|$���O��FER(&1@(EP��Z3�T0 k� ��W��W	E1 4#Q&�1D"3Q  ��    � < �xS@tn��8 �K l��|$���O��GER (1D(EP��Z3�T0 k� ��W��W	E1 4#Q&�1D"3Q  ��    � < ��S@|n��7 �K l��|$��O��HER*1D)EP��Z3�T0 k� ��V��V	E1 4#Q&�1D"3Q  ��    � < ��SE�m��7 �K l��|$��O��HER,AH*EP� Z3�T0 k� ��]��]	E1 4#Q&�1D"3Q  ��    � < !��SE�m��7 �K l��|$��O��IER-AL*EP�Z3�T0 k� ��b��b	E1 4#Q&�1D"3Q  ��    � < $��SE�l��7 �K l��|$��O��JER/AP+EP�Z3�T0 k� ��e��e	E1 4#Q&�1D"3Q  ��    � < &��SE�l��7 �K l��|$��O��JER1AT+EP�Z3�T0 k� ��h��h	E1 4#Q&�1D"3Q  ��    � < )��SE�l� 6 �K l��|$��O��KEQ�3AX,EP�Z3�T0 k� ��i��i	E1 4#Q&�1D"3Q  ��    � < +��TE�k�6 �K m�|$��O��LEQ�4A\,J��Z3�T0 k� ��k��k	E1 4#Q&�1D"3Q  ��    � < .��TE�k�6 �K m�|$��O��LEA�6A`-J��Z3�T0 k� ��l��l	E1 4#Q&�1D"3Q  ��    � < 0��TE�j�6 �K m�|$��O��MEA�8Ad-J��	Z3�T0 k� ��l��l	E1 4#Q&�1D"3Q  ��    � < 2��TE�j�6 �K m�|$��O��MEA�9Qh-J��
Z3�T0 k� ��m��m	E1 4#Q&�1D"3Q  ��    � < 4��UE�j�5 �K m�|$��O��NEA�;Ql.J�Z3�T0 k� ��m��m	E1 4#Q&�1D"3Q  ��    � < 7��U@/�i� 5 �K m�|$��O��OEA�<Qp.J�Z3�T0 k� �l�l	E1 4#Q&�1D"3Q  ��    � < 9��U@/�i�(5 �K m�!�$��O��OEA�=Qt.J�b��T0 k� �k� k	E1 4#Q&�1D"3Q  ��    � < ;��V@/�i�,4 �K m�!�$��O��PEA�?Qx/J�b��T0 k� �0j�4j	E1 4#Q&�1D"3Q  ��    � < =��W@ h�83 �K m�!�$��O��QEA�A
ф/J�$b��T0 k� �Hi�Li	E1 4#Q&�1D"3Q  ��    � < @�WE�g�@3 �K m�!�$���O��QEA�B
ш/J�,b��T0 k� �Hd�Ld	E1 4#Q&�1D"3Q  ��    � < C�XE�g�D2 �K m�!�$
���B��REA�C
ь0J�4b��T0 k� �Ha�La	E1 4#Q&�1D"3Q  ��    � < F�YE� f�L1 �K m�!�$
���B��REA�D
є0J�8b��T0 k� �L]�P]	E1 4#Q&�1D"3Q  ��    � < H�ZE�(f�P1 �K m�!�$
���B��SE1�E
ј0J�@b��T0 k� �TZ�XZ	E1 4#Q&�1D"3Q  ��    � < J�$ZE�0e�X0 �K m�!�$	���B� SE1�F
Ѡ1J�Hb��T0 k� �XY�\Y	E1 4#Q&�1D"3Q  ��    � < L�,[E�<e�`0 �K m�!�$	���B�TE1�G
Ѥ1J�Lb��T0 k� �`W�dW	E1 4#Q&�1D"3Q  ��    � < N�4\@pDd�d/ �K m#�!�$���E�TE1�G
�1J�Tb��T0 k� �hT�lT	E1 4#Q&�1D"3Q  ��    � < P�D^@pTc�p- �K m#�|$���E�UE1tI
�2J�dZ3�T0 k� �|Q��Q	E1 4#Q&�1D"3Q  ��    � < S�L_@p`b�x, �K m'�|$��E�VE1pI
�2J�hZ3�T0 k� ��N��N	E1 4#Q&�1D"3Q  ��    � < V�P`@phb߀, �K m'�|$��E�VE1hI
��2J�pZ3�T0 k� ��L��L	E1 4#Q&�1D"3Q  ��    � < Y�Xa@ppa߈+ �K m+�|$��I WE1`J��2J�xZ3�T0 k� �K��K	E1 4#Q&�1D"3Q  ��    � < [�`c@px`ߌ* �K m+�|$��I$WE1\J��3J�Z3�T0 k� �I��I	E1 4#Q&�1D"3Q  ��    � < ]�ddE�`�) �K m+�|$��I(WE1TJ��3JфZ3�T0 k� �O��O	E1 4#Q&�1D"3Q  ��    � < `�leE�_�( �K m/�|$�#�I0XE�LJ��3JьZ3�T0 k� �T��T	E1 4#Q&�1D"3Q  ��    � < b�pfE�^�' �K m/�|$�'�I4XE�HJ��3Jє Z3�T0 k� �W��W	E1 4#Q&�1D"3Q  ��    � < d�xhE�^�& �K m/�|(�/�E8YE�@J��3Jќ!Z3�T0 k� �Y��Y	E1 4#Q&�1D"3Q  ��    � < f�|iE�]�% �K m3�|(�7�E@YE�<J��3JѠ!Z3�T0 k� �Z��Z	E1 4#Q&�1D"3Q  ��    � < h��lE�\��# �K m7�!�(�C�ELZE�0J��3JѰ#bs�T0 k� ��[��[	E1 4#Q&�1D"3Q  ��    � < k��mE�[��# �K m7�!�(�K�EPZE�(J� 4JѸ$bs�T0 k� ��\��\	E1 4#Q&�1D"3Q  ��    � < n��nE�Z��" �K m7�!�(�S�EXZE�$J�4J��%bs�T0 k� ��\��\	E1 4#Q&�1D"3Q  ��    � < qєpE�Z��! �K m;�!�(�W�B�`[E� I�4J��%bs�T0 k� ��\��\	E1 4#Q&�1D"3Q  ��    � < tєqE��Y��  �K m;�!�,�_�B�d[E�I�4J��&bs�T0 k� ��[��[	E1 4#Q&�1D"3Q  ��    � < wјsE��Y�� �K m;�!�,�g�B�l[E�H�4J��'bs�T0 k� ��Y��Y	E1 4#Q&�1D"3Q  ��    � < yќtE��X�� �K m?�!�,�o�B�t\E�H�4J��(bs�T0 k� � W�W	E1 4#Q&�1D"3Q  ��    � < {ѠuE��X�� �K m?�!�,�w�B�|\E�G�4J��(bs�T0 k� �W�W	E1 4#Q&�1D"3Q  �    � < }ѠwE��X�  �K m?�!�,��B��\E�F�4J��(bs�T0 k� �W�W	E1 4#Q&�1D"3Q  ��    � < ѤxE��X� �K mC�!�,���B��\E� E�5J��(bs�T0 k� �S�S	E1 4#Q&�1D"3Q  ��    � < �ѨzE�X� �K mC�|,���B��]C��A�$5J��)Z3�T0 k� �(P�,P	E1 4#Q&�1D"3Q  ��    � < �Ѩ|E�X�  �K mC�|,���B��]C��?�(6J��)Z3�T0 k� �0M�4M	E1 4#Q&�1D"3Q  ��    � < �Ѩ}E�X�( �K mG�|,���B��^C��=�,6J��)Z3�T0 k� �8L�<L	E1 4#Q&�1D"3Q  ��    � < �Ѭ~@q$W�0 �K mG�|,ͯ�B��^C��;�06J�)Z3�T0 k� �@I�DI	E1 4#Q&�1D"3Q  ��    � < �Ѭ@q,W�8 �K mG�|,ͷ�B��^C��9�46J�)Z3�T0 k� �HF�LF	E1 4#Q&�1D"3Q  ��    � < �ᬀ@q4W�@ �K mK�|,Ϳ�B��^C��7�46J�)Z3�T0 k� �PC�TC	E1 4#Q&�1D"3Q  ��    � < �ᬀ@q<V�H �K mK�|,���B��_C��5�86J�)Z3�T0 k� �XB�\B	E1 4#Q&�1D"3Q  ��    � < �ᬀ@qDV�P �K mK�|,���B��_C��3�<6J�)Z3�T0 k� �`@�d@	E1 4#Q&�1D"3Q  ��    � < ��@qLV�X �K mK�|,���B��_C��2�@6J�)Z3�T0 k� �l?�p?	E1 4#Q&�1D"3Q  ��    � < ��@qTU�` �K mO�|,���B��`C��0�D7J� )Z3�T0 k� �t>�x>	E1 4#Q&�1D"3Q  ��    � < ��@q\T�d �K mO�|,���B��`C��.H7J�$)Z3�T0 k� �|=��=	E1 4#Q&�1D"3Q  ��    � < �1�~@qhT�l��K O�|,���B��`C��,L6J�$)Z3�T0 k� �<��<	E1 4#Q&�1D"3Q  ��    � < �1�~@qpS	�t��K S�|,���B��`C��+P7J�,)Z3�T0 k� �<��<	E1 4#Q&�1D"3Q  ��    � < �1�}@qxS	�x��K S�|,���B�aC��)X7J�0)Z3�T0 k� �;��;	E1 4#Q&�1D"3Q  ��    � < �1�}@q�R	����K W�|,��B�aC��'\6J�8(Z3�T0 k� �:��:	E1 4#Q&�1D"3Q  ��    � < �1�|@��Q	����K W�|,��B�aC�x&�`6J�<(Z3�T0 k� �;��;	E1 4#Q&�1D"3Q  ��    � < �1�{@��P	����K�[�|,��B� aC�t$�d6J�D(Z3�T0 k� �:��:	E1 4#Q&�1D"3Q  ��    � < �1�z@��O
 ���K�_�|,�'�B�0bC�d!�l6J�D(Z3�T0 k� ��9��9	E1 4#Q&�1D"3Q  ��    � < ��y@��N
 ���K�c�|,�/�B�8bC�`�t6J�L'Z3�T0 k� ��9��9	E1 4#Q&�1D"3Q  ��    � < ��x@��M
 ���K�c�|,�7�B�@bC�Xrx6J�T'Z3�T0 k� ��8��8	E1 4#Q&�1D"3Q  ��    � < ��x@��M
 ���K�g�|,�C�B�LbC�Pr|5J�X'Z3�T0 k� ��7��7	E1 4#Q&�1D"3Q  ��    � < ��w@��L
 ���K�k�|,�K�B�TcC�Lr�5J�`&Z3�T0 k� ��6��6	E1 4#Q&�1D"3Q  ��    � < ��v@��K����K�o�|,�S�B�\cC�Dr�5E�h&Z3�T0 k� ��5��5	E1 4#Q&�1D"3Q  ��    � < ��u@��J����K�s�|,�[�B�dcC�@r�5E�l&Z3�T0 k� ��4��4	E1 4#Q&�1D"3Q  ��    � < ��s@��H��
��K�{�|,�k�B�tcC�4r�4E�x%Z3�T0 k� �3�3	E1 4#Q&�1D"3Q  ��    � < ��r@��H��
��K��|,�s�B�|dE@,r�3E�x%Z3�T0 k� �2�2	E1 4#Q&�1D"3Q  ��    � < ��q@��G��
��K���|,�{�BЄdE@$r�3E�|%Z3�T0 k� �1� 1	E1 4#Q&�1D"3Q  ��    � < ��p@�F��	��K���|,���BАdE@ r�2EҀ$Z3�T0 k� �$0�(0	E1 4#Q&�1D"3Q  ��    � < ��n@�E��	��K���|,���BИdE@��2E҄$Z3�T0 k� �,/�0/	E1 4#Q&�1D"3Q  ��    � < ��|m@�D��	��K���|,���BРdE@��1E҈#Z3�T0 k� �4.�8.	E1 4#Q&�1D"3Q  ��    � < ��|l@�C��	��K���|,���E��eE0��0C�#Z3�T0 k� �@-�D-	E1 4#Q&�1D"3Q  ��    � < ��xj@�$B����K���|,���E��eE0
��0C�#Z3�T0 k� �H,�L,	E1 4#Q&�1D"3Q  ��    � < ��xi@�0A����K���|,���E��eE0��/C�"Z3�T0 k� �P+�T+	E1 4#Q&�1D"3Q  ��    � < ��th@�8@����Kͣ�|,���E��eE?��.C�"Z3�T0 k� �X*�\*	E1 4#Q&�1D"3Q  ��    � < ��pe@�H>���Kͯ�|,�ǷE��eE?��-C�!Z3�T0 k� �h(�l(	E1 4#Q&�1D"3Q  ��    � < �lc@�P=���Kͳ�|,�ϷE��fE?��,C�!Z3�T0 k� �l)�p)	E1 4#Q&�1D"3Q  ��    � < �la@�X<���Kͻ�|,�׶E��fE?���+C� Z3�T0 k� �p)�t)	E1 4#Q&�1D"3Q  ��    � < �h`@�`;� ��KͿ�|,�߶E��fE/���*C� Z3�T0 k� �x)�|)	E1 4#Q&�1D"3Q  ��    � < �h^@�h:�(�K���|,��E��fE/���*C� Z3�T0 k� �|)��)	E1 4#Q&�1D"3Q  ��    � < �h]@�p9�0�K���|,��E��fE/����)EҠZ3�T0 k� �(��(	E1 4#Q&�1D"3Q  ��    � < �h[@�x8�8�K���|,���B�fE/����(EҠZ3�T0 k� �'��'	E1 4#Q&�1D"3Q  ��    � < �dY@��7�@�K���|,��B�fE/����'EҠZ3�T0 k� �&��&	E1 4#Q&�1D"3Q  ��    � < �dX@��6�H�K���|,��B�fE/����&EҠZ3�T0 k� �%��%	E1 4#Q&�1D"3Q  ��    � < �dT@��4�\�(K���|,��B�(eE/��	� %E�Z3�T0 k� �#��#	E1 4#Q&�1D"3Q  ��    � < �                                                                                                                                                                            � � �  �  �  d A�  �K����  �      6 \��^, ]�%�%� �  �� g��   I I   � �V�     g� �U    ���             $	 Z           �`�    ���  (
	           [��  : :     �
��     [�D
��    �d             !		 Z          ֐�    ���   
	           l��   M M      �H     mr� �!    ���   	        O Z �        !��     ���   8	 

          EW            Е�     EW ��F      �   
          9  Z            p     ���  0
3
          E�z   � �
	   / ���     E�n ���    L�              < Z           @�    ���   H


          �  ��     C�	�     ��	�                             ����              �  ���    		 5 	           ����          W ��u    ���x ��    �| �            
 
 a��           �     ��@   0
&


         ���       k ��    ��� ��[    � �             
 
 \��          �P     ��@   (
 
          ��Q�        ���    ��E( ��0     �f               6��          �     ��@   0	
          �҃�        �3    �ҍ�*    �j y                     �         	 �      ��@   H	$
          z5�         � k��     z^� k�    ����             ` �         
  *p     ��J   03 
           8����     �!�#     8��!ҙ      �                    �  �              )  ��@    P		 5                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          D@�  ��        � ���     E@� �/?      � "                 x                j  �       �                          D    ��        � �       E   �           "                                                �                          �
 � � �� � � � k!�� � �   	  
            
  �   � �w ���E       ބ �c` /� \� /� \� 0 \� � _    _@ �� 0\� �  ]@ �D ]����  ����. ����< ����J ����X ����J ����X � �� ]  :d ]  
�| W� 
�\ X  �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }����� ����� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����    3���   ������  
�fD
��L���"����D"� �  " `   J jF��     �j   
��
��
���    "�j��" " �
� �  �  
�  E    ��     � �       E    ��     � �       z    ��     � k          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �3333      ��T ���        �GT ��        �        ��        �        ��        �    ��
     E d�~��        ��                         T�) ,  	�����                                     �                 ����             E ����&��   3                 20 Luc Robitaille                                                                                   2  2     �C
�:Hk �] k� �#kk n;ks ^C � � �	C0 �
C%	 �C1 � C) �C/ � C7 � C8 �C9 � C; � C< �B�+ � B�* � B�# � B�5 �J� � J�$ � J� �	� � �	� � �� � �� � �c� � � c� � � k� � �!k� � �"k� � #k� �,$"�, %"�&�'
�,("�, )"�*"�+*� � ,"N u �-"% � � ."@ � � /*N � 0*HE � 1*PmH  *'u � 3*O � 4*Sm � 5*u � 6*SM � 7*U � 8*RU � 9*Qm � :*P] �;*7m �<*+u �=*;m � >*Q}  )�m                                                                                                                                                                                                                         �� R         �     @ 
             Z P E ]  ��        
            ������������������������������������� ���������	�
���������                                                                                          ��    ���   ������������ �!�"�#�$�k�l�'�(�)�*�+�m�n�o�/�0�1�2�p�q�r�6�7�1�2�N�s�O�;�<�1�2�=�a�?�2�@�A�B�C�t�E�B�F   �4, E    3�  Q A����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             
        t    #    �� 
İJ      �                             ������������������������������������������������������                                                                                                                                        ����  �  �                                           ���������������� ���������������������   ������� ��������� ������� ������� ����������������������� � ���������� ���� ��� � ��  ������������������ �������������������  ������������� ������������������������������������ ���� ��  ������������ ������� �������                                    �    9     �� ��J      B�                             ������������������������������������������������������                                                                       
                                                                      ����  ��                                             � ������������ �������� ������ �� �� ������� ���������  �� ������������� ����������� �� ���� ������������� �������� �������� ����� �����  ���� �������������������� ����� � ������������� � ��� �����������������������  ������                                                                                                                                                                                                                                                                                                                            �              


             �  }�           �          L-           Y                                                        c      6�  K��������  �����������������������������������������������������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � �� �\                                                                                                                                                                                                                                                                                           )n)nY  
�        l            l                              m                                                                                                                                                                                                                                                                                                                                                                                                          > �  >�  Z�  @<  )#�  EZm.  �N ��� �~��H�~��� ����������������{������                 2   n q        $   �   & QW  �   W                  �                                                                                                                                                                                                                                                                                                                                        K K    �                       !��                                                                                                                                                                                                                            Z   �� �~ ���      �� M      ���������������� ���������������������   ������� ��������� ������� ������� ����������������������� � ���������� ���� ��� � ��  ������������������ �������������������  ������������� ������������������������������������ ���� ��  ������������ ������� �������� ������������ �������� ������ �� �� ������� ���������  �� ������������� ����������� �� ���� ������������� �������� �������� ����� �����  ���� �������������������� ����� � ������������� � ��� �����������������������  ������              $����������������UUUU�����UUU�U{�����������������UUUW����x�����w�����������������UUuU������wxwwww����������������WwwU�������wwwwx����������������UUUU����w�xw�w������������������Uuww���uUw��uU���Uz��uz��Wz��wzu�wYW�wxw�uxwwuW���������wx��UUwwX�xuy����u������wwww�wwwwwwwwwwwUUwWuUuu�UWW�wwwwy��x���x���ww�uwuuwwx��x�����Y����������w��www�wwwy��wyx�wyx��x�U���U���U���uy��u���u��uu��uU���wx��wxxwuW�WuuxU�uWW�UUU�uWu��W�y���wx�ww��wxx����wwwwwWwwwwwuW��ww��wx��w��xww��WwxUW�wWW�wy����w����������x�www��xwx�w��w�Ww����w��xwx�xwwwx�xwww��ww�wwwwwww�Wy�x�xuw��UwuwWwuwWwxwX�xwW�wuW�z�u�Y�u�X�u�U��yUU�Uuw�yUX��UX�uWwuWuwWwUwwUUUwUUWUUUUuUUWWUUWwwuW�WUW�XUuwx�UXx�Uxwwwxww�xww����ww��UwuwwW��ww��ww��ww��xw��xwwwwwwwwwwwwxwwwxuwwxwwwwUwwwWwwwwywX��yWx�Xxy�W��uXYwWuZ��u��w���ux���w���U���U���U���u���UZ��UWUUwWuUUU�Uu��Uw��UWx�UUW��UU��UUwwwxUwww��wx��������x���w���Ux�wx�wwwwww���w���U��ww��ww�wwwuwwwWwwxWwwywww�wwx�ww��xx��wx��w����WU��WY��uY��Wx��Wy�Uxz�Xw��Xw�W���W���U��������������������������UUW�uUUX�U�U�W�uWW��WU���u���WUUUWUUwuuwwwwx��wwx�wwwwwwwwuwwwWuwwWwwwuwwx�ww�wwwx�w�xxw��wx��xw�Uw��W���Xx�U��uW��UxwUWwwUwww�w�W�x�W�y�wx��wx�Wwx�Wyz�wz��x�q��    2      A    �  E                       M     �  ���������J'    ��     F�      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��  � ��     � ��   	 ��   p �� �� ��  � ��     �� ��  ��   	 ��   p �� ��  � ��  �` ��   ��    ��   � �� �� �z   ����� �$ ��  �� �� ��   	 �� �� ��  �� �� �  �� �� �z � ���    9  ��9       �  ��   ���� e����J   g���        f ^�         �� � 3            ��^��������J���J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                         E  �\       U TUTQ�T\�jA���̪������ UTDDEUU�����j������������������DUP UUTD�����v����������������    U�UPUDDE��\����������������        U   TE ��@ x�@ �lE �|U  E� \� �Q� _ǪE�L��\��\�������������������E�lTP��E ��P �����������UDL�_UL�_L�UL�L�̪�������U������D���EU��E��E���E���������z��Q�j�T_�z �_�  T\  E��U ��T ����|��E |P �E  @  \��\��\��Ez� Oʪ UǪ \� Eʪ�P ��E �|�P���D��lϪ�����������L��L��L�UUL�QDL�_���Ua��̪��w���E��EU��E���E��DU�����wz��   �  �E �ETOQ���j����������UO  �T  ��P ��O ��� �����O���E  T\  E   T                   ����Ǫ��\ʪ�E\ʪUE\� UDU  UT    ����������������z������DUUUUTD�������������������|���UUTDDUU�����������̧|�T�TUUDP U       ��TQ�TE TE  E                   wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwtwwwCwwt1wwCwt1wC�t1��C1����������""""���������������!���""!����,���ww��7����������������wwwwwwwwwwwwwwwwwwww7wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwws��w1wt1�wC�t1��s��s��s������"$��Gw�!������������L���q��"r��������!�����!ww�r�w�ww!�wwrwwwwwwqwwwrwwww�7ww�ww�ww��7w��w���G��'!wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  " ! " ""  "!  " ! " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  " ! " ""  "!  " ! " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  " ! " ""  "!  " ! " ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                       b}z�gg��j�� 
�� 	�� �� �� 
�� �� ��̻�"+��" 4"  4   D   H   H   �  +  ""    ��       ��  �٠ �ڛ ̸� ̻� �̽ �̀ �ɀ ��0 ��C 4�T H�T H�D �T@ �T  �C  �0  ɚ  ��� ��� �" �"  �"�                 �� �� �� {�             �   �  " � "�� � �  ��                                        �   �   �   "   "   "  !�    ��                              �                        ��"� �"� ����            �     "   "                   �     �                         � ".��".��/����  �                                                                                                                                                      � �� �������ۛ˽���� �ͼ ��+ �""�B.�R#Z�C U�D �T Z� �; � �� ��� ��  ��� ˽� �wp �&  �vp �w� ��� ˙� ̻� �۰ �ِ ��� Ш� �� >�" 3��.30" ��  �   �                �"/ "" ""  ��  ��                       .  .  "   "           �   �   �   �   �   �   �@      �    �  �   �""��""����                          �� �� ��               �  �  �     "   "                      �۰ ̽  �̰ ̻� ˸� ��U@��T@UUUJ             �  �˰ ��� �wp �&                                                                                                                                                                   ˰ ̻ ̻ �� {�  �� 
�� ��� ��� ������
���	��ܻ̍ݻ���"� 8"  8  �  D�  H�  X�  ��  �   �          "  "     �                        ��  ��� �̺�̻����ۻ�˽��̽��̝ ̙� �30 �EP �U@ �T0 EC0 T3  C:  K�  �"  �"/ ����˽� �"� "" �""� � �� ��      �   �  .�  ."  �               �                         "   "  !�    ��                ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                          �    ��                                                                                                                                                      "  "(��ȩ�ܚ��ۊ����� ��  �   �   �   �   �� ��� ̻� ˽� ��� �w� �������������������������� �̻ ���         �   �       �   �   "" �+� Ȼ� ɫ� ɨ� ��                �� �I��3 ��D 
UD 
UD TD  T�  ˸  ��  �� ̰ �+ ��"/ �"/  ����  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� �   �".  .                            �   �    �   �       �   �   �                .      ���.�                     ���                                                                                                                                                                                            "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             �"  �""� "�    �     �                                                                                                                                                                                                    �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �   �ڀ �Ͱ ��� �� �̰��˰ ��� ���                     �                               �   �   ��  ���   ˰  ̹  ��@ ��UP�EEXDTD�                                                                                                                                                                  �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �   �   �   �   �@      �    �  �   �""��""����     �"  �                        .   .   �                                      �".��".  ���    �                    ".  ".  ���     ��   �  ��  �  �  �         � ".��".��/����  �                                                                                                                                                      �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp��& ��vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �" �"" �"   �                    .   .   �                  �   �                           �� " ��   "                  �".��".  ���    � �EU �E  
�   �               �"�!/"�  �                                                                                                                                                                                 �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���            �    �  �   �""��""����         �  ��  ��  ww  &'  vv  w                   �   �                      �".��".  ���    �                    ".  ".  ���     ��   �  ��  �  �  �         � ".��".��/����  �                                �   "                                                                                                  �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���        T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ��"� �"� ����                            ".  ".  ��� ���                                                �   ���                            �   "                                                                                                    �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �"  "�  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �              .  ". ""  "    � ���                                                                                                                                                                                                                     �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ���������""��""��""�����        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                   2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD           	 
          
        ((((((( 
	(((( GwDGwqwDDwtwwww3333DDDD             ! " # $ % & '   ( $ % ) ! " # * ('(&(%($(#("(! (((""""����������A��I��I + , -   . / 9 1  	 2         3       4 (((((((2	19/(.(-(,(+""""�����A�DA�I��I� 5 6   7   8 9 1 :   $ % ) ! " #   ; ) ! " # $ % ) (#("(!()(%($ :198(((7(6(5""""��������I���I���I���I���    <     = 8 9 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>198(=((( (<MAMAMMMM�M�M����3333DDDD L  . M + , N    O P Q R S S S T S S S T S S 0 Z S ST S S ST S S SRQPO(( (N(,(+(M(.LD�����MD��M����3333DDDD  7  N 5 U V W X Y S S [ S S S _ S S S _ S S \ ] S S_ S S S_ S S S[ S SY(X(W(V(U(5(N((7���4���4���4���4���4���43334DDDD  `  V    a b c S S f g h i j i i i j i i ^ d i ij i i ij ihgf S Scb(a(((V((`""""wwwwqqqqwGwGGG 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
""""wwwwwwqqDAwG w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw������������������333DDD w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xwwM��M��D��M����������3333DDDD + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+DD��D�M��D����3333DDDD � W  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ������ ���((W(�""""������DH�H� � a � l � � � � � �������� � �� � � � � � ���	����� � � �� �������l(�(a(�""""�������H�H��D �  � y � � � � � � � � � � � � � � � �� ��������� � � � � � � � � ������y(�(�""""��������H��H��H��H� = l �  � � � � � � � � � � ��� � � � � �������� � � � ��� � � � ������((�l(=DD������L��DL����3333DDDD    �  � � � � � � � � � ������ � � � � � ���� � � � ������ � � �����((�(( L�A�AAD��DL�����3333DDDD x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���4���4���4L��4L��4���43334DDDD w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww""""���������M�MMM  � w w � � � � � � � � � ��	� � � ��� � � � � � � � � � � ��	� � � ��� �����ww�(""""�������A��AA �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((���������������333DDD ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`I��I����������������3333DDDD M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M��A���I��I���I�����3333DDDD � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(�""""������������������������ � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(�""""������D�D��� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5""""������������������������ x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�xwqwwqwwwwwqwwwDwwww3333DDDD w � � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxwwqqwwwDDwtGwwww3333DDDD � � � i i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+www4www4www4www4www4www43334DDDD W � � u u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(�""""wwwwwwqwwwqwqwq333333333333333333333333333333333333333333333333333333333333����  
�fD
��L���"���""""wwwwwwwDwGwA�D"� �  " `   J jF� ����
��� �����
���� ����
��� �����
��� 0 q�A�L�L�L��L���333DDDLDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDDC
�:Hk �] k� �#kk n;ks ^ � �	C	C!	 �
C%	 �C1 � C) �C/ � C7 � C8 �C9 � C; � C< �B�+ � B�* � B�# � B�5 �J� � J�$ � J� �	� � �	� � �� � �� � �c� � � c� � � k� � �!k� � �"k� � #k� �,$"�, %"�&�'
�,("�, )"�*"�+*� � ,"N u �-"% � � ."@ � � /*N � 0*HE � 1*PmH  *'u � 3*O � 4*Sm � 5*u � 6*SM � 7*U � 8*RU � 9*Qm � :*P] �;*7m �<*+u �=*;m � >*Q}  )�m3333DDDDAqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD������� �!�"�����������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ���#�$�k�l�'�(�)�����������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ���*�+�m�n�o�/�0�����������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE���1�2�p�q�r�6�7�����������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD���1�2�N�s�O�;�<�����������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD���1�2�=�a�?�2�@�����������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD���A�B�C�t�E�B�F�����������������������""""��������AAAHA""""�������DDA��H��������������������������������������������""""���������DAAAq""""�����ADHA��H�� �2�H�T�L���]�L�Y����������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� �� ��>�O�L�V�Y�L�U��1�S�L�\�Y�`�������8�>�7���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� ����>�L�L�T�\��=�L�S�H�U�U�L��������>��<���""""������A�D��I��""""�������D����� ����7�\�J��<�V�I�P�[�H�P�S�S�L�������8�>�7���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �>��<������A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �8�>�7�����""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,�����������DDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II�""""������D""""������IADD���I""""��������D��""""�������I��I�I�I�""""�������A�D�II�I""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            