GST@�                                                            \     �                                                ���     �  ��  y         ����e ����ʳ������������������        �g      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"��   " `  J  jF��    "�j "����
��
��     �j�� 
   ��
  d�                                                                              ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������=?  00  45  18                         
     
                ��  �4  �  ��                  �Y  	          : �����������������������������������������������������������������������������                                  0       �   @  &   �   �                                                                                 '        )n)n1n  	�Y    �0   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E 0 �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    D2D�ǻ@�?'�IS�Y|C����x_B����?7�"���T0 k� S��W�&51D"3Q��0 D 3Q ��    ��� �D2D�˼@�?'�IW�Y|C����x_B����?7�"���T0 k� S��W�&51D"3Q��0 D 3Q ��    ��� �41D�ϼ@�?'�I_�Y|C����x_B����/3�"���T0 k� O��S�&51D"3Q��0 D 3Q ��    ��� �4 1D�Ͻ@�?'�Ic�Y|C����x_B����//�"���T0 k� K��O�&51D"3Q��0 D 3Q ��    ��� �3�0D�ӽ@�?'�Ik�Y|C����x_2����//�"���T0 k� �G��K�&51D"3Q��0 D 3Q ��    ��� �3�0D�׾@�?'�I"o�Y|C����x_2�����/+�"���T0 k� �G��K�&51D"3Q��0 D 3Q ��    ��� �3�/D�ۿ@�?#�I"s�Y|C����x_2�����/+�c��T0 k� �C��G�&51D"3Q��0 D 3Q ��    ��� �C�/D���@�?#�I"�Y|C����x_2����/+�c��T0 k� �;��?�&51D"3Q��0 D 3Q ��    ��� �C�/D���A?#�I"��Y|C����x_B����/+�c��T0 k� �;��?�&51D"3Q��0 D 3Q ��    ��� �C�/D���A?#�I��Y|C���x_B���ۭ+�c��T0 k� �7��;�&51D"3Q��0 D 3Q ��    ��� �C�/D���A?#�I��Y|C��w��x_B���׭+�c��T0 k� �3��7�&51D"3Q��0 D 3Q ��    ��� �C�/E���A?#�I��Y|C��o��x_B���Ϯ+�c��T0 k� �/��3�&51D"3Q��0 D 3Q ��    ��� �C�/E���A?#�I��Y|C��g��x_B���Ǯ+�c��T0 k� �+��/�&51D"3Q��0 D 3Q ��    ��� �C�/E���A?#�I��Y|C��[��x_ ���ҿ�+�c��T0 k� �+��/�&51D"3Q��0 D 3Q ��    ��� �C�/E���A?#�I"��Y|C��S��x_ ���һ��+�c��T0 k� �'��+�&51D"3Q��0 D 3Q ��    ��� �3�/E���A?�I"��Y|C��K��x_ ���ҳ��+�c��T0 k� �#��'�&51D"3Q��0 D 3Q ��    ��� �3�0Es�A?�I"��Y|C��C��x_ ���ҫ��+�c��T0 k� ���#�&51D"3Q��0 D 3Q ��    ��� �3�0Es�A?�I"��Y|C��C��x_ ���ҫ��/�c��T0 k� ���#�&51D"3Q��0 D 3Q ��    ��� �3�0Es�A?�I"��Y|C��?��x_ ���⫰�/�c��T0 k� ���&51D"3Q��0 D 3Q ��    ��� �3�1Es�A?�I��Y|C��;��x_ ���⣰�/�c��T0 k� ���&51D"3Q��0 D 3Q ��    ��� �3�1Es�A?�I��Y|C��7��x_ ���⛰�3�c��T0 k� ���&51D"3Q��0 D 3Q ��    ��� �#�2Es�A?�I��Y|C��3��x_ ���⓱�3�c��T0 k� ���&51D"3Q��0 D 3Q ��    ��� �#�3Ec�A?�I��Y|C��/��x_ ���⋱�7�c��T0 k� ���&51D"3Q��0 D 3Q ��    ��� �#�3Ec�A?�I��Y|C��+��x_ ���R���7�c��T0 k� ���&51D"3Q��0 D 3Q ��    ��� �#�4Ec�A?�I"��Y|C��#��x_ ���R{��;�c��T0 k� ���&51D"3Q��0 D 3Q  ��    ��� �#�4Ec�A?�I"��Y|C����x_ ���Rs��;�c��T0 k� ���&51D"3Q��0 D 3Q  ��    ��� �#�5Ec�A?�I"��Y|C����x_ ���Rk��?�c��T0 k� ���&51D"3Q��0 D 3Q  -�    ��� �#�6Ec�A?�I"��Y|C����x_ ���Rc��C�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� ��7Ec�A?�I"��Y|C����x_ ���R[��C�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ��7Ec�A?�B���Y|C����x_ ����S��G�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ��8Ec�A?�B���Y|C����x_³��K��K�c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� ��9Ec�A?�B���Y|C����x_³��?��O�c��T0 k� �����&51D"3Q��0 D 3Q ��    ��� ��:Ec�A?�B���Y|C����x_³��7��S�c��T0 k� ����&51D"3Q��0 D 3Q ��    ��� ��:Ec�A?�B���Y|C����x_³��/��W�c��T0 k� ����&51D"3Q��0 D 3Q ��    ��� ��;Ec�A?�O��Y|C����x_³��'��[�c��T0 k� ����&51D"3Q��0 D 3Q ��    ��� ���;Ec�A?�O��Y|C�����x_³����_�c��T0 k� ����&51D"3Q��0 D 3Q ��    ��� ���<Eb��A?�O��Y|C�����x_¯����c�c��T0 k� ����&51D"3Q��0 D 3Q ��    ��� ���=Eb��A?�O��Y|C�����x_¯����g�c��T0 k� �ߝ��&51D"3Q��0 D 3Q ��    ��� ���=Eb��A?�O��Y|C�����x_ү����k�c��T0 k� �ߜ��&51D"3Q��0 D 3Q �    ��� ���=Eb��A?�O��Y|C�����x_ү�����s�c��T0 k� �ۛ�ߛ&51D"3Q��0 D 3Q �    ��� ���>Eb��A?�O��Y|C�����x_ҫ����w�c��T0 k� �ӛ�כ&51D"3Q��0 D 3Q ��    ��� ���>ER��A?�O��Y|C�2���x^ҫ����{�c��T0 k� �˛�ϛ&51D"3Q��0 D 3Q ��    ��� ���?ER��A?�O��Y|C�2��x^ҧ�����c��T0 k� ����Û&51D"3Q��0 D 3Q ��    ��� ���@ER��A?�O��Y|C�2��x^���ϳϋ�c��T0 k� �����&51D"3Q��0 D 3Q ��    ��� �C�@ER��A?�O��Y|C�2��x]� �ǲϏ�c��T0 k� �����&51D"3Q��0 D 3Q ��    ��� �C�AP���A?�O��Y|C�2��x]�ῲߗ�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �C�AP���A?�O��Y|C�2��x\�ᷲߛ�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �C�AP���A	?�O��Y|C�2��x[�᯲ߣ�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �C�BP���A	?�O��Y|C�2��x[�᧲ߧ�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �C�BP���A	?�O��Y|C�2��xZ�៲߯�c��T0 k� {���&51D"3Q��0 D 3Q  /�    ��� �C�CP���A
?�O��Y|C�2��xY�ᗱ߷�c��T0 k� s��w�&51D"3Q��0 D 3Q  ��    ��� �C�CP�� A
?�O��Y|C�2��xY�ዱ߻�c��T0 k� k��o�&51D"3Q��0 D 3Q  ��    ��� �C�CP��A?�O��Y|C�B��xX�ჱ���c��T0 k� c��g�&51D"3Q��0 D 3Q  ��    ��� �C�DP��A?�O��Y|C�B��xW�	�{����c��T0 k� �W��[�&51D"3Q��0 D 3Q  ��    ��� �C�DP��A ?�O��Y|C�B��xV�
�s����c��T0 k� �[��_�&51D"3Q��0 D 3Q  ��    ��� �C�DP��A ?�O��Y|C�B߯�xU��k����c��T0 k� �_��c�&51D"3Q��0 D 3Q  ��    ��� �C�EP��A ?�O��Y|C�B߮�xT��c����c��T0 k� �_��c�&51D"3Q��0 D 3Q  ��    ��� �C�EP��A ?�@��Y|C�B߮�xS"��[����c��T0 k� �[��_�&51D"3Q��0 D 3Q  ��    ��� �C�EP��A$?�@��Y|C�Bۭ�xQ"��S����c��T0 k� �W��[�&51D"3Q��0 D 3Q  ��    ��� �C�FP��A$?�@��Y|C�Bۭ�xP"|aK����c��T0 k� �C��G�&51D"3Q��0 D 3Q  ��    ��� �C�FP��	A$?�@��Y|C�B۬RxO"|aC����c��T0 k� �/��3�&51D"3Q��0 D 3Q  ��    ��� �C�FP��	A$?�@��Y|C�B׬RxN"xa;���c��T0 k� ���#�&51D"3Q��0 D 3Q  ��    ��� �C�GP��
A$?�@��Y|C�B׫RxM"xa3���c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�GC�A(?�@��Y|C�B׫RxL"ta+���c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�GC�A(?�@��Y|C�BӪRxK"ta���c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �C�HC�A(?�@��Y|C�BӪRxI"pa��#�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�HC�A(?�@��Y|C�BөRxH"pa��+�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�HC�A,?�@��Y|C�BөRxG"lQ��3�c��T0 k� �ߜ��&51D"3Q��0 D 3Q  ��    ��� �C�IAR�A,?�@��Y|C�BϩRxF"lP���;�c��T0 k� �ۡ�ߡ&51D"3Q��0 D 3Q  ��    ��� �C�IAR�A,?�@��Y|C�BϨRxE"hP���C�c��T0 k� �Ӥ�פ&51D"3Q��0 D 3Q  ��    ��� �C�IAR�A,?�@��Y|C�BϨRxD"hP��K�c��T0 k� �˦�Ϧ&51D"3Q��0 D 3Q  ��    ��� �C�IAR�A,O�@��Y|C�B˧RxC"dP��S�c��T0 k� �è�Ǩ&51D"3Q��0 D 3Q  ��    ��� �C�JAR�A0O�@��Y|C�B˧RxB"dPߥ�[�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�JAR�A0O�@��Y|C�B˧RxA"`Pפ�c�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�JAR�A0O�@��Y|C�B˦bx@"`PϤ�k�c��T0 k� ����&51D"3Q��0 D 3Q  ��   ��� �C�KAR�A0O�@��Y|C�BǦbx?"\Pǣ�s�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�KAR�A0O�@��Y|C�Bǥbx?"\P���{�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�KAR�A4O�@��Y|C�Bǥbx>"XP��
@��c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�KAR�A4O�@��Y|C�Bǥbx="XP��
@��c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �C�LAR�A4O�@��Y|C�Bäbx<"TP��
@��c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �C�LAR�A4�@��Y|C�Bäbx;"T@��
@��c��T0 k� �{���&51D"3Q��0 D 3Q  ��   ��� �C�LAR�A4�@��Y|C�Bäbx:"P@��
@��c��T0 k� �s��w�&51D"3Q��0 D 3Q  ��    ��� �C�LAR�A4�@��Y|C�Bãbx9"P @��0��c��T0 k� �k��o�&51D"3Q��0 D 3Q  ��    ��� �C�LAR�A8�@��Y|C�Bãbx9"P @��0��c��T0 k� �c��g�&51D"3Q��0 D 3Q  ��    ��� �C�MAR�A8�@��Y|C�B��bx8"L!@{�0��c��T0 k� �[��_�&51D"3Q��0 D 3Q  ��    ��� �C�MAR�A8�@��Y|C�B��bx7"L!@s�0��c��T0 k� �S��W�&51D"3Q��0 D 3Q  ��    ��� �C�MAR�A8�@��Y|C�B��bx6"H"@k�0��c��T0 k� �G��K�&51D"3Q��0 D 3Q  ��    ��� �C�MAR�A8�@��Y|C�B��bx5"H#`c�0��c��T0 k� �?��C�&51D"3Q��0 D 3Q  ��    ��� �C�NAR�A8�@��Y|C�B��bx5"D#`[�0��c��T0 k� �7��;�&51D"3Q��0 D 3Q  ��    ��� �C�NAR�A8 �@��a�C�B��bx4"D$`S�0��c��T0 k� �/��3�&51D"3Q��0 D 3Q  ��    ��� �C�NAR�A< �@��a�C�B��bx3"D$`K�@��c��T0 k� �'��+�&51D"3Q��0 D 3Q  ��    ��� �C�NAR�A< �@��a�C�B��bx2"@%`C�@��c��T0 k� ���#�&51D"3Q��0 D 3Q  ��    ��� �C�NAR�A< �@��a�C�B��bx2"@%`;�@��c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�OAR�A< �@��a�C�2��bx1"@&P3�@��c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�OAR|A< �@��a�C�2��bx0"<'P/�@��c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�OAR|A< �@��a�C�2��bx0"<'P'�@��c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�OAR| A< �@��a�C�2��bx0"8(P�A�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �C�OARx A@ �@��a�C�2��bx0"8(P�A�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �C�PARx A@ �@��a�C�2��bx08)@�A�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�PARx A@ �@��a�C�R��bx04)@�A�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�PARt A@ �@��Y|C�R��bx04*@�A�c��T0 k� �ߪ��&51D"3Q��0 D 3Q  ��    ��� �C�PARt A@ �@��Y|C�R��bx04*O��A'�c��T0 k� �ת�۪&51D"3Q��0 D 3Q  ��    ��� �C�PARt A@ �@��Y|C�R��bt00*O��A+�c��T0 k� �Ӫ�ת&51D"3Q��0 D 3Q  ��    ��� �C�QARp A@ �@��Y|C�R��bt00+o�A3�c��T0 k� �˩�ϩ&51D"3Q��0 D 3Q  ��    ��� �C�QARp AD �@��Y|C�B��bt0�0+o�A;�c��T0 k� �ǩ�˩&51D"3Q��0 D 3Q  ��    ��� �C�QARp AD �@��Y|C�B��bt0�,,o�AC�c��T0 k� ����é&51D"3Q��0 D 3Q  ��   ��� �C�QARp AD �@��Y|C�B��bt0�,,oߚAG�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �C�QARl AD �@��Y|C�B��bt0�(-oךAO�c��T0 k� ������&51D"3Q��0 D 3Q �    ��� �C�QARl AD �@��Y|C�B��bt0�(-ӚQW�c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�QARl AD �@��Y|C����bt0�$-˙Q_�c��T0 k� �{���&51D"3Q��0 D 3Q ��    ��� �C�RARh AD �@��Y|C����bt0�$-ǙQc�c��T0 k� �g��k�&51D"3Q��0 D 3Q ��    ��� �C�RARh AD �@��a�C����bt0� .��Qk�c��T0 k� �S��W�&51D"3Q��0 D 3Q ��    ��� �C�RARh AD �@��a�C����bt0�.��Qs�c��T0 k� �?��C�&51D"3Q��0 D 3Q ��    ��� �C�RARh AH �@��a�C����bt0�.���Q{�c��T0 k� �+��/�&51D"3Q��0 D 3Q ��    ��� �C�RARd AH �@��a�C����bt0�.���Q�c��T0 k� ����&51D"3Q��0 D 3Q	 ��    ��� �C�RARd AH �@��a�C����Rt0�.���Q��c��T0 k� ����&51D"3Q��0 D 3Q ��    ��� �C�SARd AH �@��a�C����Rt0�.���Q��c��T0 k� ����&51D"3Q��0 D 3Q ��    ��� �C�SARd AH �@��a�C����Rt0�-���Q��c��T0 k� �ۻ�߻&51D"3Q��0 D 3Q ��   ��� �C�SAR` AH �@��a�C����Rp0�-���
џ�c��T0 k� �˽�Ͻ&51D"3Q��0 D 3Q ��    ��� �C�SAR` AH �@��a�C����Rp0�-���
ѣ�c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�SAR`AH �@��a�C����Rp0�,���
ѫ�c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�SAR`AH �@��a�C�����p0�,���
ѳ�c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�SAR`AH �@��Y|C�����p0�,���
ѻ�c��T0 k� �{���&51D"3Q��0 D 3Q ��    ��� �C�SAR\AL �@��Y|C�����p0�+���
�úc��T0 k� �g��k�&51D"3Q��0 D 3Q ��    ��� �C�TAR\AL �@��Y|C�����p/�+��
�˹c��T0 k� �S��W�&51D"3Q��0 D 3Q ��    ��� �C�TAR\AL �@��Y|C�����p/� *�{�
�ϸc��T0 k� �?��C�&51D"3Q��0 D 3Q ��    ��� �C�TAR\AL �@��Y|C�����p/� )�w�
�׸c��T0 k� �+��/�&51D"3Q��0 D 3Q ��    ��� �C�TAR\AL �@��Y|C�����p/��)�s�
�߷c��T0 k� ����&51D"3Q��0 D 3Q ��    ��� �C�TARXAL �@��Y|C����p/��(�k�
��c��T0 k� ����&51D"3Q��0 D 3Q ��    ��� �C�TARXAL �@��Y|C����p/��'�g�
��c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�TARXAL �@��Y|C����p.��&�c���c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�TARTAL �@��Y|C����p.��&�_���c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�UARTAL �@��Y|C����p.��%�[��c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�UARTAL �@��Y|C����p.��$�W��c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�UARTAL �@��Y|C����p-��#S��c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�UARPAP �@��Y|C�R���p-��"O��c��T0 k� �w��{�&51D"3Q��0 D 3Q ��    ��� �C�UARPAP �@��Y|C�R���p,��!K��c��T0 k� �c��g�&51D"3Q��0 D 3Q ��    ��� �C�UARPAP �@��Y|C�R���p+��K�'�c��T0 k� �O��S�&51D"3Q��0 D 3Q ��    ��� �C�UARPAP �@��Y|C�R���p+��G�+�c��T0 k� �;��?�&51D"3Q��0 D 3Q ��    ��� �C�UARLAP �@��Y|C�R��Rp+��C�3�c��T0 k� �'��+�&51D"3Q��0 D 3Q ��    ��� �C�UARLAP �@��Y|C�R��Rt*��?�7�c��T0 k� ����&51D"3Q��0 D 3Q ��    ��� �C�VARLAP  �@��Y|C�R��Rt*���;�?�c��T0 k� �����&51D"3Q��0 D 3Q ��    ��� �C�VARHAP  �@��Y|C�R��Rt)���7�C�c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�VARHAP  �@��Y|C�R��Rt)���3�K�c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�VARHAP  �@��Y|C�R��Rt(���/�"O�c��T0 k� ������&51D"3Q��0 D 3Q ��    ��� �C�VARDAP  �@��Y|C�R��Rt(���/�"W�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �C�VARDAP  �@��Y|C�R��Rt'���+�"[�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �C�VARDAP  �@��Y|C�R��Rt&���'�"c�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �C�VARDAP  �@��Y|C�R��Rt&���#�"g�c��T0 k� �s��w�&51D"3Q��0 D 3Q! ��    ��� �C�VAR@AT  �@��Y|C�R��Rt%����"g�c��T0 k� �_��c�&51D"3Q��0 D 3Q! ��    ��� �C�VAR@AT  �@��Y|C�R��Rx%����"g�c��T0 k� �K��O�&51D"3Q��0 D 3Q! ��    ��� �C�VAR@AT! �@��Y|C�R��Rx$���"k�c��T0 k� �7��;�&51D"3Q��0 D 3Q! ��    ��� �C�WAR@AT! �@��Y|C�R��Rx$��
�"o�c��T0 k� �#��'�&51D"3Q��0 D 3Q! ��    ��� �C�WAR<AT! �@��Y|C�R��bx#��	�"s�c��T0 k� ����&51D"3Q��0 D 3Q! ��    ��� �C�WAR<AT! �@��Y|C�R��bx#���"w�c��T0 k� ������&51D"3Q��0 D 3Q" ��    ��� �C�WAR<AT! �@��Y|C�R��bx"���"{�c��T0 k� ������&51D"3Q��0 D 3Q" ��    ��� �C�WAR<AT! �@��Y|C�R��bx"���"{�c��T0 k� ������&51D"3Q��0 D 3Q" ��    ��� �C�WAR8AT! �@��Y|C�R��bx!���"�c��T0 k� ������&51D"3Q��0 D 3Q" ��    ��� �C�WAR8AT! �@��Y|C�R��bx!�� �"��c��T0 k� ������&51D"3Q��0 D 3Q" ��    ��� �C�WAR8AT! �@��Y|C�R��bx!���"��c��T0 k� �� �� &51D"3Q��0 D 3Q" ��    ��� �C�WAR8AT! �@��Y|C�R��bx ����"��c��T0 k� ����&51D"3Q��0 D 3Q! ��    ��� �C�WAR4AT! �@��Y|C�R��bx �����"��c��T0 k� �l �&51D"3Q��0 D 3Q! ��    ��� �C�WAR4AT" �@��Y|C�R��bx�����"��c��T0 k� �X �&51D"3Q��0 D 3Q! ��    ��� �C�WAR4AT" �@��Y|C�R��b|�����"��c��T0 k� �D �&51D"3Q��0 D 3Q! ��    ��� �C�WAR4AT" �@��Y|C���b|�����"��c��T0 k� �0 �&51D"3Q��0 D 3Q! ��   ��� �C�XAR4AT" �@��Y|C���b|�����"��c��T0 k� �
 �&51D"3Q��0 D 3Q! ��    ��� �C�XAR0AT" �@��Y|C���b|����"��c��T0 k� � �&51D"3Q��0 D 3Q! ��    ��� �C�XAR0AX" �@��Y|C���b|����"��c��T0 k� �� �&51D"3Q��0 D 3Q  ��    ��� �C�XAR0AX" �@��Y|C���b|����"��c��T0 k� �� �&51D"3Q��0 D 3Q  ��    ��� �C�XAR0AX" �@��Y|C� ���b|����"��c��T0 k� �� �&51D"3Q��0 D 3Q  ��    ��� �C�XAR0AX" �@��Y|C� ���b|����"��c��T0 k� �� �&51D"3Q��0 D 3Q ��    ��� �C�XAR,AX" �@��Y|C� ���b|����"��c��T0 k� �� �&51D"3Q��0 D 3Q ��    ��� �C�XAR,AX" �@��Y|C� ���b|����"��c��T0 k� �� �&51D"3Q��0 D 3Q ��    ��� �C�XAR,AX" �@��Y|C� ���b|����"��c��T0 k� �| �&51D"3Q��0 D 3Q ��    ��� �C�XAR,AX" �@��Y|C�ҋ�b|q���"��c��T0 k� �h �&51D"3Q��0 D 3Q ��    ��� �C�XAR,AX" �@��Y|C�ҋ�b|q��ߓ"��c��T0 k� �T �&51D"3Q��0 D 3Q ��    ��� �C�XAR(AX# �@��Y|C�ҋ�b|q��ߓ"��c��T0 k� �@ �&51D"3Q��0 D 3Q ��    ��� �C�XAR(AX# �@��Y|C�ҋ�b|q��ۓ"��c��T0 k� �, �&51D"3Q��0 D 3Q ��    ��� �C�XAR(AX# �@��Y|C�ҋ�b|q��ۓ"��c��T0 k� � �&51D"3Q��0 D 3Q ��    ��� �C�XAR(AX# �@��Y|C�ҋ�b�q��ד"��c��T0 k� �  �&51D"3Q��0 D 3Q ��    ��� �C�XAR(AX# �@��Y|C�ҋ�b�q��ד"��c��T0 k� ��" �&51D"3Q��0 D 3Q ��    ��� �C�YAR(AX# �@��Y|C�ҋ�b�q��Ӓ"��c��T0 k� ��$ �&51D"3Q��0 D 3Q ��   ��� �C�YAR(AX# �@��Y|C�ҋ�b�q��Ӓ"ëc��T0 k� ��% �&51D"3Q��0 D 3Q ��    ��� �C�YAR$AX# �@��Y|C�ҋ�b�q��ϒ"ǫc��T0 k� ��) �&51D"3Q��0 D 3Q ��    ��� �C�YAR$AX# �@��Y|C�ҋ�b�q��˒ǫc��T0 k� ��* �&51D"3Q��0 D 3Q ��    ��� �C�YAR$AX# �@��Y|C�⋛b�q��˒˫c��T0 k� ��, �&51D"3Q��0 D 3Q ��   ��� �C�YAR$AX# �@��Y|C�⋛b����˒˫c��T0 k� ��. �&51D"3Q��0 D 3Q ��    ��� �C�YAR$AX# �@��Y|C�⋛b����ǒϫc��T0 k� ��/ �&51D"3Q��0 D 3Q ��    ��� �C�YAR AX# �@��Y|C�⋛b����ǒϫc��T0 k� ��1 �&51D"3Q��0 D 3Q ��    ��� �C�YAR A\# �@��Y|C�⋛b����Òӫc��T0 k� ��2 �&51D"3Q��0 D 3Q ��    ��� �C�YAR A\# �@��Y|C�⋛b����Ò
�ӫc��T0 k� ��4 �&51D"3Q��0 D 3Q ��    ��� �C�YAR A\$ �@��Y|C�⋛b����Ò
�׫c��T0 k� ��6 �&51D"3Q��0 D 3Q ��    ��� �C�YAR A\$ �@��Y|C�⋛b������
�׫c��T0 k� ��7 �&51D"3Q��0 D 3Q ��    ��� �C�YAR A\$ �@��Y|C�⋛R������
�۫c��T0 k� ��9 �&51D"3Q��0 D 3Q ��    ��� �C�YAR A\$ �@��Y|C�⋛R�����
�߫c��T0 k� ��; �&51D"3Q��0 D 3Q ��    ��� �C�YAR A\$ �@��Y|C�⋛R������߫c��T0 k� ��< �&51D"3Q��0 D 3Q ��    ��� �C�YARA\$ �@��Y|C�⋛R�������c��T0 k� ��> �&51D"3Q��0 D 3Q ��    ��� �C�YARA\$ �@��Y|C�⋜R�������c��T0 k� ��@ �&51D"3Q��0 D 3Q ��    ��� �C�YARA\$ �@��Y|C�⋜R�������c��T0 k� ��A �&51D"3Q��0 D 3Q
 ��    ��� �C�YARA\$ �@��Y|C�⋜��������c��T0 k� ��C �&51D"3Q��0 D 3Q	 ��    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��D �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��F �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��H �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��I �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��K �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��M �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��N �&51D"3Q��0 D 3Q  ��    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��P �&51D"3Q��0 D 3Q  ,�    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��R �&51D"3Q��0 D 3Q  ��    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��S �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\$ �@��Y|C�⋜��������c��T0 k� ��U �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\% �@��Y|C�⋜��������c��T0 k� ��V �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\% �@��Y|C�⋜��
�������c��T0 k� ��X �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\% �@��Y|C�⋜��	������ߪc��T0 k� ��Z �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\% �@��Y|C�⋜��������ߪc��T0 k� ��[ �&51D"3Q��0 D 3Q ��   ��� �C�ZARA\% �@��Y|C�⋜��������۪c��T0 k� ��] �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\% �@��Y|C�⋜��������۪c��T0 k� ��_ �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\% �@��Y|C�⋜�������תc��T0 k� ��` �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\% �@��Y|C�⋜�������Ӫc��T0 k� ��b �&51D"3Q��0 D 3Q ��    ��� �C�ZARA\% �@��Y|C�⋜�������Ӫc��T0 k� ��c �&51D"3Q��0 D 3Q ��    ��� �C�ZARA`% �@��Y|C�⋜�������Ϫc��T0 k� ��e �&51D"3Q��0 D 3Q ��    ��� �C�ZARA`% �@��Y|C�⋜��������˪c��T0 k� ��g �&51D"3Q��0 D 3Q ��    ��� �C�ZARA`% �@��Y|C�⋝��������Ǫc��T0 k� ��h �&51D"3Q��0 D 3Q ��    ��� �C�ZARA`% �@��Y|C�⋝��������êc��T0 k� ��j �&51D"3Q��0 D 3Q ��   ��� �C�ZARA`% �@��Y|C�⋝����������c��T0 k� ��l �&51D"3Q��0 D 3Q ��    ��� �C�ZARA`% �@��Y|C�⋝����������c��T0 k� ��m �&51D"3Q��0 D 3Q ��    ��� �C�ZARA`% �@��Y|C�ҋ�����������c��T0 k� ��o �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�ҋ����q������c��T0 k� ��p �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�ҋ����q������c��T0 k� ��r �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�ҋ����q������c��T0 k� ��t �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�ҋ����q������c��T0 k� ��u �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�҇����q������c��T0 k� ��w �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�B�����q������c��T0 k� ��y �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�B�����������c��T0 k� ��z �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�B����������c��T0 k� ��| �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�B����������c��T0 k� ��} �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�B����������c��T0 k� �� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�B����������c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`% �@��Y|C�B����������c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C�B�����������c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C�B�����������c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C�B�����������c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C�B�����������c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C�B�����������c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C�R�����������"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C�R�����������"���T0 k� ��� �&51D"3Q��0 D 3Q ��   ��� �C�[ARA`& �@��Y|C�R�����������"���T0 k� ��� �&51D"3Q��0 D 3Q ��   ��� �C�[ARA`& �@��Y|C�R�����������"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C�R���������R��"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C�R������#���R��"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C� �������#���R��"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C� �������'���R��"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C� �������+���R��"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C� �������/���R��"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C� �������3���R��"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C���	ҋ��7���R��c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C���	ҋ��;���R��c��T0 k� ��� �&51D"3Q��0 D 3Q  ��    ��� �C�[ARA`& �@��Y|C��	ҋ��?���R��c��T0 k� ��� �&51D"3Q��0 D 3Q  -�    ��� �C�[ARA`& �@��Y|C��	ҋ��C���R��c��T0 k� ��� �&51D"3Q��0 D 3Q  ��    ��� �C�[ARA`& �@��Y|C��	ҋ��G��R��c��T0 k� ��� �&51D"3Q��0 D 3Q  ��    ��� �C�[ARA`& �@��Y|C��	ҋ��G��R��c��T0 k� ��� �&51D"3Q��0 D 3Q  ��    ��� �C�[ARA`& �@��Y|C��	⋻�K����c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C��	⋺�O����c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�[ARA`& �@��Y|C��	⋺BS����c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�\ARA`& �@��Y|C��	⋹BW����c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�\ARA`& �@��Y|C��	⋹B[����c��T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�\ARA`& �@��Y|C��	ҋ�B[����"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�\ARAd& �@��Y|C��	ҋ�B_�{���"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� �C�\ARAd& �@��Y|C��	ҋ�Bc�{���"���T0 k� ��� �&51D"3Q��0 D 3Q ��    ��� ����B���E���p(E���Y|C��,� �/��h:^s�3��T0 k� ����&51D"3Q��0 D 3Q ��    ��� ����B���E���x(E���Y|C��4 ��7��p9^s�3��T0 k� ����&51D"3Q��0 D 3Q ��    ��� ����B���E����(E��Y|C��?���?��x9^s�3��T0 k� ����&51D"3Q��0 D 3Q ��    ��� ����B���E��܈(E��Y|C��G���G�р9^w�3��T0 k� ����&51D"3Q��0 D 3Q ��    ��� ����B���E��܌(E��Y|C��O�� �O�ш9^w�3��T0 k� ����&51D"3Q��0 D 3Q ��    ��� ����B��E��ܔ(E��Y|C��W��(�[�ѐ8^w�3��T0 k� �����&51D"3Q��0 D 3Q ��    ��� ����B��E��ܜ(E��Y|C��_��4�c�ќ8^w�3��T0 k� ������&51D"3Q��0 D 3Q ��    ��� ����B��E��ܤ(E��Y|C��g��<�k��8^w�3��T0 k� ������&51D"3Q��0 D 3Q ��    ��� ����B�'�E��ܬ(E��Y|C��o��D�s��7^{�3��T0 k� ������&51D"3Q��0 D 3Q ��    ��� ����B�/�E��	ܴ(E�#�Y|C��w��L�{��7^{�3��T0 k� ������&51D"3Q��0 D 3Q ��    ��� ����B�;�E��ܸ'E�'�Y|C���T����6^{�3��T0 k� ������&51D"3Q��0 D 3Q ��    ��� ���B�C�E����'E�+�Y|C����\�����6^{�3��T0 k� ������&51D"3Q��0 D 3Q ��    ��� ���B�O�E����'E�3�Y|C����d���5^{�3��T0 k� ������&51D"3Q��0 D 3Q ��    ��� ���B�W�E����&E�7�Y|C����p���5^�3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ���B�_�E����&E�;�Y|C����x����4^�3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ��#�B�k�E����&E�C�Y|C���������4^�3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ��+�B�s�E�� ��%E�G�Y|C���������3^�3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ��/�B��E�����%E�O�Y|C���������3^�3��T0 k� ������&51D"3Q��0 D 3Q  /�    ��� ��7�B���E����$E�S�Y|C��������� 2^�3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ��?�B���E����$E�[�Y|C���������2^��3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ��C�B���E���#E�_�Y|C���������1^��3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ��K�B���E���#E�g�Y|C����������0^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��O�B���E���"E�k�Y|C������ ���� 0^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��W�B���E���!E�s�Y|C������  ���(/^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��[�B���E���$!E�w�Y|C������! ���0.^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��_�E���E���, E�{�Y|C������!�r8.^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��c�E���E���4E���Y|C������"�r@-^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��k�E���C���DCM��Y|C�����#�rP+^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��o�E���C���LCM��Y|C�����##�rX*^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��s�E���C���TCM��Y|C���� $+�r`)^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��w�E��C���\CM��Y|C����$3�rh)^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��{�E��C���dCM��Y|C����%;�rl(^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ���E� C���lCM��Y|C��'��%C�rt'^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ���E�  C���tCM��Y|C��/�  &K�r|%^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �Ӄ�E�( E���|CM��Y|C��7� ('S���$^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �Ӄ�E�4 E��}�CM��Y|C��;� 0'[���#^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� Ӈ�E�H E��}�CM��Y|C��K� @)o���!^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �Ӌ�E�P E��}�CM��Y|C��S� H)w��� ^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �S��E"X E��}�C]��Y|C��[� P*���^��3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �S��E"g�E��}�C]��Y|C��_� X+���%���3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �S��E"o�E����C]��Y|C��g� `+����%���3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �S��E"{�E����C]��Y|C��o� h,����%���3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �S��E"��E����C]��Y|C��w� p-����%���3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �C��E"��E����E-��Y|C���x-����%���3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �C��E"��A���E-��Y|C�����/����%���3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �C��E"��A���
E-��Y|C�����/����%���3��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �C��E���A���	E-��Y|C�����0����%���3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ����E���A���E-��Y|C�����1����%���3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ����E���A���E.�Y|C�����1�����%���3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ����E���E����E.�Y|C�����2�����%���3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ����E���E����E.�Y|C�����3�����%���3��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �C��E���E���E�Y|C�����4����	%���3��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C��E���E��� E#�Y|C������5���	�	%���3��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C��E���F ���E'�Y|C������5��	�%���3��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C��E��F ���#�E/�Y|C������6��	�%���3��T0 k� ���#�&51D"3Q��0 D 3Q  ��    ��� �C��E��F ���'�E3�Y|C������7��	�$%���3��T0 k� �+��/�&51D"3Q��0 D 3Q  ��    ��� �C�E��F ���/�E;�Y|C������7��	�(%���3��T0 k� �'��+�&51D"3Q��0 D 3Q  ��    ��� �C�E��F ���7�EC�Y|C������8�#�
0%���3��T0 k� �'��+�&51D"3Q��0 D 3Q  ��    ��� �3{�E�/�@���G�B�O�Y|C����9�3�
0%���3��T0 k� �/��3�&51D"3Q��0 D 3Q  ��    ��� �3x E�7�@���K�B�W�Y|C����:�;�
0%���3��T0 k� �3��7�&51D"3Q��0 D 3Q  ��    ��� �3|E�?�@���S�B�_�Y|C����;�?�
0%���3��T0 k� �7��;�&51D"3Q��0 D 3Q  ��    ��� �3|E�G�@���S�B�g�Y|C����$<�G�	�0%���3��T0 k� �;��?�&51D"3Q��0 D 3Q  ��    ��� �3�E�O�@���W�B�o�Y|C��'��,<�O�	�4%���c��T0 k� �C��G�&51D"3Q��0 D 3Q  ��    ��� �ÀE�W�@���[�B�w�Y|C��3��4=�S�	�4%���c��T0 k� �K��O�&51D"3Q��0 D 3Q  ��    ��� �ÄE�_�@���_�B�{�Y|C��;��<>�W�	�8%���c��T0 k� �S��W�&51D"3Q��0 D 3Q  ��    ��� �ÄE�o�@���g�B���Y|C��K��L@�c�
8%���c��T0 k� �_��c�&51D"3Q��0 D 3Q  ��    ��� �È	E�s�B����k�B���Y|C��S��T@�k�
<%���c��T0 k� �g��k�&51D"3Q��0 D 3Q  ��    ��� �ÈE�{�B����o�B���Y|C��[��\A�o�
@%���c��T0 k� �k��o�&51D"3Q��0 D 3Q  ��    ��� ���EÃ�B����s�B���Y|C��c��dB�s�
@%���c��T0 k� �o��s�&51D"3Q��0 D 3Q  ��    ��� ���EÇ�B����s�B���Y|C��o��lC�w�
D%���c��T0 k� �s��w�&51D"3Q��0 D 3Q  ��    ��� ���EÏ�B���w�B���Y|C��w��tD�{��D%���c��T0 k� �{���&51D"3Q��0 D 3Q  ��    ��� ���EÓ�B���{�B���Y|C����|E���H%���c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ���EÛ�B����B���Y|C���F҃��L%���c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �3�Eã�B�����B���Y|C���Hҋ��P %���c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �3�Eç�B�����B���a�C����Hҋ��W�%���c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �3�Eï�B�����B���a�C����Iҏ��[�%���c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �3�Eó�B�����B���a�C����Jғ��_�%���c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �3�E÷�B�����B���a�C����Kғ��_�%���c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �3�Eû�B�#����B���a�C�ý�LҔ�c�%���c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�Eÿ�B�+����B���a�C�˽�MҔ�g�%���c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�!Eÿ�B�/����B��a�C�ӽ�NҔ�k�%���c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�$E���B�7����B��a�C���PҘ�s�%������T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �C�&E���B�?����B��a�C���QҘ�w�%������T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �	S�'E���B�C����B�#�a�C����R�s{�%������T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �	S�)E���E�K����B�+�Y|C����S�
s�%������T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �	S�*E�ϿE�O����B�3�Y|C���T�s��%������T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �	S�-E�ӼE�[����B�?�Y|C��	2V�s��%������T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �	c�.E�ӺE�c����B�G�Y|C���	2W2�s��%������T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �	c�0E�׸E�g����B�O�Y|C��'�	2X2�s��%������T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �	c�1E�׶E�o����B�W�Y|C��/�	2X2�s��%������T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �	c�2E�׵E�w����B�_�Y|C��7�	2Y2�s��%�����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �	c�3E�׳E�{����B�g�Y|C��?�	B Z2����%�����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �3�5E�ױE������B�o�Y|C�	G�	B(Z2����%�����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �3�6E�װDы����B�w�Y|C�	O�	B,[����%�����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �3�9E�ӭDї����B߇�a�C�	[�	B8\����%�����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �3�:E�ӫDџ����Bߋ�a�C�	c�	2<\�s��%�����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �3�;E�ӪDѧ����Bߓ�a�C�	"k�	2@]�s��%�����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �3�=E�өDѫ����Bߛ�a�C�	"s�	2D]�s��_����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� 3�?E�ϧDѳ����B���a�C�	"w�	2H]�s��_����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� 3�@E�ϦDѻ����B���a�C�	"�	2L^�s��_����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�CA�ˤD������B���a�C����	BT^�s��_����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�EA�ˣD������B���a�C����	BX^�s��%�����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�GA�ǢD������B���a�C����	BX_��s��%�#����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�HA�ǡD������B���Y|C����	B\_�|c��%�#����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�JA�àD������B���Y|C����	B`_�|c��%�'����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�ME㿟D������B���Y|C��ÿ	2d_�xc��%�+����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�OE㻞D������B���Y|C��˿	2h_�tc��%�/����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�QE㷝D�����B���Y|C��ӿ	2h_�tc��%�3����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�SE㳝D�����B���Y|C��߿	2l_�tc��%�3����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�UE㳜D�����B��Y|C���	2l_�pc��%�7����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� #�VE�D�����B��Y|C����	Bp_�pc��%�7����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �XE�D�'����B��Y|C����	Bp_�lc��%�;����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �\E�D�7����B�'�Y|C���	Bt_�lc��%�?����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �]E�D�?����B�/�Y|C���	Bt_�hc��%�C����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �_E�D�C����B�7�Y|C���	2t_�h	���%�G����T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �aE�D�K���B�?�Y|C��#�	2x_�d	���%�G����T0 k� ����&51D"3Q��0 D 3Q  �� 	   ��� �cE�D�S���B�G�Y|C��+�	2x_�d	�Ͼ%�K����T0 k� ����&51D"3Q��0 D 3Q  �� 	   ��� �dE�D�[���B�O�Y|C��3�	2x_�d	�ϼ%�K����T0 k� ����&51D"3Q��0 D 3Q  �� 	   ��� �fEs��D�c���B�W�Y|C��;�	2x_�`	�ϻ%�O����T0 k� ����&51D"3Q��0 D 3Q  �� 	   ��� �gEs��D�k���B�_�Y|C��C�	Bx_�`	�Ϲ%�O����T0 k� ����&51D"3Q��0 D 3Q  �� 	   ��� �iEs��D�s���B�g�Y|C��K�	Bx_�`	�ϸ%�S����T0 k� ����&51D"3Q��0 D 3Q  �� 	   ��� �jEs��D�{���B�o�Y|C��S�	Bx_�\	�˵%�W����T0 k� ����&51D"3Q��0 D 3Q  �� 	   ��� ��mEs��D����B��Y|C��g�	Bx_�\		�ñ%�[����T0 k� ����&51D"3Q��0 D 3Q  �� 	   ��� ��oEc��E����B���Y|C��o� bx_�X	ÿ�%�[����T0 k� �����&51D"3Q��0 D 3Q  �� 	   ��� ��pEc�E����B���Y|C�w� bx_�X#��%�_����T0 k� �o��s�&51D"3Q��0 D 3Q  �� 	   ��� ��qEc{�E����B���Y|C�� bx_�X#��%�_����T0 k� �c��g�&51D"3Q��0 D 3Q  �� 	   ��� ��rEc{�E����B���Y|C��� bx_�T#��%�c����T0 k� �[��_�&51D"3Q��0 D 3Q  �� 	   ��� ���tEcw�E����B���Y|C��� bx_�T#��%�c����T0 k� �S��W�&51D"3Q��0 D 3Q  �� 	   ��� ���uA�o�I���#�BЫ�Y|C��� x_�P#��%�g����T0 k� �G��K�&51D"3Q��0 D 3Q  �� 
   ��� ���vA�k�I���#�Bг�Y|C���� x_�P c��%�g�c��T0 k� �?��C�&51D"3Q��0 D 3Q  �� 
   ��� ���wA�c�I���'�Bл�Y|C���� x_�S�c��%�k�c��T0 k� �7��;�&51D"3Q��0 D 3Q  �� 
   ��� ���xA�_�I����'�B�úY|C���� x_�O�c��%�k�c��T0 k� �3��7�&51D"3Q��0 D 3Q  �� 
   ��� �t xA�W�I�� �+�B�˹Y|C���� x_�O�c��%�o�c��T0 k� �+��/�&51D"3Q��0 D 3Q  �� 
   ��� �tyE�S�J� �+�B�ӹY|C���� x_�O�c��%�o�c��T0 k� �7��;�&51D"3Q��0 D 3Q  �� 
   ��� �tzE�K�J��+�B�۹Y|C���� x_�K�c��%�o�c��T0 k� �;��?�&51D"3Q��0 D 3Q  �� 
   ��� �tyE�G�J��/�B��Y|C���� x_�K�c��%�s�c��T0 k� �?��C�&51D"3Q��0 D 3Q  �� 
   ��� �txE�C�J��/�B��Y|C���� x_K�c��%�s�c��T0 k� �?��C�&51D"3Q��0 D 3Q  �� 
   ��� ��xE�;�J��3�B��Y|C���� x_K�c��%�w�c��T0 k� �?��C�&51D"3Q��0 D 3Q  ��    ��� ��wH�7�I���3�B���Y|C���� x_K�c��%�w�c��T0 k� �3��7�&51D"3Q��0 D 3Q  ��    ��� ��vH�3�I���7�B��Y|C����Bx_G�c��%�{�c��T0 k� �#��'�&51D"3Q��0 D 3Q  ��    ��� ��uH�+�I���7�B��Y|C����Bx_G�c��%�{�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� ��tH�'�I���7�B��Y|C����Bx_G�c��%�{�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� ��sH�#�I���;�B��Y|C���Bx_G�c��%��c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �� rH��J��;�B�#�Y|C���Bx_G�c��_�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� ��$qHs�J��?�B�+�Y|C���Bx_G�c��_�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� ��$pHs�J��?�B�3�Y|C���Bx_G�c��_��c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �t(oHs�J��C�B�;�Y|C��#�Bx_�K�c��_��c��T0 k� ����&51D"3Q��0 D 3Q  �    ��� �t(nHs�J �?�B�C�Y|C��#�Bx_�K�c��_�c��T0 k� ����&51D"3Q��0 D 3Q  ��   ��� �t,mHs�I��?�IG�Y|C��'�Bx_�K�c��_�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �t,kHb��I��?�IO�Y|C��+�Bx_�K�c��_{�c��T0 k� ����&51D"3Q��0 D 3Q  ��    ��� �t0jHb��I�?�IW�Y|C��+�Bx_�O�c��_{�c��T0 k� �߿��&51D"3Q��0 D 3Q  ��    ��� �t4iHb��I�?�I_�Y|C��/��x_�O�c��_{�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �t4gHb�I�;�Ic�Y|C��/��x_�S�c��_w�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �t8fHb�J;�Ik�Y|C��3��x_�S�c��_w�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �t8eHR�J;�I!o�Y|C��3��x_�W�c��_w�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �t<cHR�J/;�I!w�Y|C��3��x_�[�c��_s�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �d<bHR�J/;�I!{�Y|C��7��x_�[�c��_s�c��T0 k� ������&51D"3Q��0 D 3Q  ��    ��� �d<`HR߳J/7�I!��Y|C��7��x_�_�c�_s�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �d@^HR۳I�/7�I!��Y|C��7��x_�c�S�_o�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �d@]Hb״I�/7�I��Y|C��7��x_�g�S�_o�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �d@[HbӴI�/7�I��Y|C��7��x_�g�S{�_o�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �dDZHbϵI�/7�I��Y|C��7��x_�k�S{�_o�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �dDXHb˶I�?7�I��Y|C��7��x_�o�S{�_k�c��T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �dDWHbǶ@?3�I��Y|C��3��x_�s�Cw�_k�"���T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �dDUHr÷@?3�E��Y|C��3��x_�w�Cw�_k�"���T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �dDSHr÷@?3�E��Y|C��3��x_�{�Cs�_g�"���T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �dDRHr��@?3�E��Y|C��/��x_���Cs�_g�"���T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �dDPHr��@?3�E��Y|C��/��x_���Co�_g�"���T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �TDNHr��@?3�E��Y|C��+��x_���Ck�_g�"���T0 k� �����&51D"3Q��0 D 3Q  �    ��� �TDMH���@?3�E�öY|C��+��x_���3k�_c�"���T0 k� �����&51D"3Q��0 D 3Q  ��    ��� �T@KH���@?/�E�˶Y|C��'��x_���3g�_c�"���T0 k� �����&51D"3Q��0 D 3Q ��    ��� �T@IH���@?/�E�϶Y|C��#��x_���3g�_c�"���T0 k� �����&51D"3Q��0 D 3Q ��    ��� �T@HH���@?/�E�׷Y|C����x_���3c�__�"���T0 k� �����&51D"3Q��0 D 3Q ��    ��� �T<FH���@?/�E�۷Y|C����x_���3_�__�"���T0 k� �����&51D"3Q��0 D 3Q ��    ��� �T<EBB��@c?/�E��Y|C����x_����[�__�c��T0 k� ҇����&51D"3Q��0 D 3Q ��    ��� �T8CBB��@c?/�E��Y|C����x_����[�_[�c��T0 k� ҃����&51D"3Q��0 D 3Q ��    ��� �T8BBB��@c?/�E��Y|C����x_����W�_[�c��T0 k� �����&51D"3Q��0 D 3Q ��    ��� �T4@BB��@c?+�F��Y|C����x_����S�_W�c��T0 k� �{���&51D"3Q��0 D 3Q ��    ��� �T4?BB��@c?+�F��Y|C����x_����O�OW�c��T0 k� �{���&51D"3Q��0 D 3Q ��    ��� �D0>BB��@c?+�F�Y|C���x_����K�OS�c��T0 k� �w��{�&51D"3Q��0 D 3Q ��    ��� �D,<BB��@c?+�F�Y|C����x_����G�OS�c��T0 k� �s��w�&51D"3Q��0 D 3Q ��   ��� �D(:BB��@c?+�F�Y|C����x_����?�OO�c��T0 k� �o��s�&51D"3Q��0 D 3Q ��    ��� �D$9Dһ�@c?+�F#�Y|C����x_����;�OK�c��T0 k� �k��o�&51D"3Q��0 D 3Q ��    ��� �D 8Dһ�@c?+�F'�Y|C����x_��7�OG�c��T0 k� g��k�&51D"3Q��0 D 3Q ��    ��� �D7Dһ�@c?+�E�/�Y|C����x_£��3�?G�"���T0 k� c��g�&51D"3Q��0 D 3Q ��    ��� �D6Dҿ�@�?'�E�7�Y|C����x_£��/�?C�"���T0 k� _��c�&51D"3Q��0 D 3Q ��    ��� �D5Dҿ�@�?'�E�?�Y|C����x_£��'�??�"���T0 k� _��c�&51D"3Q��0 D 3Q ��    ��� �D4D�ú@�?'�E�G�Y|C����x_§��#�?;�"���T0 k� [��_�&51D"3Q��0 D 3Q ��    ��� �D3D�ǻ@�?'�E�K�Y|C����x_B����?;�"���T0 k� W��[�&51D"3Q��0 D 3Q ��    ��� �                                                                                                                                                                            � � �  �  �  d A�  �K����   �      6 \��f� ]��� � �� \�   $ $      � ��     \> �~H     Q    	                . �          ۰     ���   0	&
          �        � ��'     �G ��    �v�z                  �         &�     ���   0
           &�          ��     &� � �     Z :                 	  �         `      ���   (	          ��Q    \	     ��I�    �����I�          
                �o           @�     ���   H
$
         ��o�         / �}m    ��m� �}m                        ��o           �p     ���   0
3           ���� ��	      C���    �������                             ���E              \  ���    P		 5             ���-        W ��n    ���	 ��n    ��                  6	�� �          R0     ��@    		�          ���l  � �	    k �bS    ���� �c�    �\��                	�� �          P�   	  ��@  (
	          ����  4 4     �w�    ��{� ���    ��               '�� ��        ��     ��@   8	 

         ���5   u      ����J    ���"����    ���S             	 �� �         	 \�     ��H   H


         ���a  � �  	   � �f�    ��9� �<    �I�               8	�� �         
 ��     ��`   0
3
         ��b� **      � ��    ��b� ��                            ���s               ��@   		 5 	                 ��      �                                                                           �                               ��        ���          ��                                                                 �                          ��� ��        ��h�� �' ��<�h�� �0F   �                 x                j  ^  �	   �                                �        ���         ��                                                               �                          � � ��� �� � � ��� � ����h��        	   
      
  [   i �� s��J       �d �m` �d n` ��  n� �� n� �D 0w` �� @w� �D 0x@ ��  n� �� n� ڄ �w` ۤ x� �� x����J ����X � �D _  �d  _@ Hd _� H� _� ;� q  �� t� �� �u  �� v  
�\ W� 
� W� 
�\ X  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }����� ����� � �� _` � �c` � d` �� h` � �h� �$ i� $ �m` $ n` D  n� �� �`� �� a� �D `j� � 0k� �d 0l  �� l` � �o� � p� ��  }����� � 
�\ W  
�\ W� 
�< W� 
�| X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���� � �����d  ������  
�fD
��L���"����D"� �  " `   J jF��    "�j "���
��
���     �j��  
  �
� �  �  
� ����  ��     ���  �        ��     � �      ����  ��     ���          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �      �� �T ���        � �T ��        �        ��        �        ��        � 	 	 4�    ������        ��                         T�) , ��� �                                      �                 ����	            	���� 	���&��  �� � 2               13 Teemu Selanne       3:30                                                                        5  5     �C
� � �J�> J�> �c � � c� � �c� � � c� � �cW � �	c_ � �
ck � � s � �ct � � cv � �c� � � c� � �K/ �KY �KI �c� �c� �c�' i	�# i	�: y�! y�L"�: "�L"�6*�E |"; � � "F � �  "B � � !"Q � � "" � #"F �<  " {L  "! {L  "! {  "F � �(" � �)!� {  "F � +"K �L  "! {L  "+ {<  " {� /"� �{0� �{1
� � � 2"D �  "I � � 4"D �  "I � � 6"P � � 7"' �  "L �  "L � � :" � ;"F �<  " {<  " { � >"Q �  "G �@� 
�( 
�! 
�                                                                                                                                                                                         �� P        �     @ 
        �     U P E _  ��        	            ������������������������������������� ���������	�
���������                                                                                          ��    �rh�� ��������������������������������������������������������   �4, 0   * l� ���� � ��@	��@ւ��A�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          0    (    �� �D�J     O�  	                           ������������������������������������������������������                                                                        	                                                                     ������                                             ��������������������������������� ������������������������������ � �� ������ ������ ��� ����������������� ������������������� ���� ������� �  ��������������� ����������� ������� ����� ������������ ������������������ ����������                             	        G    0      �  �\�J      �                             ������������������������������������������������������                                                                                                                                         ����  �  �                                           �������������������� �������������� ���������������� ������� ���� ������� ����������� ������������� ����������� ����������� ���������������� ������ ���������������  ������������� ��������������������� ������������� ����� ��� ����                                                                                                                                                                                                                                           
          	                                                                       �              


             �  }�         ���%      #%����  8�����  �����������������������������������������������������������������������������      .�      6�     O     O                                                      ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � %�d �\        0                                                                                                                                                                                                                                                                 )n)n1n  	�Y                a      a      b                  c      c                                                                                                                                                                                                                                                                                                                                                                                                                  > �  >�  J�  0  �  Jc�  ���������|��(����� ��˶�A�˖�r�˖������H                      ��        $   �   & QW  �  g                  �                                                                                                                                                                                                                                                                                                                                      0 K K   �                       !��                                                                                                                                                                                                                            Z   �� �� Ѱ��      �� f      ��������������������������������� ������������������������������ � �� ������ ������ ��� ����������������� ������������������� ���� ������� �  ��������������� ����������� ������� ����� ������������ ������������������ ������������������������������ �������������� ���������������� ������� ���� ������� ����������� ������������� ����������� ����������� ���������������� ������ ���������������  ������������� ��������������������� ������������� ����� ��� ����             $����������������˪�������������������������������������f��ff��ff�������̺�ff�fffffffffffffffffff����ƹ��ffʻfff�fffjffffffffffff��������������������ʺ��l���f˪������������������������������������������������������������������fff�fff�fff�ffk�ffi�ff��ff��ff�ffffffff�fff�x�����w��xx�������wfffffff�ffff�fffww��ww�x����wx��fk��ff��ff��ffʹffj��fʪ�f�ˊ�k������������ʚ��������������������������������������������˫��ʫ��ff��fl��fl��ff̫fff�ffʬ�f���f�����������wu���w��l������f����W��������xww��Wy�l����x������k���W�fi���j���j���f����˘�����y�y�y����������������������������������������������������ʻ����ʫɚ�����l���ƨ�lƘ�j���k���̜i���j���kxx���wx������wx������������ƈx����������������wW����w�������������������������z����������˫��̺������������������������������������������������������������ʺ������k������������������������������������������x�j���˙�x�˘��̩�x������x���xx�x������x������wx���˫��ʫ����������˪�����ʻ��������������������������������������ʻ�ʻ�����ʪ̫����˺��������������������˪�����f���k��f��fǶW�g���k���̻���f������������������x�������˩f̺�����uw�����w��x�wXx��˪�����������l����l���i��ƹx�f�������������������ʫUW��UUU�UUUX      7      D   �C �                       \     �  ���������J'      ��     b�   �         �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ��  � ��     � ��   	 ��   p �� �� ��    ����  ��  �| >�������J J���|����  ��  �|  ��  �1   ��   ��  � ��   � �� �� �z   � � �$ ��   T ��  �� ��   ��  �� �� �  �� �� �z � ��� �$  � �  �� �  �      �  ��   y���� e�����  g���  �     f ^�         �� ���      y      ��f����2�������J��f����      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                                                  U  T   T   T     T UDUDDUDDDDDDDDDDDDDDDP   E�  DU� DDU�DDDUDDDDDDDDDDDD                UP  E�  E   E                                           ���U�UTD�DDDDDDTDD TDD   �   U_ DEU�DDDUDDDDD��DZT�DDDDDDDDDDDDTDDDDDDDDUTU�����DDDDDDDDDDDEDDDEDDDDTUTU�Ԫ���Z_   P   � �U�UTDUDDDDUTD�DT��D        U_��DEU_DDD_DDDPDDE�DDE  �DD DD DD �DD �UD  �U       DZTDEDDDDE�DDE�DDE�TDDT�DE�TE���DDTU�ZD���������DDTDD��ZT�T���ZTDDE��D��T�T��DUTTT��Z��TQTDDUTD�DDDTDDD�DDDDDDE�DD_TDE�DD_ DDP DDP DD_ DU_ U�  �                                       TE�DDD�UUU                    ���DDDUUUTD  D  D  D  D  U��D�TDDDDEUUDP  DP  DP  DP  UP  TDE�DDDPUUU_                                                    wwwwtDDDt""$t"""t"w"t"w"t"w"t""$wwwwtDGtD"GtD"GtD"GtD"GtD"GtD"GtwwwwDDDD"D"""D"""DD""Gt""Gt""Gt"wwwwDDDD"B"""B""DDD"GwD"GwB$GtB$wwwwDwww$www$wwt$wwtGwwtGwwwwwwwwwwwtDDDD�DLL�D���D�D�D�t�D�t�D�wwwwDDww��Gw��Gww�Gww�Gww�Gww�Gwt"""t"w"t"w"t"w"t"""t""$tDDDwwwwD"GtD"GtD"GtD"DDD""$D""$DDDDwwww"Gt""Gt""Gt""Gt""Gt""Gt"DGtDwwwwGt"DGD"DGB$GGB$DGB""GB""GDDDwwwwwwwwwwwwwwwwDwww$www$wwwDwwwwwwwt�D�t�D�t�D�t�D�t�D�t�DMtDDDwwwww�Gww�Gww�Gww�Gw��Gw��GwDDwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 " ""   "" !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  "!  " ! " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                            " ""   "" !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                             �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   �   " � ��      �    �   �   �"  ""  !� �� ��  �               �   " ��.�  ��   ����   �       �                                   �    ��"  �"                    ".  ".  ��� ���                                                                                                                                                                                             	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��   ��  �    �  �  ��                 �   �   �"  �.  .   �                 �                        ��"� �"� ����                              �   �      ��   �  ��  �  �  �         � ".��".��/����  �                                                                                                                                                      �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp��& ��vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �" �"" �"   �                    .   .   �   ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                            �".��".  ���    �                    �   O   T     ��                                 � "�"  �    � � �                                                                                                                                                           ̙ �ɪ���˭�̻� �� �   ""  ""  .         �� ̻ �� ��w �rb �wg���z�����ٙ�����ˍ�ݙ8����DD��3D��33L�3� �3+ ��" �" ""  ".  �  �   �                        �T  �U  �D  +�� ��� 
�  �"" �"" ��"/��� ��� �  ��               �   �   �   �   �   �   �@      �    �  �   �""��""����    �   "    �  /   /   �   �                       �                        ��"� �"� ����                                     	�  ���� �                               ""  "".  . �    �                                                                                                                                        �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �               0   0   �   �" �""��        "   "   "   �   �               �   " ��.�  ��                   �                        ��"� �"� ����                            �   ���                                                                                                                                                                                                            �  �  �  �  w  �  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �       �   �                   �           �   �                     �     �                                      � ����ݼ� ����                                                                                                                                                                               �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp��& ��vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �" �"" �"   �                    .   .   �     .  " "" ��� "                                                                �               �     "   "                                 ���                                                                                                                                                                                        �   �   w   b   g     
�  �� �� �� �̻ ������ɨ�-�ݼ-ݍ�"Չ� X���DDX�TCZES3�T3�@ ��"��"�� ""� �"/��/��        �   ��  ��  ��  {�  wp  ��� ���������̻��̽��̽���ؚ��ڨ��؛˻��˸� ��  �C  D0  3   0   0   �   �   �    �  /   ���                     2�  2   1   �                  �    � .� .  �� 	  
  �  ",  ""  �"   "                      �"  �"  �� "            � "�",�"+� ",                       "  .���"    �     �                                       �   ���                            �   "                                                                                                                   � ̻ �ۼͺ�	ۚ����C�˽T;��UJ��ET�35J�D3T�  ̰ ̻	�̻���w���&��wv��wpʨ� ��� ��� ��  "�� .� "�� ��0 "          .  .  "   "             �  �� ʝ ,��+� "" "��CEJ�D5J� J�  �� 
�� �  �� �+� �"" """����    �                   � ˹ Y�����
�ڛ��٩ �� �̽���ݪ۽w�}�&��vv���p���              �                             ���                         �"  �"                    ���.�                     P   P   P   P   U   E   ��  �ɠ ��� ���  �"  " ��"�""��"! � �  �   �   �   �                                                                                                                     �  �� 
����ݜ��ש˙��ܻ��ݼ��ۼ �"+ ". B"( �"# JUC ZTD 
TC 
�D 
�D JD@ �T 
�@ �� � "��"/��""��"� �  �    �    �   ̰  ��  ��  �z� wy� w�� �̸ �۪��ة��
��� �����3>��33 33 33  �� �� 
�  "" "" ��"/����  �  �                           �   �   "   �"  ""� " �                        � ���             �  "� "  "  "  �                         �                      �".��".  ���    �       �  �  �  �                                      "  "  "           �  � �                       � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                           �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��  .�"." "."   /�  �  �              � ��         �� �� �� g} &' vw                     ".  ".  ���                                                                                                                                                                                                     �  �  � 	� 
� ɭ �� 蘰 ��� ��������  ��  �   �      �  �   �   �             ��  �ͻ�������ڛ��z���z��ڊ���� 3���34ۍ�5��������ݘ ��������������������� �������� ��"/�".� .�  �                       �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� ���                         �� ��                  �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                   2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ DD D@                     �� ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD l � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=GwDGwqwDDwtwwww3333DDDD  � �!�aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( """"����������A��I��I X � �!�aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx""""�����A�DA�I��I� w � �!�aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""��������I���I���I���I��� � � �!�aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(MAMAMMMM�M�M����3333DDDD  � �!�aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�D�����MD��M����3333DDDD m � �!�a�a� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� Sa��m(`���4���4���4���4���4���43334DDDD � � �!�aa � � � �!i!j � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� Sa��(M""""wwwwqqqqwGwGGG � � �!�aa � � � �!m!n � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� Sa�� 
(�""""wwwwwwqqDAwG � u!�!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� S)��(-(�������������������333DDD!�!�!�!�!�!� �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5M��M��D��M����������3333DDDD + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+DD��D�M��D����3333DDDD � W  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ������ ���((W(�""""������DH�H� � a � l � � � � � �������� � �� � � � � � ���	����� � � �� �������l(�(a(�""""�������H�H��D �  � y � � � � � � � � � � � � � � � �� ��������� � � � � � � � � ������y(�(�""""��������H��H��H��H� = l �  � � � � � � � � � � ��� � � � � �������� � � � ��� � � � ������((�l(=DD������L��DL����3333DDDD    �  � � � � � � � � � ������ � � � � � ���� � � � ������ � � �����((�(( L�A�AAD��DL�����3333DDDD x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���4���4���4L��4L��4���43334DDDD w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww""""���������M�MMM  � w w � � � � � � � � � ��	� � � ��� � � � � � � � � � � ��	� � � ��� �����ww�(""""�������A��AA �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((���������������333DDD ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`I��I����������������3333DDDD M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M��A���I��I���I�����3333DDDD � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(�""""������������������������ � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(�""""������D�D��� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5""""������������������������ x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�xwqwwqwwwwwqwwwDwwww3333DDDD w � � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxwwqqwwwDDwtGwwww3333DDDD � � � i i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+www4www4www4www4www4www43334DDDD W � � u u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(�""""wwwwwwqwwwqwqwq a � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(�""""wwwwwwwDwGwA  � �!�aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(��A�L�L�L��L���333DDDLDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDDC
� � �J�> J�> �c � � c� � �c� � � c� � �cW � �	c_ � �
ck � � s � �ct � � cv � �c� � � c� � �K/ �KY �KI �c� �c� �c�' i	�# i	�: y�! y�L"�: "�L"�6*�E |"; � � "F � �  "B � � !"Q � � "" � #"F �<  " {L  "! {L  "! {  "F � �(" � �)!� {  "F � +"K �L  "! {L  "+ {<  " {� /"� �{0� �{1
� � � 2"D �  "I � � 4"D �  "I � � 6"P � � 7"' �  "L �  "L � � :" � ;"F �<  " {<  " { � >"Q �  "G �@� 
�( 
�! 
�3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD��������������������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ��������������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ��������������������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE��������������������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD��������������������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD��������������������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD��������������������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� ����7�\�J��<�V�I�P�[�H�P�S�S�L�������8�>�7���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� ��!��-�V�I��0�Z�Z�L�U�Z�H����������8�>�7���""""������A�D��I��""""�������D����� ����>�L�L�T�\��=�L�S�H�U�U�L��������>��<���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �8�>�7���!���A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �>��<�����""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,��,��,�D�,���#333DDDDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II�""""������D""""������IADD���I""""��������D��""""�������I��I�I�I�""""�������A�D�II�I""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            