GST@�                                                            \     �                                               �   �                        ����e ��	 ʳ������������������        i      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    "�j* ,  �����
�"     �j@ �    ��
  �                                                                               ����������������������������������      ��    bb QQb  114 44c c   c      		 

       	   
       ��G �   ( (                 nhp ))1         888�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                ��  �       ��   @  #   }   �                          �                                                     'w w  )n)h1p  �    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��D>hEE�?����	�+�|3����E.|F������3�T0 k� ������SXD"!U2d    ��    ����B��D>`FE�;����	�'�|3����E.|F������3�T0 k� ������SXD"!U2d    ��    ����A��D>XGE�7����	�#�|3����E.|F������3�T0 k� ������SXD"!U2d    ��    ����@�D>PHE�3����	��|7����E.�F������3�T0 k� ������SXD"!U2d    ��    ����?�D>HHE�+����	��|7����E.�F��� ���3�T0 k� ������SXD"!U2d    �8    ����>�D>4JE��	��	��|;����E.�G�� ���3�T0 k� �o��s�SXD"!U2d   ��?    ����=�DN,KE��	��	��|;����E��G�� ���x3�T0 k� �c��g�SXD"!U2d   ��?    ����< �DN$LE��	��	��|?�Λ�E��G�� ��p3�T0 k� �S��W�SXD"!U2d   ��?    ����; �DNME��	��^�|?�Λ�E��G�� ۿ�d3�T0 k� �G��K�SXD"!U2d   ��?    ����: �DNNE��	��^�|?�Λ�E��G� Ӿ�\3�T0 k� �7��;�SXD"!U2d   ��?    ����9 �DNNE��	��^�|C�Λ�E��G-{� ˽�T3�T0 k� �+��/�SXD"!U2d   ��?    ����8 �I�OE������^�|C�Η�E��G-w� ý�L3�T0 k� ���#�SXD"!U2d   ��?    ����8��I� PE������^�|C�ޗ�E��G-s� ���D3�T0 k� ����SXD"!U2d   ��?    ����8��I��QE������]��|G�ޓ�E��
G-k� ���43�T0 k� ������SXD"!U2d   ��? 	   ����8��I��QE������]��|G�ޏ�E��	G-g����,3�T0 k� ������SXD"!U2d   ��? 	   ����8��I��RE������]��|G�ޏ�E��G-c����$3�T0 k� ������SXD"!U2d   ��? 	   ����8��I��RE������]��|K�E��G-[����3�T0 k� ������SXD"!U2d   ��? 	   ����8��I��SE���������|K�EΘG-W����3�T0 k� ������SXD"!U2d   ��? 	   ����8���I��SE���������|K�EΘG-S����3�T0 k� ������SXD"!U2d   ��? 	   ����8���I��SE���������|K�EΘG-O��� 3�T0 k� ������SXD"!U2d   ��? 	   ����8���I��SE���������|K���EΘG-K�P{���3�T0 k� ������SXD"!U2d   ��? 	   ����8���I��TE��������|G��w�EΜ G-C�Pk���3�T0 k� �{���SXD"!U2d   �? 	   ����8���I��TE��������|D �s�EΟ�G-?�Pc� �3�T0 k� <{���SXD"!U2d   ��? 	   ����8���I��TE��������|D �o�EΟ�G-?�P[� �3�T0 k� <{���SXD"!U2d   ��? 	   ����8���I͸TE��������|D�k�EΟ�G-C�PS� �3�T0 k� <{���SXD"!U2d   ��? 	   ����8���IʹTE��������|D�g�EΟ�G-C�PK� �3�T0 k� <{���SXD"!U2d   ��? 	   ����8���IͰTE�������|@�c�EΟ�G-C�PG� �3�T0 k� <{���SXD"!U2d   ��? 	   ����8���IͬTE�������|@�[�Eޟ�G-C�P?�P�3�T0 k� �{���SXD"!U2d   ��? 	   ����8���IͨTE��������|@�W�Eޟ�E�G�P7�P�3�T0 k� �{���SXD"!U2d   ��? 	   ����8���E�TE��������|@�S�Eޟ�E�G�P/�P�3�T0 k� �{���SXD"!U2d   ��? 	   ����8���E�TE�{������|@�O�Eޟ�E�G�@'�P�3�T0 k� �{���SXD"!U2d   ��? 	   ����8���E�UE�o�����|@�C�Eޛ�E�G�@�P�3�T0 k� ,{���SXD"!U2d   ��? 	   ����8���E�UE�k�����|@�;�Eޛ�E�K�@�P�3�T0 k� ,{���SXD"!U2d   ��?    ����8���E�UFg�����|@�7�Eޗ�E�K�@�@x3�T0 k� ,{���SXD"!U2d   ��?    ����8���E�UF_�����|@�/�Eޗ�E�G�O��@p3�T0 k� ,{���SXD"!U2d   ��?    ����8���E��VF[�����|@�+�Eޓ�E�G�O��@h3�T0 k� ,{���SXD"!U2d   ��?    ����8���E��VFW��݇�|@�#�Eޓ�E�G�O�@`3�T0 k� L{���SXD"!U2d   �?    ����8���E��WFS��݇�|@�E��TC�O�@X3�T0 k� L{���SXD"!U2d   ��?    ����8���E�|XD�G����|<�E��TC��ۯ@H3�T0 k� L{���SXD"!U2d    ��?    ����8��E�xXD�C����|<�E��TC��ӯ@@3�T0 k� L{���SXD"!U2d    ��?    ����8��E�tYD�C��]�|<��E��TC��˯@43�T0 k� ,{���SXD"!U2d    ��?    ����8��E�tZD�?��]�|<��E��TC��ï@,3�T0 k� ,{���SXD"!U2d    .�?    ����8��E�pZD�;��]{�|<��D>�TC�����$3�T0 k� ,{���SXD"!U2d    ��?    ����8��E�l[D�;��]w�|<��D>{�T-?�����3�T0 k� ,{���SXD"!U2d    ��?    ����8��E�h\D�;��]w�|<��D>w�T-;�����3�T0 k� ,{���SXD"!U2d    ��?    ����8��E�d]D�7��]s�|<��D>s�T-;�����3�T0 k� �{���SXD"!U2d    ��?    ����8��E�`^D�7���]o�|<��D>o�T-7�����3�T0 k� �{���SXD"!U2d    ��?    ����8�߲F\`D�3���]k�|<��D>g�T-3������3�T0 k� �{���SXD"!U2d   ��?    ����8�۴FXaD�3���]g�|<��D>c�T-/������3�T0 k� �{���SXD"!U2d   ��?    ����8�׶FXbD�3� l��]g�|<��D>_�T=/�����3�T0 k� �{���SXD"!U2d   ��?    ����8�ӷFTcD�3� l��]g�|<��D>[�T=/��w���3�T0 k� �{���SXD"!U2d   ��?   ����8�ϹFPdD�3� l��]g�|<��D>W�T=/��o���3�T0 k� ,{���SXD"!U2d   �?    ����8�˺FPfD�3� l��c�|<]��D>S�T=+��g���3�T0 k� ,{���SXD"!U2d    ��?    ����8�˼FPgD�3� l��_�|8]��DNO�T=+��_���3�T0 k� ,{���SXD"!U2d    ��?    ����8�ǾFLhD�3���[�|8]��DNK�T=+��W���3�T0 k� ,{���SXD"!U2d    ��?    ����8�ÿFLiD�3���W�|8]��DNG�T=+��O���3�T0 k� ,{���SXD"!U2d    ��?    ����8���E�LjD�3���O�|8]��DNC�T=+��G���3�T0 k� �{���SXD"!U2d    ��?    ����8���E�LlD�3���O�|8	]��DN;�T=+��?���3�T0 k� �{���SXD"!U2d    ��?    ����8���E�HmD�7���O�|8	]��DN7�T=+��7���3�T0 k� �{���SXD"!U2d    ��?   ����8γ�E�HnD�7� ��K��8	]��DN3�T=+��/���3�T0 k� �{���SXD"!U2d    ��?    ����8Ϋ�E�HoD�7� ��-G��8	]��DN/�T='��+���3�T0 k� �{���SXD"!U2d    ��?    ����8Σ�E�HqD�7� ��-?��8]{�DN#�T='����t3�T0 k� �{���SXD"!U2d    ��?    ����8Ο�E�LrD�7� ��-?��8]w�DN�T='����l3�T0 k� �{���SXD"!U2d    ��?    ����8Λ�E�LtD�7�L��-;��8]o�D^�T=#����d3�T0 k� �{���SXD"!U2d    ��?    ����8Η�E�LuD�7�L��-7��8]o�D^�T=�O��\3�T0 k� �{���SXD"!U2d    ��?    ����8Ώ�E�PvD�7�L��-7��8]o�D^�T=�N���T3�T0 k� �{���SXD"!U2d    ��?    ����8΋�E�PwD�7�L��=3��8]o�D^�T=�N��L3�T0 k� �{���SXD"!U2d    ��?    ����8΃�E�TxE7�|��=/��8]o�D]��T=�N��<3�T0 k� �{���SXD"!U2d    ��?    ����8�{�E�TyE7�|��=+��8]k�D]��T=�N߹�43�T0 k� �{���SXD"!U2d    ��?    ����8�w�B�XzE7�|��='��8]k�D]��T=�N׺�,"��T0 k� �{���SXD"!U2d    ��?    ����8�s�B�X{E7�|��='��8]k�D]��T=�NϺ� "��T0 k� �{���SXD"!U2d    ��?    ����8�o�B�\{E7�|��=#��8 ]k�D]��T=�Nǻ�"��T0 k� �{���SXD"!U2d    ��?    ����8�g�B�`|E7����=��;�]g�D]��T=�>ü�"��T0 k� �{���SXD"!U2d    ��?    ����8�c�B�`|E7����=��;�]g�Dm��T=�>���"��T0 k� �{���SXD"!U2d    ��?    ����8�W�E�h}E7����=��7�]g�Dm��T<��>����"��T0 k� �{���SXD"!U2d    ��?    ����8�O�E�h~E7����=��7�Mg�Dm��T<��>����"��T0 k� �{���SXD"!U2d    ��/    ����8�K�E�l~E}7����=��7�Mc�Dm��T<��>���� "��T0 k� �{���SXD"!U2d    ��/    ����8�G�E�p~E}7����=��7�Mc�Dm��T<��>����!"��T0 k� �{���SXD"!U2d    ��/    ����8�?�E�tE}7����=��7�Mc�Dm��T<��>��N�""��T0 k� �{���SXD"!U2d    ��/    ����8�7�E�xE}7����=��7�M_�Dm��T<��>��N�"3�T0 k� �{���SXD"!U2d    ��/    ����8�3�E�xE}7����=��3��_�Dm��T<��>��N�#3�T0 k� �{���SXD"!U2d    ��/    ����8�'�E��Em7����=��3��[�Dm��T<��Nw�N�%3�T0 k� �{���SXD"!U2d    ��/    ����8��E��Em7����=��3��[�D=��T<��Ns�N�&3�T0 k� �{���SXD"!U2d    ��/    ����8��CM�Em7���=��3��W�D=��T<��Nk�N�'3�T0 k� �{���SXD"!U2d    ��/    ����8��CM�~Em3���<���3��W�D=��T<��Ng�N�(3�T0 k� �{���SXD"!U2d    ��/    ����8��CM�~Em3���<���3��S�D={�T<��N_�N�(3�T0 k� �{���SXD"!U2d    ��/    ����8��CM�~Em3���<���3��O�D=s�T<��>[�N�)3�T0 k� �{���SXD"!U2d    ��/    ����8���CM�}E]/���<���3��K�D=c�T<��>O�N�+3�T0 k� �{���SXD"!U2d    ��/    ����8���CM�}E]/���<���/��G�E�_�T<��>K�>|,"s�T0 k� �{���SXD"!U2d    ��/    ����8���CM�|E]/���<���/��C�E�W�T<��>C�>t-"s�T0 k� �{���SXD"!U2d    ��/    ����8���CM�{E]+���<���/��?�E�O�T<��>?�>l."s�T0 k� �{���SXD"!U2d    ��/    ����8�� CM�{E]+���<���/��?�E�G�T<��>7�>h0"s�T0 k� �{���SXD"!U2d    ��/    ����8��C]�zE�'���<���/��;�E�C�T<��>3�>`1"s�T0 k� �{���SXD"!U2d    ��/    ����8��C]�yE�#���<���/��7�E�;�T<��>/�>X2"s�T0 k� �{���SXD"!U2d    ��/    ����8�C]�xE����<���/��/�E�+�T<��.#�>L4"s�T0 k� �{���SXD"!U2d    ��/    ����8�C]�wE����<���/��+�E�'�T<��.�>D6"s�T0 k� �{���SXD"!U2d    ��/    ����8�E��vE����<���/��'�E�T<��.�><7"s�T0 k� �{���SXD"!U2d    ��/    ����8�E��uE����<���/��#�E�T<��.�>89"s�T0 k� �{���SXD"!U2d    ��/    ����8�E��tD=���<���+���E�T<��.�>0:3�T0 k� �{���SXD"!U2d    ��/    ����8�E��sD=�L�<���+���E�T<��.�.,<3�T0 k� �{���SXD"!U2d    ��/    ����8��E��rD=�L�<���+���E� T<��.�.$=3�T0 k� �{���SXD"!U2d    ��/    ����8��	EͼpD=�L�<���+���E��T<��.�. ?3�T0 k� �{���SXD"!U2d    ��/    ����8�x
EͼnE��L�<���+���E��	T<��.�.B3�T0 k� �{���SXD"!U2d    ��/    ����8�p
E��mE�� �<���'���E��
T<��-��.C3�T0 k� �{���SXD"!U2d    ��/    ����8�h
E��lE�� �<���'���E��T<��-��.E3�T0 k� �{���SXD"!U2d    ��/    ����8�d
E��jE�� �<���'���E��T<����.F3�T0 k� �{���SXD"!U2d    ��/    ����8�\E��iE�� �<���'���D��T<����. H3�T0 k� �{���SXD"!U2d    ��/    ����8�TE��hE��� �<���'���D��T<����-�J3�T0 k� �{���SXD"!U2d    ��/    ����8�HE��eE��� l�<���'�m�D��T<����-�M3�T0 k� �{���SXD"!U2d    ��/    ����8�@E��dE��� l�<���'�m�D��T<�����N3�T0 k� �{���SXD"!U2d    ��/    ����8�<
E��bE��� l�<���'�m�D��T<�����P3�T0 k� �{���SXD"!U2d    ��/   ����8�4
E��aD��� l�<���'�l��D��T<�����R3�T0 k� �{���SXD"!U2d    ��/    ����8�0
E��_D��� l�<���'�l��D��T<�����R3�T0 k� �{���SXD"!U2d    ��/    ����8� 	Eݼ^D��� ��<���'����D��T<�����S3�T0 k� �{���SXD"!U2d    ��/    ����8�	Eݸ^D��� ��<���'����D��T<�����S3�T0 k� �{���SXD"!U2d    ��/    ����8�Eݴ]El�� ��<���'����D��T<���� �S3�T0 k� �{���SXD"!U2d    ��/    ����8�Eݰ]El�� ��<���'����D�� T<�����T3�T0 k� �{���SXD"!U2d    ��/    ����8�Eݨ\El���<���'�l��D��#T<������T3�T0 k� �{���SXD"!U2d    ��/    ����8� Eݠ\El���<���'�l��D��%T<������T3�T0 k� �{���SXD"!U2d    ��/    ����8��Eݜ[El���<���'�l��D�|'T<������T3�T0 k� �{���SXD"!U2d    ��/    ����8��Eݘ[El���<���'�l��E�x(T<������T3�T0 k� �{���SXD"!U2d    ��/    ����8�EݐZEl���<���'�l��E�t*T<������T3�T0 k� �{���SXD"!U2d    ��/    ����8�E�ZEl��|�<���'�l��E�l-T<����
� T3�T0 k� �{���SXD"!U2d    ��/    ����8�E�YEl��|�<���'�l��E�d/T<��� �T3�T0 k� �{���SXD"!U2d    ��/    ����8� E�|YEl��|�<���'�l��E�`1T<��~ �T3�T0 k� �{���SXD"!U2d    ��/    ����8��E�tYEl��|�<���'�l��E�\2T<��~�T3�T0 k� �{���SXD"!U2d    ��/    ����8��E�pYEl��|�<���'�l��E�X4T<��~�T3�T0 k� �{���SXD"!U2d    ��/    ����8��E�dYEl����<���'�l��FP8T<��~�S3�T0 k� �{���SXD"!U2d    ��/    ����8���E�\YEl����<���'�l��FL9T<����S3�T0 k� ������SXD"!U2d    ��&    ����8���E�TYE\���<���'�l��FH;T<����S3�T0 k� ������SXD"!U2d    ��&    ����8���E�PYE\{���<���'�l��FD=T<����R3�T0 k� ������SXD"!U2d    ��&    ����8���E�HYE\s���<���'�l��FD?T<���� R3�T0 k� ������SXD"!U2d    ��&    ����8���E�<YE\g�|�<���#�l��F<BT<����(Q3�T0 k� �����SXD"!U2d    ��&    ����8���E�4ZE\_�|�<���#�\��F8DT<����,P3�T0 k� ������SXD"!U2d    ��&    ����8���E�0ZE\[�|�<���#�\��F8FT<����0P3�T0 k� ������SXD"!U2d    ��&    ����8���E�(ZE\S�|�<���#�\��F4HT<���~4O3�T0 k� ������SXD"!U2d    ��&    ����8���E� [P�K�|�<���#�\��F4JT<���~8O3�T0 k� �����SXD"!U2d    ��&    ����8���E�[P�C��<���#�\��F0LTL���~<N3�T0 k� �����SXD"!U2d    ��&    ����8���E�\P�C��<���#���E�0PTL��� ~DL3�T0 k� �s��w�SXD"!U2d    ��&    ����8���E�]P�?��<������E�,RTL��� �DL3�T0 k� �o��s�SXD"!U2d    ��&    ����8���E�^P�;��<������E�,STL��� �HK3�T0 k� �k��o�SXD"!U2d    ��&    ����8���E� ^P�7�%|�<������E�,UTL���$�LK3�T0 k� �c��g�SXD"!U2d    ��&    ����8���E��`P�7�%|�<�����{�E�,YTL���(�TI3�T0 k� �W��[�SXD"!U2d    ��&    ����8���E��aP�7�%|�<�����w�E�,[TL���(�TI3�T0 k� �S��W�SXD"!U2d    ��&    ����8���F�bP�3�%|�<�����o�E�,\U\���(�XH3�T0 k� �G��K�SXD"!U2d    ��&    ����8���F�cP�3�%|�<�����k�E�,^U\���,�\H3�T0 k� �?��C�SXD"!U2d    ��&   ����8���F�dP�/�%|�<�����c�E�,`U\���,�\H3�T0 k� �7��;�SXD"!U2d    ��&   ����8���F�fP�'�%|�<�����W�E�0cU\���0
�`G3�T0 k� �+��/�SXD"!U2d    ��&    ����8���F�gP�'�%|�<�����O�E�0eU\���0	�dG3�T0 k� �'��+�SXD"!U2d    ��&    ����8���F�hP�#�%|�<�����K�E�0fU\���0�dG3�T0 k� �'��+�SXD"!U2d    ��&    ����8���F�iP��%|�<�����C�E�4hU\���4�dF3�T0 k� ���#�SXD"!U2d    ��&    ����8��F�lP��%|�<�����7�E�8jU\���4�hE3�T0 k� ����SXD"!U2d    ��&    ����8}�F�mE��%|�L�����/�E�8lU\���8�lE3�T0 k� ����SXD"!U2d    ��&    ����8}�F�nE��%|�L�����'�E�<mU\���8�lD3�T0 k� ����SXD"!U2d    ��&    ����8}�E��pE��%|�L������E�<nU\���8�pD3�T0 k� ������SXD"!U2d    ��&   ����8}�E��rE��%|�L������E�@qU\��< �pB3�T0 k� ����SXD"!U2d    ��&    ����8}�E��sE��%|�L������E�DrU\��?��tA3�T0 k� �����SXD"!U2d    ��&    ����8}�E��tE���%|�L������E�HsU\��?��tA3�T0 k� ������SXD"!U2d    ��&   ����8}�E��vE���%|�L�������E�LtU\��C��x@3�T0 k� ������SXD"!U2d    ��&    ����8}�E��wE���%|�L�������E�LtU\��C��x?3�T0 k� ������SXD"!U2d    ��&    ����8�#�E��yE���%|�\������E�TvA���G��|=3�T0 k� �����SXD"!U2d    ��&    ����8�'�B��zE���%|�\������E�TwA���G��|<3�T0 k� �����SXD"!U2d    ��&    ����8�+�B��{E���%|�\�����߯E�XwA���G��|;3�T0 k� ����SXD"!U2d    ��&    ����8�+�B��|E���%|�\�����ۮCL\xA���G���:3�T0 k� ����SXD"!U2d    ��&    ����8�/�B��}E���%|�\�����ӬCL\xA���K���93�T0 k� �ߕ��SXD"!U2d    ��&    ����8�/�B��~E����\�����ϫCL`yA���K���73�T0 k� �۔�ߔSXD"!U2d    ��&    ����8�3�E��E����\����˩CLdyA���K���63�T0 k� �ߔ��SXD"!U2d    ��&    ����8�7�E���E����\����çCLdyA���K���53�T0 k� ����SXD"!U2d    ��&    ����8�;�E���E����������CLlzA���O���23�T0 k� �ۑ�ߑSXD"!U2d    ��&    ����8�;�E���F��L�������CLlzA���O���13�T0 k� �ې�ߐSXD"!U2d    ��&    ����8�?�E��F��L�������CLpzBL��O���03�T0 k� �ې�ߐSXD"!U2d    ��&    ����8}C�E��F��L�������CLpzBL��S�	ތ/3�T0 k� �׎�ێSXD"!U2d    ��&    ����8}C�E��F��L�������C\tzBL��S�	ތ.3�T0 k� �׌�یSXD"!U2d    ��&    ����8}G�E��~F��L�,������C\xzBL��S�	ތ-3�T0 k� �ӊ�׊SXD"!U2d    *�&    ����8}G�E��~P���L�,������C\xzBL��S�	ތ,3�T0 k� �׊�ۊSXD"!U2d    ��&    ����8}K�E��}P���L�,������C\|zBL��W�	ތ+3�T0 k� �Ӊ�׉SXD"!U2d    ��&    ����8}O�E��|P���L�,������C\�y@��W�	�)3�T0 k� �ۈ�߈SXD"!U2d    ��&    ����8}O�E��|P���L�l�������C\�y@��W�	�(3�T0 k� �׋�ۋSXD"!U2d    ��&    ����8}S�E��{P���L��l�������C\�x@��W�	�'3�T0 k� �׎�ێSXD"!U2d    ��&    ����8}S�E��{Q��\��l�������C\�x@��[�	�'3�T0 k� �׏�ۏSXD"!U2d    ��&    ����8}W�E��zQ��\��l�������C\�w@��[�	�&3�T0 k� �א�ېSXD"!U2d    ��&    ����8mW�E��yQ��\��l�������C\�wB���[�	ތ&3�T0 k� �ې�ߐSXD"!U2d    ��&    ����8m[�E��xQ��\��l�����ǔCl�uB���_�	ތ$3�T0 k� ����SXD"!U2d    ��&    ����8m[�E��wQ��\��l�����˓Cl�uB���_�	ތ$3�T0 k� ����SXD"!U2d    ��&    ����8m_�E��vQ��\��l�����ӓCl�tB���_�	ތ#3�T0 k� ����SXD"!U2d    ��&    ����8m_�E��uQ��\��l�����גCl�sD���_�	�#3�T0 k� ����SXD"!U2d    ��&    ����8m_�E��tQ��\��l�����ߒCl�rD���_�	�#3�T0 k� ������SXD"!U2d    ��&    ����8m_�E��sP���\��l������Cl�qD���_�	�"3�T0 k� ������SXD"!U2d    ��&    ����8m_�E��qP���\��l������Cl�pD���c�	�"3�T0 k� ����SXD"!U2d    ��&    ����8m_�E��oP���l��l�������Cl�nD���c�	ތ"3�T0 k� ����SXD"!U2d    ��&    ����8m_�E��nP���l��l�������Cl�mD���c�	ތ!3�T0 k� ����SXD"!U2d    ��&    ����8]_�E� m@��l��l������C|�lD���c�	ތ!3�T0 k� ����SXD"!U2d    ��&    ����8]_�E� k@��l��l������C|�kD���g�	ތ!3�T0 k� �#��'�SXD"!U2d    ��&    ����8]_�E� j@��l��l������C|�jD���g�	ތ!3�T0 k� �+��/�SXD"!U2d    ��&    ����8]_�E�i@��l��l������C|�iD���g�	�!3�T0 k� �/��3�SXD"!U2d    �&    ����8]_�I}g@��l��l������C|�gD���g�	�!3�T0 k� �3��7�SXD"!U2d    ��/    ����8][�I}fE���<��l�����#�C|�fD���g�	�!3�T0 k� �7��;�SXD"!U2d    ��/    ����8][�I}dE���<��������/�C|�cD��	�g�	�!3�T0 k� �?��C�SXD"!U2d    ��/    ����8]W�I}cE���<��������3�C|�bD��	�k���!3�T0 k� �G��K�SXD"!U2d   ��/    ����8]W�EMbE���<��������;�C|�aD��	�k���!3�T0 k� �K��O�SXD"!U2d   ��/    ����8]S�EMaE���<��������?�C|�_D��	�k���!3�T0 k� �O��S�SXD"!U2d   ��/    ����8]S�EM_E���<��������G�CL�^D��	�k���!3�T0 k� �S��W�SXD"!U2d   ��/    ����8]O�EM^E���<��������K�CL�\D��	�k���!3�T0 k� �W��[�SXD"!U2d   ��O    ����8MK�EM]E���<��������S�CL�ZD��	�k���!3�T0 k� �[��_�SXD"!U2d   ��O    ����8MG�E=ZE;��<��������[�CL�WH��	�k���!3�T0 k� �g��k�SXD"!U2d   ��O    ����8MC�E=YE;��<��������c�CL�UH��	�k���!3�T0 k� �k��o�SXD"!U2d   ��O    ����8MCE=XE;��,��<�����g�CL�TH��	�k���!3�T0 k� �o��s�SXD"!U2d    ��O    ����8M?�E=VE;��,��<�����k�CL�RH��	�k���!3�T0 k� �s��w�SXD"!U2d    ��O    ����8M;�E=UE;��,��<�����s�CL�PH��	�k���!3�T0 k� �w��{�SXD"!U2d    ��O    ����8M7�CMSE+��,��<�����w�CL�NH��	�k���!3�T0 k� �{���SXD"!U2d    ��O    ����8M3�CMRE+��,��<�����{�CL�MH��	�k���!3�T0 k� ������SXD"!U2d    ��O    ����8M/�CMNE+��,�������̇�CL�IH��	�k���!3�T0 k� ������SXD"!U2d    /�O    ����8=+�CMME+Ͽ,�����#�̋�C\�GH��	�k���!3�T0 k� ������SXD"!U2d    ��O    ����8='�CMKE+Ͼ,�����#�̏�C\�EH��	�k���!3�T0 k� ������SXD"!U2d    ��D    ����8=#�CMIEӽ,�����#�̓�C\�CBL�	�k���!3�T0 k� ������SXD"!U2d    ��D    ����8=�CMFE׻,�����#�̟�C\�?BL�	�k���!3�T0 k� ������SXD"!U2d    ��D    ����8M�CMDE׺,� ���!��̣�C\�=BL�k���!3�T0 k� ������SXD"!U2d    ��D    ����8M�CMBE۹����!��̧�C\�;BL�k���!3�T0 k� ������SXD"!U2d    ��D    ����8M�C]@E߸�L��!��̫�C\�9D��k���!3�T0 k� ������SXD"!U2d    ��D    ����8M�C]<E��L��!��̳�C\�5D��k���!3�T0 k� ������SXD"!U2d    ��D    ����8=�C]<B�� 	L��|�̷�I\�3D��o���!3�T0 k� ������SXD"!U2d    ��D    ����8=�C]:B�� L��|#�̻�I\�1D��o���!3�T0 k� ������SXD"!U2d    ��D    ����8=�E=8B��\��|#�̿�I\�/O��o�N�!3�T0 k� ������SXD"!U2d    ��D    ����8<��E=4B��\��|#�̿�I\�,O����s�N�!3�T0 k� ������SXD"!U2d    ��D    ����8<��E=2B���\��|#����I\�*O����w�N�!3�T0 k� ������SXD"!U2d    ��D    ����8<��E=0B���\��|#����Il�)O����w�N�!3�T0 k� ������SXD"!U2d    ��D    ����8<��E=,B��|��|#��ÏIl�&O����{�N�!3�T0 k� ������SXD"!U2d    ��D    ����8<��E=*B��� |��|#��ÏIl�$O�����N�!3�T0 k� ������SXD"!U2d    ��D    ����8<��E=*B���$|��|#�,ÐIl�#O������ �!3�T0 k� ������SXD"!U2d    ��D    ����8	\��E=*B���0|��!�#�,ÑI\� O������ �!3�T0 k� ������SXD"!U2d    ��D    ����8	\��@m*B���8��!�#�,ǒI\�O������ �!3�T0 k� ������SXD"!U2d    ��D    ����8	\��@m)B���<��!�#�,ǒI\�O������ �!3�T0 k� ������SXD"!U2d    ��D    ����8	\��@m)B�#��D��!�#�%<ǓI\�O�������� 3�T0 k� ������SXD"!U2d    ��D    ����8	\��@m(B�+��P��##�%<˔Il�O�������� 3�T0 k� ������SXD"!U2d    ��D    ����9	l��E-(E3��X��##�%<˔Il�O�������� 3�T0 k� ������SXD"!U2d    ��D    ����:	l��E-'E7��\��##�%<˕Il�O�������� 3�T0 k� ������SXD"!U2d    ��D    ����;	l��E-&EC��l��##�%<˖Il�O�������� 3�T0 k� ������SXD"!U2d    ��D    ����<	l��E-&EK��p����#�%<ϖI\�O�������� 3�T0 k� ������SXD"!U2d    ��D    ����=	\��E%EO�}x����#�%<ϗI\�O�������� 3�T0 k� ������SXD"!U2d    ��D    ����>	\��E%EW�}�����#�%<ϗI\�O�������� 3�T0 k� ������SXD"!U2d    ��D    ����?	\��E $Ec�}�����#�%<ϘI\�D܏��Ǆ�� 3�T0 k� ������SXD"!U2d    ��D    ����A	\��E$#E�k�}�����#�%<әIl�D܏��τ�� 3�T0 k� ������SXD"!U2d    ��D    ����C	l��B�$#E�o�}�����#�%<әIl�D܏��ӄ�� 3�T0 k� ������SXD"!U2d    ��D    ����E	l��B�("E�w�}�����#�%<ӚIl�Dܓ��ۄ�� 3�T0 k� ������SXD"!U2d    ��D    ����G	l��B�0"E���}�����#�%<ӛIl�Dܓ����� 3�T0 k� �����SXD"!U2d    �D    ����G	l��B�4!E���}� ,���#�%<כCL�Dܗ�	��� 3�T0 k� ����SXD"!U2d    �D    ����G ���@8!E����� ,���#�%<כCL�Dܗ�	��� 3�T0 k� �#��'�SXD"!U2d    ��D    ����G ���@8 BL���� ,���#�%<לCL�Dܗ�	���� 3�T0 k� �3��7�SXD"!U2d    ��D    ����G ���@@ BL���� ,���#�%<۝CL�Dܛ�	���3�T0 k� �C��G�SXD"!U2d    ��D   ����G ���@DBL���� -��#�%<ߝCL�
Dܟ�	���"s�T0 k� �O��S�SXD"!U2d    ��D    ����G ���@DBL���� -��#�%<ߞCL�
D��	/���"s�T0 k� �W��[�SXD"!U2d    ��D    ����G ���@HBL���� -��#�%<�CL�	D��	/���"s�T0 k� �c��g�SXD"!U2d    ��D    ����G ���@LBL���� -��#�%<�CL�D��	/���"s�T0 k� �k��o�SXD"!U2d    ��D    ����G ���@PBL�������#�%<�CL�D��	/���"s�T0 k� �c��g�SXD"!U2d    ��D    ����G ���@PBL�����#��#�%<�CL�D��	/�~�"s�T0 k� �[��_�SXD"!U2d    ��D    ����G ���@TBL�����'��#�%<�CL�M|��	�~�"s�T0 k� �[��_�SXD"!U2d    ��D    ����G ���@XBL�����/��#�%<�C\�M|��	#�~�"s�T0 k� �[��_�SXD"!U2d    ��D   ����G ���@XBL�����7��#�%<�C\�M|��	'�"s�T0 k� �[��_�SXD"!U2d    ��D    ����G ���@\BL�����;��#�%<�C\�M|��	+�"s�T0 k� �_��c�SXD"!U2d    ��D    ����G ���@`BL��� �C��#�%<�C\��M|��	/�"s�T0 k� �c��g�SXD"!U2d    ��D    ����G ���@`BL����K��#�%<��C\��M|��	//�3�T0 k� �g��k�SXD"!U2d    ��D    ����G ���@dBL����O��#�%<��C\��M���	/3�3�T0 k� �k��o�SXD"!U2d    ��D    ����G ���@hBL���
�W��#�%<��C\��M���	/7�3�T0 k� �s��w�SXD"!U2d    ��D    ����G ���@hBL���
 _��#�%<��C\��M���	/7�3�T0 k� ������SXD"!U2d    ��D    ����G ���@lBL���
 g��#�%<��C\��M���	/;�$3�T0 k� ������SXD"!U2d    ��D    ����G ���@lBL���	 k��#�%<��C\��M����;�o(3�T0 k� ������SXD"!U2d    ��D    ����G ���@pBL��� 	 s��#�%<��C\��M����?�o,3�T0 k� ������SXD"!U2d    ��D    ����G ���@tBL���$ w��#�%<��Cl��M����?�o,3�T0 k� ������SXD"!U2d    ��D    ����G ���@tBL���( ��#�%<��Cl��M����C�o03�T0 k� ������SXD"!U2d    ��D    ����G ���@xBL���, ���#�%<��Cl��M����C�o43�T0 k� ������SXD"!U2d    ��D    ����G ���@xBL���0 ���#�%<��Cl��M|���C�o83�T0 k� ������SXD"!U2d    ��D   ����G ���@|BL���4 ���#�%<��Cl��M|���G�o<"��T0 k� ������SXD"!U2d    ��D    ����G ���@|BL���8 ���#�%<��Cl��M|���G�o<"��T0 k� ������SXD"!U2d    ��D    ����G ���@�BL���< ���#�%<��Cl��M|���K�o@"��T0 k� ������SXD"!U2d    ��D    ����G ���@�BL���@ ���#�%<��Cl��M|���K�?@"��T0 k� ������SXD"!U2d    ��D    ����G ���@�BL���D ���#�%<��Cl��M|���O�?D
"��T0 k� ������SXD"!U2d    ��D    ����G ���@�BL���H ���#� l��Cl��M|���O�?D	"��T0 k� ������SXD"!U2d    ��D    ����G ���@�BLÙ�L ���#� l��Cl��M|���S�?H"��T0 k� ������SXD"!U2d    ��D    ����G ���@�BLÙ�P ���#� l��C|��M|���S�?H"��T0 k� �����SXD"!U2d    ��D    ����G ���@�BLÙ�T ���#� l��C|��BL���S�?L"��T0 k� ����SXD"!U2d    ��D    ����G ���@�BLØ�X ���#� l��C|��BL���W�?L"��T0 k� ����SXD"!U2d    ��D    ����G ���@�BLØ�X ���#� l��C|��BL���W�?P"��T0 k� ����SXD"!U2d    ��D    ����G ���@�BLØ�\ ���#� l��C|��BL���[�?P3�T0 k� ����SXD"!U2d    ��D    ����G ���@�BLØ�` ���#� l��C|��BL���[�?P3�T0 k� ����SXD"!U2d    ��D    ����G ���@�BLØ�d ���#� l��C|��BL���[�?T 3�T0 k� ���#�SXD"!U2d    ��D    ����G ���@�BLØ�h ���#� l��C|��BL���_�?W�3�T0 k� �#��'�SXD"!U2d    ��D    ����G ���@�BL×�h ���#� l��C|��BL���_�?[�3�T0 k� �'��+�SXD"!U2d    ��D    ����G ���@�BL×�l ���#� l��C|��BL���_�?[�3�T0 k� �+��/�SXD"!U2d    ��D    ����G ���@�BLǗ�p ���#� l��C|��BL���c�?[�3�T0 k� �/��3�SXD"!U2d    ��D    ����G ���@�BLǗ�t  ���#� l��CL��BL���c�?_�3�T0 k� �7��;�SXD"!U2d    ��D    ����G ���@�BLǗ�t  ���#� l��CM�BL���g�?_�3�T0 k� �;��?�SXD"!U2d    ��D    ����G ���@�BLǗ�x  ���#� l��CM�BL���g�Oc�3�T0 k� �?��C�SXD"!U2d    ��D    ����G ���@�BLǗ�� ���#� ��CM�BL���g�Oc�3�T0 k� �C��G�SXD"!U2d    ��D    ����G ���@�BLǖ��� ���#� ��CM�BL���k�Oc�3�T0 k� �G��K�SXD"!U2d    ��D    ����G ���@�BLǖ��� ��#� ��CM�BL���k�Og�3�T0 k� �K��O�SXD"!U2d    ��D    ����G ���@�BLǖ��� ��#� ��CM�BL���k�Og�3�T0 k� �O��S�SXD"!U2d    ��D    ����G ���@�BL˖��� ��#� ��CM�BL���o�Og�3�T0 k� �S��W�SXD"!U2d    ��D    ����G ���@�BL˖��� ��#� ��CM�BL���o�Ok�3�T0 k� �W��[�SXD"!U2d    ��D    ����G ���@�BL˖��� ��#� ��CM�BL���o�Ok�3�T0 k� �[��_�SXD"!U2d    ��D    ����G ���@�BL˖��� ��#����CM�BL���o�Ok�3�T0 k� �_��c�SXD"!U2d    ��D    ����G ���@�BL˕��� ��#����CM�BL���s�Oo�3�T0 k� �c��g�SXD"!U2d    ��D    ����G ���@�BL˕��� ��#����C]�BL���s�Oo�3�T0 k� �g��k�SXD"!U2d    ��D    ����G ���@�BL˕��� #��#����C]�BL���s�Oo�3�T0 k� �k��o�SXD"!U2d    ��D    ����G ���@�BL˕��� #��#����C]�BL���w�Os�3�T0 k� �o��s�SXD"!U2d    ��D    ����G ���@�BLϕ��� '��#����C]�BL���w�Os�3�T0 k� �s��w�SXD"!U2d    ��D    ����G ���@�BLϕ��� +��#����C]�BL���w�Os�3�T0 k� �w��{�SXD"!U2d    ��D    ����G ���@�BLϕ��� /��#����C]�BL���w�Os�3�T0 k� �w��{�SXD"!U2d    ��D    ����G ���@�BLϕ��� 3��#����K��BL���{�Ow�3�T0 k� �{���SXD"!U2d    ��D    ����G ��@�BLϕ��� 7��#����K��BL���{�Ow�3�T0 k� �����SXD"!U2d    ��D    ����G ��@�BLϔ��� ;��#����K��BL���{�Ow�3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLϔ��� ;��#����K��BL���{�O{�3�T0 k� ������SXD"!U2d    ��D   ����G ��@�BLϔ��� ?��#����K��BL����O{�3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLϔ��� C��#����K��BL����O{�3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLϔ��� G��#����K��BL����O{�3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӔ��� G��#����K�#�BL����O�3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӔ��� K��#����K�#�BL�����O�3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӔ��� O��#����K�#�BL�����O�3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӔ��� S��#����K�'�BL�����O�3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӓ��� S��#����K�'�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӓ��� W��#����K�+�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӓ��� [��#����K�+�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӓ��� [��#����K�+�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӓ��� _��#����K�/�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӓ��� c��#����K�/�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLӓ��� c��#����K�/�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLד��� g��#����K�/�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLד��� k��#����K�3�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLד��� k��#����K�3�BL�����O��3�T0 k� ������SXD"!U2d    ��D   ����G ��@�BLד��� o��#����K�3�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLד��� s��#����K�7�BL�����O��3�T0 k� ������SXD"!U2d    ��D    ����G ��@�BLג��� s��#����K�7�BL�����O��3�T0 k� ����óSXD"!U2d    ��D   ����G ��@�BLג��� w��#����K�7�BL�����O��3�T0 k� ����òSXD"!U2d    ��D   ����G ��@�BLג��� w��#����K�;�BL�����?��3�T0 k� �ò�ǲSXD"!U2d    ��D    ����G ��@�BLג��� {��#����K�;�BL�����?��3�T0 k� �ò�ǲSXD"!U2d    ��D    ����G ��@�BLג��� {��#����K�;�BL�����?��3�T0 k� �ǲ�˲SXD"!U2d    ��D    ����G ��@�BLג��� ��#����K�;�BL�����?��3�T0 k� �˲�ϲSXD"!U2d    ��D    ����G ��@�BLג��� ��#����K�?�BL�����?��3�T0 k� �˱�ϱSXD"!U2d    ��D    ����G ��@�BLג��� ���#����K�?�BL�����?��3�T0 k� �ϱ�ӱSXD"!U2d    ��D    ����G ��@�BLے��� ���#����K�?�BL�����?��3�T0 k� �ϱ�ӱSXD"!U2d    ��D    ����G ��@�BLے��� ���#����K�?�BL�����?��3�T0 k� �ӱ�ױSXD"!U2d    ��D    ����G ��@�BLے��� ���#����K�C�BL�����?��3�T0 k� �ӱ�ױSXD"!U2d    ��D    ����G ��@�BLے��� ���#����K�C�BL�����?��3�T0 k� �ױ�۱SXD"!U2d    ��D    ����G �߰@�BLے��� ���#����K�C�BL�����?��3�T0 k� �װ�۰SXD"!U2d    ��D    ����G �߰@�BLے��� ���#����K�C�BL�����o��3�T0 k� �۰�߰SXD"!U2d    ��D    ����G �߰@�BLے��� ���#����K�G�BL�����o��3�T0 k� �۰�߰SXD"!U2d    ��D    ����G �߰@�BLے��� ���#����K�G�BL�����o��3�T0 k� �߰��SXD"!U2d    ��D    ����G �߯@�BLۑ��� ���#����K�G�BL�����o��3�T0 k� �߰��SXD"!U2d    ��D    ����G �߯@�BLۑ��� ���#����K�G�BL�����o��3�T0 k� ����SXD"!U2d    ��D    ����G �߯@�BLۑ��� ���#����K�K�BL�����_��3�T0 k� ����SXD"!U2d    ��D    ����G �ۯ@�BLۑ��� ���#����K�K�BL�����_��3�T0 k� ����SXD"!U2d    ��D    ����G �ۮ@�BLۑ��� ���#����K�K�BL�����_��3�T0 k� ����SXD"!U2d    ��D    ����G �ۮ@�BLۑ��� ���#����K�K�BL�����_��3�T0 k� ����SXD"!U2d    ��D    ����G �ۮ@�BLۑ��� ���#����K�K�BL�����_��3�T0 k� ����SXD"!U2d    ��D    ����G �ۮ@�BLߑ��� ���#����K�O�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �ۮ@�BLߑ��� ���#���K�O�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �ۭ@�BLߑ��� ���#���K�O�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �׭@�BLߑ��� ���#���K�O�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �׭@�BLߑ��� ���#���K�O�BL������{�3�T0 k� �����SXD"!U2d    ��D    ����G �׭@�BLߑ��� ���#���K�S�BL������w�3�T0 k� �����SXD"!U2d    ��D    ����G �׭@�BLߑ��� ���#���K�S�BL������s�3�T0 k� ������SXD"!U2d    ��D    ����G �׬@�BLߑ��� ���#���K�S�BL������o�3�T0 k� ������SXD"!U2d    ��D    ����G �׬@�BLߑ��� ���#���K�S�BL������k�3�T0 k� ������SXD"!U2d    ��D    ����G �׬@�BLߑ��� ���#���K�S�BL������g�3�T0 k� ������SXD"!U2d    ��D    ����G �Ӭ@�BLߑ��� ���#� �K�S�BL������c�3�T0 k� ������SXD"!U2d    ��D    ����G �Ӭ@�BLߑ��� ���#� �K�W�BL������_�3�T0 k� ������SXD"!U2d    ��D    ����G �Ӭ@�BLߑ��� ���#� �K�W�BL������[�3�T0 k� �����SXD"!U2d    ��D    ����G �ӫ@�BLߐ��� ���#� �K�W�BL������W�3�T0 k� �����SXD"!U2d    ��D    ����G �ӫ@�BLߐ��� ���#� �K�W�BL������S�3�T0 k� �����SXD"!U2d    ��D    ����G �ӫ@�BLߐ��� ���#� �CMW�BL������O�3�T0 k� ����SXD"!U2d    ��D    ����G �ӫ@�BLߐ��� ���#� �CMW�BL������K�3�T0 k� ����SXD"!U2d    ��D    ����G �ӫ@�BLߐ��� ���#� �CM[�BL������C�3�T0 k� ����SXD"!U2d    ��D    ����G �ӫ@�BLߐ��� ���#� �CM[�BL������?�3�T0 k� ����SXD"!U2d    ��D    ����G �ϫ@�BLߐ�� ���#� �CM[�BL������;�3�T0 k� ����SXD"!U2d    ��D    ����G �Ϫ@�BLߐ�� ���#� �CM[�BL�����3�3�T0 k� ����SXD"!U2d    ��D    ����G �Ϫ@�BL��� ���#� �CM[�BL�����/�3�T0 k� ����SXD"!U2d    ��D    ����G �Ϫ@�BL��� ���#� �CM[�BL�����+�3�T0 k� ����SXD"!U2d    ��D    ����G �Ϫ@�BL��� ���#� �E�_�BL�����#�3�T0 k� ����SXD"!U2d    ��D    ����G �Ϫ@�
BL��� ð�#� �E�_�BL������3�T0 k� ����SXD"!U2d    ��D   ����G �Ϫ@�
BL��� ð�#� �E�_�BL������3�T0 k� ����SXD"!U2d    ��D    ����G �Ϫ@�
BL��� ð�#� �E�_�BL������3�T0 k� ����SXD"!U2d    ��D   ����G �ϩ@�
BL��� ǰ�#� �E�_�BL������3�T0 k� ����SXD"!U2d    ��D    ����G �ϩ@�
BL��� ǰ�#� �E�_�BL������3�T0 k� ����SXD"!U2d    ��D    ����G �ϩ@�
BL��� ǰ�#� �E�_�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �˩@�
BL��� ǰ�#� �E�_�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �˩@�
BL��� ˰�#� �E�_�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �˩@�
BL��� ˯�#� �E�_�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �˩@�
BL��� ˯�#� �E�_�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �˩@�
BL��� ˯�#� �E�_�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �˨@�
BL��� ϯ�#� �E�_�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �˨@�
BL��� ϯ�#� �E�_�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �˨@�
BL��� ϯ�#� �E�[�BL�������3�T0 k� ����SXD"!U2d    ��D    ����G �˨@�
BL��� ӯ�#� �E�[�BL�� o����3�T0 k� ����SXD"!U2d    ��D    ����G �˨@�
BL��� ӯ�#� �E�[�BL�� o����3�T0 k� ���#�SXD"!U2d    ��D    ����G �˨@�
BL��� ӯ�#� �E�W�BL�� o����3�T0 k� ���#�SXD"!U2d    ��D    ����G �˨@�
BL��� ӯ�#� �E�W�BL�� o��3�T0 k� ���#�SXD"!U2d    ��D    ����G �Ǩ@�
BL��� ӯ�#� �E�S�M|�� o��3�T0 k� ���#�SXD"!U2d    ��D    ����G �Ǩ@�
BL��� ׯ�#� �E�S�M|�� ���3�T0 k� �#��'�SXD"!U2d    ��D    ����G �ǧ@�
BL��� ׮�#� �E�O�M|�� ���3�T0 k� �#��'�SXD"!U2d    ��D    ����G �ǧ@�
BL��� ׮�#� �E�O�M|�� ����{�3�T0 k� �#��'�SXD"!U2d    ��D    ����G �ǧ@�
BL��� ׮�#� �E�K�M|�� ����s�3�T0 k� �#��'�SXD"!U2d    ��D    ����G �ǧ@�
BL��� ׮�#� �E�G�M|�� ����k�3�T0 k� �#��'�SXD"!U2d    ��D    ����G �ǧ@�
BL��� ۮ�#� �E�C�M|�����_�3�T0 k� �'��+�SXD"!U2d    ��D    ����G �ǧ@�
BL��� ۮ�#� �E�C�M|�����W�3�T0 k� �'��+�SXD"!U2d    ��D    ����G �ǧ@�
BL��� ۮ�#� �E�?�M|�����O�3�T0 k� �'��+�SXD"!U2d    ��D    ����G �ǧ@�
BL��� ۮ�#� �E�;�M|�����G�3�T0 k� �'��+�SXD"!U2d    ��D    ����G �ǧ@�	BL��� ۮ�#� �E�7�M������?�3�T0 k� �'��+�SXD"!U2d    ��D    ����G �ǧ@�	BL��� ߮�#� �E�3�M������7�3�T0 k� �+��/�SXD"!U2d    ��D    ����G �ǧ@�	BL��� ߮�#� �E�/�M���_���/�3�T0 k� �+��/�SXD"!U2d    ��D    ����G �Ǧ@�	BL��� ߮�#� �E�+�M���_���'�3�T0 k� �+��/�SXD"!U2d    ��D    ����G �Ǧ@�	BL��� ߮�#� �E�'�M���_����3�T0 k� �+��/�SXD"!U2d    ��D    ����G �Ǧ@�	BL��� ߮�#� �E�#�M���_����3�T0 k� �+��/�SXD"!U2d    ��D    ����G �Ǧ@�	BL��� ߮�#� �E��M���_����3�T0 k� �+��/�SXD"!U2d    ��D    ����G �æ@�	BL��� ��#� �E��M�����3�T0 k� �/��3�SXD"!U2d    ��D    ����G �æ@�	BL��� ��#� �E��M������3�T0 k� �/��3�SXD"!U2d    ��D    ����G �æ@�	BL��� ��#� �E��M|����3�T0 k� �/��3�SXD"!U2d    ��D    ����G �æ@�	BL��� ��#� �D��M|����3�T0 k� �/��3�SXD"!U2d    ��D    ����G �æ@�	BL��� ��#� �D��M|���߸3�T0 k� �/��3�SXD"!U2d    ��D    ����G �æ@�	BL��� ��#� �D��M|���׸3�T0 k� �/��3�SXD"!U2d    ��D    ����G �æ@�	BL��� ��#� �D��M|�����ϸ3�T0 k� �3��7�SXD"!U2d    ��D    ����G �æ@�	BLߑ�� ��#� �D��M|����=Ƿ3�T0 k� �3��7�SXD"!U2d    ��D    ����G �æ@�	BLߑ�� ��#� �D��M|����=��3�T0 k� �3��7�SXD"!U2d    ��D    ����G �æ@�	BLߑ�� ��#� �D��M|���=��3�T0 k� �3��7�SXD"!U2d    ��D    ����G �å@�	BLے�� ��#� �D��M|���=��3�T0 k� �3��7�SXD"!U2d    ��D    ����G �å@�	BLے�� ��#� �D��BL��{�=��3�T0 k� �3��7�SXD"!U2d    ��D    ����G �å@�	BLے�� ��#� �D��BL��{�=��3�T0 k� �3��7�SXD"!U2d    ��D    ����G �å@�	BLד�� ��#� �D��BL��w�=��3�T0 k� �7��;�SXD"!U2d    ��D    ����G �å@�	BLד�� ��#� �D��BL��w�=��3�T0 k� �7��;�SXD"!U2d    ��D    ����G �å@�	BLӔ�#� ��#� �D��BL��s�=��3�T0 k� �7��;�SXD"!U2d    ��D    ����G �å@�	BLӔ�#� ��#� �D��BL��s�=��3�T0 k� �7��;�SXD"!U2d    ��D    ����G �å@�	BLӔ�#� ��#� �D��BL��o�={�3�T0 k� �7��;�SXD"!U2d    ��D    ����G �å@�	BLϕ�#� ��#� �D��BL��o�=w�3�T0 k� �7��;�SXD"!U2d    ��D    ����G �å@ 	BLϕ�#� ��#� �D��BL��o�=o�3�T0 k� �7��;�SXD"!U2d    ��D    ����G �å@ 	BL˕�#� ��#� �D��BL��/k�=g�3�T0 k� �;��?�SXD"!U2d    ��D    ����G �å@ 	BL˕�#� ��#� �D��BL��/k�M_�3�T0 k� �;��?�SXD"!U2d    ��D    ����G �å@ 	BL˕�#� ��#� �D��BL��/g�M[�3�T0 k� �;��?�SXD"!U2d    ��D    ����G ���@ 	BL˕�#� ��#� �D��BL��/g�MS�3�T0 k� �;��?�SXD"!U2d    ��D    ����G ���@ 	BLǕ�#� ��#� �D��BL��/g�MO�3�T0 k� �;��?�SXD"!U2d    ��D    ����G ���@ 	BLǕ�#� ��#� �D��BL��/c�MG�3�T0 k� �;��?�SXD"!U2d    ��D    ����G ���@ 	BLǕ�'� ��#� �D��BL��/c�MC�3�T0 k� �;��?�SXD"!U2d    ��D    ����G ���@ 	BLÕ�'� ��#� �D��BL��/c�M;�3�T0 k� �;��?�SXD"!U2d    ��D    ����G ���@ 	BLÕ�'� ��#� �D��BL��/_�M7�3�T0 k� �;��?�SXD"!U2d    ��D    ����G ���@ 	BLÕ�'� ��#� �D��BL��/_�M/�3�T0 k� �?��C�SXD"!U2d    ��D   ����G ���@ 	BLÕ�'� ��#� �D��BL��/[�M+�3�T0 k� �?��C�SXD"!U2d    ��D    ����G�+�C� 9C���s�nt�+�~��@lE>���<$3�T0 k� �3��7�SXD"!U2d    ��    ����[�'�C��9C���w�np|+�~��@lE>���4#3�T0 k� �+��/�SXD"!U2d    ��    ����X�#�C��:C���w�nl|/�~��@lE>���,#3�T0 k� �#��'�SXD"!U2d    ��    ����V��C��:C���w�nd |/�~��@nlE>���$"3�T0 k� ����SXD"!U2d    ��    ����T��C��;C��{�nc�|/�~��@nlE=���w�!3�T0 k� ����SXD"!U2d    ��    ����R��E��<C�{�{�n_�|/����@nlE=���o�!3�T0 k� ����SXD"!U2d    ��    ����P��E��<C�w���n[�|/����@npE=���g� 3�T0 k� �����SXD"!U2d    ��    ����N��E��=E�o���nS�|/����@npE����c� 3�T0 k� ������SXD"!U2d    ��    ����L��E�?E�g����nK�|/����E�pE����S��3�T0 k� ������SXD"!U2d    ��    ����J��E�?E�c����nG�|/����E�tE����K��3�T0 k� ������SXD"!U2d    ��    ����H���D>�@E�_����nC�|/����E�tE����G��3�T0 k� ������SXD"!U2d    ��    ����G���D>�AE�W����n?�|/����E�tG���?��3�T0 k� ������SXD"!U2d    ��    ����F���D>�BE�S����n;�|/����E�tG���7��3�T0 k� ������SXD"!U2d    ��    ����E���D>|CE�K����	�3�|/����E.xG���+��3�T0 k� ������SXD"!U2d    ��    ����D���D>pDE�G����	�/�|/����E.xG���#��3�T0 k� ������SXD"!U2d    ��    ����C                                                                                                                                                                            � � �  �  �  c A�  �J����  �      � \���4 ]�$$ � �����s     	   ��/�2    ��k�/�G    ��;                  Y��           	�  �  ���   (
          	Uv        ����O     	X�����    �� �                A��           �  �  ���   8�          ����  $ $      �0*c    ����0lC    |�                ��          �     ���   	@

          ��+�         ��P*    ��1��<�    ��"                    �$          c       ���   H
$
         ���`           .��4    ������_    ���                   �$           ��     ���  H
	!         ����  ��
     B���    �������                              ���}               ���      0            ����        V�@Pb    ��|��@Pb    �               	���G�         �        ��@   0
 
         ��ơ J J
    j�A�N    �����A�N    �                 	���G�        ���    ��@   0	%          ���: $ $      ~�/��    �����/��    ��               ���G         ��  �  ��H   8
          ��̏  � �
	   ����M    ��̏��V|      ��                ���G         	 &0�    ��`   8         ����  � �	    ��J3�    �����K��    ���g               9���G         
 @�    ��`  P
	
          �� �$	    � ��<     �� ��<                             ���O             N  ��@    P                   ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��{�  ��        ���47    ���W��1    ��� "                x                j  �       �                         ��    ��        ���      ��  ��           "                                                 �                         �/���0������@�A�/���J �������    
 	            
  �   i �z  ���J       �� �r@ �� s@ � s` �$ s� �D s� �d s� �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0� ���� � 
� U� 
�� V  
�| V ���� ����� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����G������ �  ������  
�fD
��L���"����D" � j  "  B   J jF�"    "�j * , ����
��"     �j @�    �
� �  �  
� ��    ��     ���      ��    ��     ���      ��    ��     ��/          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �D!!      �� � �  ��        �6T ���        �        ��        �        ��        �    ��    ������        ��                         �w� $ ��� ��                                    �                ����            �������%��  ���G ���`            6 Adam Burt k n h     6:02                                                                        3  3     � �
"� �)�)�2CBCD  CL �k~ � � k� �	B� � 
B� � �K � � K � �cV � �kj � �kr � � kt � �c� � � c� � �c� � �c� � � c� � �J�3 bC. � WC l C" a � � ` � � Ac� � A c� � B c� � : c� � 2  c� � * !c� � �""� � � #"� � v$� � v%
� � �&"� � � '"� � v("� � v)*� �*"� � +"�,� �-
� .* s �/!� s �0"8 � � 1"E { � 2"G �3* s 4"P �5" � 6"F �7!� s?8"6 sG 9"D �_  "C � � ;"A � � <" s � ="P � �>"* s "< �                                                                                                                                                                                                                         �� P @            @ 
        �     U P E Y  ��                    	�������������������������������������� ���������	�
��������                                                                                          ��    ��� 	  ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, $   p�� � � ���@���&�                                                                                                                                                                                                                                                                                                                                            �@���                                                                                                                                                                                                                                     
      	        ��   H�J                                     ������������������������������������������������������                                                                                                                                          �      �      h        �    ��              
 	  
	 
 	 	 ��������� ��� ���������������  �� ����������� ���� ���������� ������ ���� ����������� �������� ������� �������������� ����������������������������� � � �� ����� ��������������������������������������� ���������������������������� � ����������                                  j    )    ��  D�J    	  �  	                           ������������������������������������������������������                                                                      
                                                                    �      �      �        �        �  �          	  
 	 
 	 	 ������������ � �� ��������� ������ ������� ���������� ���� ��������������� ���������� ����� ������������ �������������� ������������� �������� ���� ����������� �� ����������������������������� ��������� ����������� ��������  �           �                                                                                                                                                                                                                                                                                                             �             


           �   }�        ��������   	��������   	������������   	����������������    ��������   	��������������������������������              '�           +                              '                      �ww�ww333wwwwwwww�ww�ww�ww�ww333wwww 4 G =                	                 � �y�h �\                                                                                                                                                                                                                                                                                     )n)h1p  �              k      `         W       k            a                                           ��                                                                                                                                                                                                                                                                                                                                                           � � �  � ��  � ��  � 2��  � 2��  � 7��  �����������g�����������h�����g�����E�����d����\�                ���@ : / z        	  	�   & AG� �   �   
              �                                                                                                                                                                                                                                                                                                                                      p C B   �      ��   #             !��                                                                                                                                                                                                                            Y��   �� � ��      �� Z      ��������� ��� ���������������  �� ����������� ���� ���������� ������ ���� ����������� �������� ������� �������������� ����������������������������� � � �� ����� ��������������������������������������� ���������������������������� � ���������������������� � �� ��������� ������ ������� ���������� ���� ��������������� ���������� ����� ������������ �������������� ������������� �������� ���� ����������� �� ����������������������������� ��������� ����������� ��������  �             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    &      2   � ��                       B     �  �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$ ^h  ��     �f ��     �f �$ ^$ �@      ����� ��   �����    ���� ��   ���� �$ ^$   �   �                      ������� 
� � ��� �� � ��� �$  � �  �� �  �      �   d   O���� e����� g��� 	 �     f ^�         �� ���      O      �������2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �   3       �  �3 3�=������<��̼��� �3 33==ƙ�<ə�ƙ�3ƙ��ƙ���i� 3= ��3=�l�ә��<��l<��l<��l<���<    �   3=  �30 ��� ���=��������                        +   3     0  �<  3� 3� =� =� 0� 0������������������3�33033�0�3�0��;f��;��̽�������3��3��<���<�f���̳=�=�������3303<�<00�<30�3����������������=��=��3�3�=�3�0  �=  �3  �3� ��0 ̳0 �0 �0  0� =� =� 3�  3�  �<  0  33�0�3�0�3�0�3303�303�303�303303��<���0<��0<033<033003300330033030�30�<00�<0330333033303330333033�0��<���0�03303303=03=03��0 ̳0 ��0 �3� �3� �=  0  3�     �                           <�03=��3=�� 3��  �=  �        033003300330�330��303= ��33    330333033303330333<��333ݰ    0=�0<3���;�3 �=  3�             �                           wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         7v` weV "fff"O�p"��p"��p"�p3�}p-��p=��p|� }�  }�  ��  ��  ��  ��  �  �  �  �  �  "              `  eV  fff O�  ��  ��  �  �} �� �� ��  |�  }�  ��    =   }   =   =              �������}�}�}�ww~r�� ∈�������������������}�� }�� ��� ��� ����   �   �   �   �   �   �   �   C""42""#2""#2""#2""#s3342"""3333    p   p   p   p   p   p   p    ��������� ��� }�� ��  ��  ����  ��  ��  ��  ��  ��  ��  ��                          � �� ��    "               wvf wfU 7Of`w��f"�� "�p-�}p���� ��� ����x��	�� �� �� "�        f  U` f` f` �p w���� `  eV  ff  O�  ��  �� ����}�                �  �  ��  �            �  �  �   �  ��  �                     �  �  �   � `  eV  ff  O�  ��  ��  ����}���������������p	���         `  eV  ff  O�  ��  ��  ���}�     �  �  �   �  ��  �   �            ��  ��  �   ��  �   ���������������p	���                    3333UUUU                        wwww                    333333333333333333333   w  G� ws@ ws� ws$7w@wwww"                               ����������� ��� �� ��  �    `  eV  ff  O�  ��  ��  � ��}�            """"                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "" "  """               "  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """               "  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  ""   "! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                      �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                 " �/����      �             "�"�����   �� �          ����   �       �                                   �    ���  ��                    ��  ��  ���   ���� �                                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �              "      �           �  �   �   ��  �                                        ��                     �   �                      �������  ���    �                    ��  ��  ���   ���� �                       ��� ���  �"  " ��"�""��"! � �  �   �   �   �                                                                                                                 �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   �   �"  ""  !� �� ��  �               �   ������  ��                      �   �                      �������  ���    �       �  �  �  �                �  �  �   �   ��  �                            �   ���                            �   �                                                                                                  �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ���� ��� ����                      �  �� ��  �    � ���                                                                                                                                                                                              �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �                "  "     �      �                         ���  +"  "" ���������                   �                        ���� ��� ����               �  �  �  �                 �       �                        �   ��  ���  � �    �                               �   �                                                                                                              �  ��� ��� ��� �ݪ�                       �   �    �z� 
�� ������������ ˍ� ��� ���������ˉ����� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��                    ˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                                         �  ��  �� ��  ��                    �   �   ��  ��  ��  ɀ  �   ��  ��  ���   �   �   �                                                       �         �  �� �  �� ��                                                       �  �  ��  �                                                                     �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   ��  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �   �   �                .                �  �� �� �� ��                         ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                   �  �˰ ��� w�� k}� gg��j�� ���
���	������ ��� ���˸�,̽�+�ӊ��8� �D 8�U�E �@ �� 	��  ��  � "" """/���  �                                 �   ��  ��  ��  ��� ̽� ̉  ɘ  �40 DD@ EU@ S3C  4M  ��  ��  *�  "�  "  ����� � �  �                          �   �                           �   �  "������"    /   �  �   ��                                �   �                      �������  ���    �    �  �  ��  �   �   �       ���                                  � ���� ��   � � �                                                                                                                                        �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �       /�      �                           �   �   �   �   �   �           �   �       �    �                     �   �  �  ��   �   ��� ������ �   �      �       �                        �   ��  ���  � �    �                                                                                                                                            �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��                     ��  ��  ���                                                    �   ���                            �   �                                                                                                     �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                �   ��  ��  ��  �  �   ��  ��                                                                                                                                                                                     �  ���ͻو  �� �˚̻��̽�����鋼�^���^�٘U�:�^��^�� U�( D�) �) �) �) ʹ� ˛� ț�+��,��,����  ��� ��� �ٝ ��ݨ��ډ�݊�� ��D@ �D�  ��� ��� ɫ� �۽ �ک ɺ��̻���諑���������������� �            �� ��� ��  �             �   ��  ��  ��  ��  ��                        �   �                         �   �          �  � � �� ��     �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(����������������� � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(����������������� 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5���������������� x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x���������������� w w x y�������H���������������������������������H������yxww����������������  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(���������������� , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,���������������� +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+���������������� 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5���������������� =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=����������������     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( ���������������� � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � ����������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
"� �)�)�2CBCD  CL �k~ � � k� �	B� � 
B� � �K � � K � �cV � �kj � �kr � � kt � �c� � � c� � �c� � �c� � � c� � �J�3 bC. � WC l C" a � � ` � � Ac� � A c� � B c� � : c� � 2  c� � * !c� � �""� � � #"� � v$� � v%
� � �&"� � � '"� � v("� � v)*� �*"� � +"�,� �-
� .* s �/!� s �0"8 � � 1"E { � 2"G �3* s 4"P �5" � 6"F �7!� s?8"6 sG 9"D �_  "C � � ;"A � � <" s � ="P � �>"* s "< �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������#� ��9�K�Z�X��5�R�O�S�G� � � � � � � � � � �/�.�7�����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�����������������������������������������!��+�J�G�S��,�[�X�Z� � � � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������2�0�.� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������/�.�7� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                