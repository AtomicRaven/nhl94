GST@�                                                           Zq     Z�                                               x&            �   H         � h� 2���J����������    ����        Ā      #    ����                                d8<n    �  ?    R�����  �
fD�
�L���"����D"� j   " B   J  jF�"    
 �j, 
���
��
�"    B�jl �   B ��
                                                                                  ����������������������������������      ��    =b 0Qb 4 114  4c  c  c      	 
      	   
       ��G �� � ( �(                 Enn )1         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                �   D       �   @  &   �   �                                                                                 'w w  E)n1n  �    �0   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E D �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��D2P�4  D�D6�PҜ8E��,� R	���Z<8T0 k� ������1d�'Qe1�t B  ��    ��� ����D2L�0  D�D6�L�8E��,��R	���Z<8T0 k� ������1d�'Qe1�t B  ��    ��� ����D2L�,  D�D6�H�8E��-��R	���Z<8T0 k� ������1d�'Qe1�t B  ��    ��� ����D2D�(  D�D6�@�8E��-���	���Z<8T0 k� ������1d�'Qe1�t B  ��    ��� ����D2@�$  D�D7�<�7E��-�{�� ���Z<8T0 k� ������1d�'Qe1�t B  ��    ��� ����D2<�$  D�D7�8��7E��-�s������Z<8T0 k� ������1d�'Qe1�t B  ��    ��� ����D28�   D�D7�4��7E��-�k������Z<8T0 k� ������1d�'Qe1�t B  ��    ��� ����D24�  D�D8�4��7E��-�_������Z<8T0 k� ������1d�'Qe1�t B  ��    ��� �b��DB0�  D�D8�0��7E��-�W�	�����Z<8T0 k� ������1d�'Qe1�t B  ��    ��� �b�DB( �  D�D:�(��7E��-�C�	�����Z<8T0 k� �� �� 1d�'Qe1�t B  ��    ��� �b�DB$ �  D�D:�$��7E��,�;�	���� Z<8T0 k� ����1d�'Qe1�t B  ��    ��� �b�DB !�  D�D;� ��7E��,�3�	����Z<8T0 k� �|��1d�'Qe1�t B  ��    ��� �b�DB!�   D�D;��7E��,�'�	����Z<8T0 k� �t�x1d�'Qe1�t B  ��    ��� �b�	DB"�   D�D<��7E��+��	����Z<8T0 k� �d�h1d�'Qe1�t B  ��    ��� ~b�DB#��  D�H<� 6E��+��	����Z<8T0 k� �\	�`	1d�'Qe1�t B  ��    ��� {b�DB#��  D�L=�6E� +��	����Z<8T0 k� �T
�X
1d�'Qe1�t B  ��    ��� xb�DB $��  D�P=�6ED +@������Z<8T0 k� �P�T1d�'Qe1�t B  ��    ��� ub�DQ�%��  D�P>�5ED *@������Z<8T0 k� �H�L1d�'Qe1�t B  ��    ��� rr�DQ�&��  D�X?�5ED *@�����	Z<8T0 k� �@�D1d�'Qe1�t B  ��    ��� or�DQ�'��  D�X?�4ED )@�����
Z<8T0 k� �<�@1d�'Qe1�t B  ��    ��� lr�DQ�(��  D�\@� $4ED )@�����
Z<8T0 k� �8�<1d�'Qe1�t B  ��    ��� ir|DQ�)��  D�\@���(4ED (@����Z<8T0 k� �4�81d�'Qe1�t B  ��    ��� frtDQ�)��  D�`@�� �03ED (@����Z<8T0 k� �0�41d�'Qe1�t B  ��    ��� crlDQ�*��  D�`@�� �43ED '@����Z<8T0 k� �(�,1d�'Qe1�t B  ��    ��� `�hDQ�+��  D�d@�� �<2EC�'@��� �Z<8T0 k� �(�,1d�'Qe1�t B  ��    ��� ^�`DQ�,��  D�dA�� �D2C��&���� �Z<8T0 k� �,�01d�'Qe1�t B  ��    ��� [�TDQ�.�  D�dA����P1C��$���� �Z<8T0 k� � �$1d�'Qe1�t B  ��    ��� Y�LDa�/�  D�hAr���X0C��$�{�� �Z<8T0 k� � �$1d�'Qe1�t B  ��    ��� V�HDa�0�  D�hAr���\/C��#�s�� �Z<8T0 k� �� 1d�'Qe1�t B  ��    ��� T�@Da�1ќ  D�hAr���d/C��"@g��| �Z<8T0 k� ��1d�'Qe1�t B  ��    ��� R�8 Da�2ј  D�hAr���l.C��!@_��t �Z<8T0 k� ��1d�'Qe1�t B  ��    ��� P�4!Da�3ѐ  D�hAr���p-C�� @S��l �Z<8T0 k� ��1d�'Qe1�t B  ��    ��� N�,"Da�5ш  D�hAr��sx,C��@K��h �Z<8T0 k� � � 1d�'Qe1�t B  ��    ��� Lb$#Da�6р  D�hAr��s�+C��@C��` �Z<8T0 k� ��!��!1d�'Qe1�t B  ��    ��� Jb%Da�8�p  A�hA���s�*C��@/��PxZ<8T0 k� ��#��#1d�'Qe1�t B  ��    ��� Hb&Da|9�h  A�hA���s�)C��@#�HtZ<8T0 k� ��$��$1d�'Qe1�t B  ��    ��� Eb'Dat;�`  A�hA���s�'C��@�DlZ<8T0 k� ��%��%1d�'Qe1�t B  ��    ��� B�(D1p<�X  A�hA���s�&C��0�<hZ<8T0 k� ��%��%1d�'Qe1�t B  ��    ��� @��)D1h=�P  A�hA��s�%C��0�4`Z<8T0 k� ��&��&1d�'Qe1�t B  ��    �   >��*D1`>�H  A�hA��s�$C��?��,\Z<8T0 k� ��'��'1d�'Qe1�t B  ��    �  <��*D1\?�@  A�hA��s�$C��?��$TZ<8T0 k� ��(��(1d�'Qe1�t B  ��    �  :��+D1TA�8  A�hA��s�#C��?��PZ<8T0 k� ��)��)1d�'Qe1�t B  ��    �  8��,D1LB�4  A�hA��c�"C��?��HZ<8T0 k� ��%��%1d�'Qe1�t B  ��    �  6��-D1HC�,  A�hA��c�!C��?��DZ<8T0 k� ��!��!1d�'Qe1�t B  ��    �  4��-D1@D�$  A�hA��c� C��?�� �<Z<8T0 k� ����1d�'Qe1�t B  ��    �  2��.D18F�  A�hA��c�C��?�� ��4Z<8T0 k� ����1d�'Qe1�t B  ��    �  0��/D14G�  A�hA��c�C��
?����0Z<8T0 k� ����1d�'Qe1�t B  ��    �  .��/D1,H�  A�hA��c�C��/� ��(Z<8T0 k� ����1d�'Qe1�t B  ��    �  ,��0D1$I�  A�hA��c�C��/���$Z<8T0 k� ����1d�'Qe1�t B  ��    �  )��0DA K��   A�hAs�c�C��/��	�Z<8T0 k� �� �� 1d�'Qe1�t B  ��    �  &��1DAL��   A�hAs�S�C��/��	�Z<8T0 k� �x!�|!1d�'Qe1�t B  ��    � 	 $��1DAM���  A�hAs�S�EӴ/��	�Z<8T0 k� �p"�t"1d�'Qe1�t B  ��    � 	 "Q�2DAN���  A�hAs�S�Eӳ�/��	�Z<8T0 k� �l(�p(1d�'Qe1�t B  ��    � 
  Q�2DAP���  A�hAs�S�Eӯ�/��	� Z<8T0 k� �h-�l-1d�'Qe1�t B  ��    � 
 Q�2EP�Q���  AShAs�S�Eӫ�/��	� Z<8T0 k� �d0�h01d�'Qe1�t B  ��    � 
 Q�3EP�R���  AShAs�S�Eӧ�/��	�  Z<8T0 k� �`3�d31d�'Qe1�t B  ��    �  Qx3EP�S���  AShAs�S�Eӣ�/�
�	�� Z<8T0 k� �X5�\51d�'Qe1�t B  ��    �  Qp4EP�T���  AShAs�S�Eӛ�/|��	�� Z<8T0 k� �P7�T71d�'Qe1�t B  ��    �  Qh4EP�V���  AShAs#���Eӗ�/x��	�� Z<8T0 k� �H8�L81d�'Qe1�t B  ��    �  Q`5EP�W��  AShAs#���C��t��	�� Z<8T0 k� �@:�D:1d�'Qe1�t B  ��    �  QX5EP�X ��  AShAs#���C��p�x	�� Z<8T0 k� �8;�<;1d�'Qe1�t B  ��    �  QP5EP�Y ��  AShAs'��C��l�p	�� b�8T0 k� �0;�4;1d�'Qe1�t B  ��    �  QH6C��Z ��  AShAs'��C��h�h	�� b�8T0 k� �(<�,<1d�'Qe1�t B  ��    �  A@6C��[ ��  AShAs+��C�{�d�\	�� b�8T0 k� � ?�$?1d�'Qe1�t B  ��    �  	A87C�\ ��  AShAs/��C�w�`�T	�� b�8T0 k� �B�B1d�'Qe1�t B  ��    �  A07C�]p��  AShAs/��C�o�\�L	�� b�8T0 k� �C�C1d�'Qe1�t B  ��    �  A(8C�^p��  AShAs3��C�g��\�D	�� b�8T0 k� �E�E1d�'Qe1�t B  ��    �  A$8E�_p��  AShAs7��C�c��X�<	�� b�8T0 k� � F�F1d�'Qe1�t B  ��    �  9E��`p��  AShAs;��C�[��X�4	�� b�8T0 k� ��G��G1d�'Qe1�t B  ��    � ��9E��bp��  AShA�?��
C�S��T�,	�� b�8T0 k� ��G��G1d�'Qe1�t B  ��    � ��:E��cp��  AShA�?��	C�K��T� 	�� b�8T0 k� ��H��H1d�'Qe1�t B  ��    � ��:E��dp�  AShA�?��	C�G��T�	�� b�8T0 k� ��H��H1d�'Qe1�t B  ��    � ���;E��epw�  AShA�?��C�?��T�	�� Z<8T0 k� ��I��I1d�'Qe1�t B  ��    � ���<E�xf`s�  AShA�?��C�7� oP�	��!Z<8T0 k� ��J��J1d�'Qe1�t B  ��    � ���<D0pg`o�  AShAs?��C�/� oP���!Z<8T0 k� ��J��J1d�'Qe1�t B  ��    � ���=D0lh`k�  AShAs?��C�'� oP���!Z<8T0 k� ��K��K1d�'Qe1�t B  ��    � ���>D0di`g�  AShAs?��C�#� oP � ��!Z<8T0 k� ��L��L1d�'Qe1�t B  ��    � ���>D0\k`_�  AShAs?��C�� oP!��ϼ!Z<8T0 k� ��L��L1d�'Qe1�t B  ��    � ���?D0Tl`[�  AShAs?��C���P"��ϸ"Z<8T0 k� ��M��M1d�'Qe1�t B  ��    � ���@D0Pm`W�  AShAs?��|C���L#����"Z<8T0 k� ��N��N1d�'Qe1�t B  ��    � �� �@D0Hn`S�  AShAs?�SxC���L%���"Z<8T0 k� ��N��N1d�'Qe1�t B  ��    � �� �AD0@o`K�  AShAs?�StC����L&���"Z<8T0 k� ��O��O1d�'Qe1�t B  ��    � �� �BD0<p`G�  AShAs?�StD���L'���"Z<8T0 k� ��P��P1d�'Qe1�t B  ��    � �� �BD04rPC�  AShAs;�StD���L)���"b|8T0 k� �xP�|P1d�'Qe1�t B  ��    � �� �CD0,sP?�  AShAs;�SpD���H*���"b|8T0 k� �pQ�tQ1d�'Qe1�t B  ��    � ��МDD0$tP7�  AShAs;�SlD���H,���!b|8T0 k� �lN�pN1d�'Qe1�t B  ��    � ��ДDD@ uP3�  AShAs;�SlD���H-���!b|8T0 k� �hK�lK1d�'Qe1�t B  ��    � ��ЌED@vP/�  AShAs;�ChD���D/���!b|8T0 k� �dI�hI1d�'Qe1�t B  ��    � ��ЄFD@xP'�  AShAs;�ChD���D0���!b|8T0 k� �\H�`H1d�'Qe1�t B  ��    � ���|FD@yP#�  AShAs;�CdD���D2���!b|8T0 k� �TG�XG1d�'Qe1�t B  ��    � ��@xGD@zP�  AShAs;�CdD���@3���!b|8T0 k� �TL�XL1d�'Qe1�t B  ��    � ��@pHE_�{P�  AShAs;�C`D���@5���!b|8T0 k� �LP�PP1d�'Qe1�t B  ��    �  ��@hHE_�|P�  AShAs;��\D���<7��� b|8T0 k� �@R�DR1d�'Qe1�t B  �    � !��@XJE_�~P�  AShA�;��XD���8:��t b|8T0 k� �,W�0W1d�'Qe1�t B  ��   � "��`TKE_�_��  AShA�?��TD���4;��p Z<8T0 k� � Y�$Y1d�'Qe1�t B  ��   � #��`LKE_؀_��  AShA�?��PD���0=��l Z<8T0 k� �[�[1d�'Qe1�t B  ��   � $��`DLE_ԀO��  AShA�C��LD{��0?�
d Z<8T0 k� �]�]1d�'Qe1�t B ��   � %��`<LE_̀O��  AShA�C��HDs��,@�
` Z<8T0 k� � `�`1d�'Qe1�t B ��   � &��`8ME_ĀO��  AShA�G��DDk��(A�
XZ<8T0 k� ��b��b1d�'Qe1�t B ��   � '��p0NE_�O��  AShA�K��<Dc�	�(C�
TZ<8T0 k� ��d��d1d�'Qe1�t B ��   � (��p(NE_�O��  AShA�K��8D[�	�$D�
LZ<8T0 k� ��f��f1d�'Qe1�t B ��   � )��p$OE_�O��  AShA�O��4DS�	�$E�|
HZ8T0 k� ��i��i1d�'Qe1�t B ��   � *��pPE_�OϿ  AShA�S��0DK�	� F�t
@Z8T0 k� ��k��k1d�'Qe1�t B ��   � +��pPE_�~Oǿ  AShA�W��(C�C�	� H�l
<Z8T0 k� ��m��m1d�'Qe1�t B ��   � ,���QE_�~O��  AShA�[��$C�;�	� I�h
4Z8T0 k� ��o��o1d�'Qe1�t B �� 	  � -���QE_�~O��  AShA�_�� C�3�	�J�`
/0Z8T0 k� ��r��r1d�'Qe1�t B  �� 	  � .���RE_�~O��  AShA�c��C�+�	�K�X
/(Y�8T0 k� ��t��t1d�'Qe1�t B  �� 	  � /��� RE_�}?��  AShA�g��C�#�	�L�P
/ Y�8T0 k� ��u��u1d�'Qe1�t B  �� 	  � 0����SAo�}?��  AShA�k��C��	�M�H
/Y�8T0 k� �lv�pv1d�'Qe1�t B  �� 	  � 1����SAox}?��  AShA�s��C��ON�<
/Y�8T0 k� �Tw�Xw1d�'Qe1�t B  �� 	  � 2����UAoh|?��  AShA�{���C���OP�,
/Y|4T0 k� �<w�@w1d�'Qe1�t B  /� 	  � 3����UAo`|?��  AShA�����C���OQ�$
/ Y|4T0 k� �(x�,x1d�'Qe1�t B  �� 	  � 4����VAo\|O��  AShA�����C��OS�
.�Y|4T0 k� �x�x1d�'Qe1�t B  �� 	  � 5����VE_T|O�  AShA�����C��OT�
.�Y|4T0 k� �v�v1d�'Qe1�t B  �� 	  � 6����WE_L{O{�  AShA�����C�߷OU�
.�Y|4T0 k� �u�u1d�'Qe1�t B  �� 	  � 7����WE_D{Os�  AShA�����C�׶	V�
�Z�4T0 k� �t�t1d�'Qe1�t B  �� 	  � 8����XE_<{Oo�  AShA�����C�϶	X��
�Z�4T0 k� �s�s1d�'Qe1�t B  �� 
  � 9����XE_4{Ok�  AShA���B�	C�ǵ	Y��
�Z�4	T0 k� �r�r1d�'Qe1�t B  �� 
  � :����YE_ zO_�  AShA���B�	C�	 [��
�Z�4	T0 k� ��q� q1d�'Qe1�t B  �� 
  � ;����YEOzOW�  AShA���B�
C�	~�\��
�Z�4	T0 k� ��n��n1d�'Qe1�t B  �� 
  � <�}��ZEOzOS�  AShA���B�
C�	��]��
�Z�4
T0 k� ��k��k1d�'Qe1�t B  �� 
  � <�{��ZEOyOO�  AShA���B�C�	��^��
�Z�4
T0 k� ��j��j1d�'Qe1�t B  �� 
  � <�x��[EO yOG�  AShA���B�C�	��^�
�Z�4
T0 k� ��i��i1d�'Qe1�t B  �� 
  � <�vO�[EN�y_C�  AShA�����C�	��_�

�Z�4
T0 k� ��h��h1d�'Qe1�t B  �� 
  � <�tO�\A�x_?�  AShA�����D��	��`�

�Z�4
T0 k� ��g��g1d�'Qe1�t B  �� 
  � <�rO�]A�x_3�  AShA����xDo���b�

>�Z�4
T0 k� ��f��f1d�'Qe1�t B  �� 
  � <�pO�]A�w_/�  AShA����pDg���c^�	
>�Z�4
T0 k� ��f��f1d�'Qe1�t B  �� 
  � <�nO�^A�w_+�  AShA����hD_���c^�	
>xZ�4
T0 k� ��f��f1d�'Qe1�t B  ��   � <�kO�_A�v_'�  AShA����\DW���d^�	
>pZ�4
T0 k� ��e��e1d�'Qe1�t B  ��   � <�iO�_A�v_#�  AShA����TDO���e^x	
>hZ�0
T0 k� ��e��e1d�'Qe1�t B  ��   � <�gO|`A�u_�  AShA����LDG���f^p
>`Z�0
T0 k� ��d��d1d�'Qe1�t B  ��   � <�eOxaA�u_�  AShA����DD;���g^h
>XZ�0
T0 k� �xd�|d1d�'Qe1�t B  ��   � <�c?pbA�t_�  AShA����<D3���h^`
>PZ�0
T0 k� �lc�pc1d�'Qe1�t B  ��   � <�a?lbA.�to�  AShA����4D+���i^X
>HZ�0T0 k� �hc�lc1d�'Qe1�t B  ��   � <�_?hcA.�so�  AShA����,D#���j^P
>DZ�0T0 k� �db�hb1d�'Qe1�t B  ��   � <�]?ddA.�so�  AShA����$D���kNH
<Z�0T0 k� �\a�`a1d�'Qe1�t B  ��   � <�[?\eA.�ro�  AShA����D���lN@
4Z�0T0 k� �Ta�Xa1d�'Qe1�t B  ��   � <�Y?TgA.xq���  AShA����D����nN,
$Z�0T0 k� �D_�H_1d�'Qe1�t B  ��   � <�W?PhA.pp���  AShA���� D����nN$
Z�0T0 k� �<_�@_1d�'Qe1�t B  ��   � <�U?LiA.hp���  AShA�����D���oN
Z�0T0 k� �4^�8^1d�'Qe1�t B  ��   � <�S?DjA.`o���  AShA�����D���pN
Z�0T0 k� �,^�0^1d�'Qe1�t B  ��   � <�Q?@lA.Xn���  AShA�����Dߧ��qN
Z�0T0 k� �$]�(]1d�'Qe1�t B  ��   � <�O?<mA.Pn���  AShA�����DӦ��qN
 Z�0T0 k� �\� \1d�'Qe1�t B  ��   � <�M/8nA>Hm���  AShA�����D˦�rM�
�Z�0T0 k� �Z�Z1d�'Qe1�t B  ��   � <�K/4oA>@l���  AShA�����C�æ�sM�
�Z�0T0 k� �Y�Y1d�'Qe1�t B  ��   � <�I/0qA>8k���  C�hA�����C໥>�s=�
�Z�0T0 k� �X�X1d�'Qe1�t B  ��   � <�G/,rA>0k���  C�hA����C೥>�t=�
-�Z�0T0 k� � W�W1d�'Qe1�t B  ��   � <�F/(sA>(j���  C�hA����C૤>�t=�
-�Z�0T0 k� ��V��V1d�'Qe1�t B  ��   � <�E/$tEN i޻�  C�hA����C���>�t=�
-�Z�0T0 k� ��V��V1d�'Qe1�t B  ��   � <�D/$vENh޷�  C�dA����C���>�u=�	
-�Z�0T0 k� ��U��U1d�'Qe1�t B  ��   � <�C/yENgޫ�  C�dA����C����u=�	
-�Z�0T0 k� ��S��S1d�'Qe1�t B  ��   � <�B/xENfޣ�  C�`A����C���u=�
-�Z�0T0 k� ��R��R1d�'Qe1�t B  ��   � <�A/xEM�e��  C�`A����C�w��u=�-�Z�0T0 k� ��R��R1d�'Qe1�t B  ��   � <�@xEM�d��  C�\A����xC�k��uM�-�Z�0T0 k� ��Q��Q1d�'Qe1�t B  ��   � <�?wE=�c��  C�\A����pC�c��|uM�-�Z�0T0 k� ��O��O1d�'Qe1�t B  ��   � <�>wE=�b��  C�XA����hC�[��tuM�-�Z�0T0 k� ��N��N1d�'Qe1�t B  ��   � <�=wE=�a��  C�TA���`C�S��puM�-�Z�0T0 k� ��M��M1d�'Qe1�t B  ��   � <�<vE=�`��  C�TA���XC�K��huM�-�Z�0T0 k� ��L��L1d�'Qe1�t B  ��   � <�;�vE=�_�w�  C�PA���LC�?��duM�-�Z�0T0 k� ��K��K1d�'Qe1�t B  ��   � <�:�uE=�^�o�  C�LA���DC�7��\uM|-�Z�0T0 k� ��J��J1d�'Qe1�t B  ��   � <�9�uE=�]�k�  C�HA���<C�/��XuMx-�Z�0T0 k� ��I��I1d�'Qe1�t B  ��   � <�8�uE=�\�c�  C�DA���4C�'��PtMx
MxZ�0T0 k� ��G��G1d�'Qe1�t B  ��   � <�8�tE=�[�[�  C�@A���, C���Lt=p
MpZ�0T0 k� ��F��F1d�'Qe1�t B  ��   � <�8�sE=�X�O�  C�<A��� C���@s=d
M`Z�0T0 k� ��D��D1d�'Qe1�t B  ��   � <�8�rE=�W�K�  C�4A���!C���8r=\
M\Z�0T0 k� ��B��B1d�'Qe1�t B  ��   � <�8�rE-�V�C�  C�0A���!D���4r=XTZ�0T0 k� ��B��B1d�'Qe1�t B  ��   � <�8�qE-�T�;�  D,A��� !D��,q=PL Z�0T0 k� ��A��A1d�'Qe1�t B  ��   � <�8�qE-�S�3�  D(A����"D��(p=HL Z�0T0 k� ��A��A1d�'Qe1�t B  ��   � <�8�pE-�R�/�  D$A����"Dߝ�$p=HL Z�0T0 k� ��A��A1d�'Qe1�t B  ��   � <�8�oE-�P�'�  D A����"Dל�o=@D!Z�0T0 k� ��?��?1d�'Qe1�t B  ��   � <�8�nF�|O��  DA����#DϜ�n-<	@!Z�0T0 k� ��>��>1d�'Qe1�t B  ��   � <�8�nF�xN��  DA����#Dǜ�m-4	<!Z�0T0 k� ��=��=1d�'Qe1�t B  ��   � <�8�mF�tM��  DA����#D���l-4	8"Z�4T0 k� ��<��<1d�'Qe1�t B  ��   � <�8�lF�lK��  DA����$D���k-0	4"Z�4T0 k� ��:��:1d�'Qe1�t B  ��   � <�8�kF�hJ��  DA����$D���j-,	,#Z�4T0 k� ��9��91d�'Qe1�t B  ��   � <�8�jF�dI��  D�A����$D��� i�(	-,#Z�4T0 k� ��8��81d�'Qe1�t B  ��   � <�8�iF�\H��  D�A����$D����h� 	-(#Z�4T0 k� ��7��71d�'Qe1�t B  ��   � <�8�hF�XG��  D�A����%D����f�	-$#Z�4T0 k� ��6��61d�'Qe1�t B  ��   � <�8� gF�TF��  D�A�����%D����e�	- $Z�4T0 k� �x5�|51d�'Qe1�t B  ��   � <�8� fF�PD��  D�A�����%D���d�	-$Z�4T0 k� �t4�x41d�'Qe1�t B  �   � <�8�(eF�DB���  D�A�����&Do���a-%Z�4T0 k� �l1�p11d�'Qe1�t B  �   � <�8O(dF�@A���  AR�A���Px&A_g���`-%Z�4T0 k� �d0�h01d�'Qe1�t B  ��   � <�8O,cF�<@���  AR�A���Pp&A__���_-%Z�8T0 k� �`/�d/1d�'Qe1�t B  ��   � <�8O,bF�8?ݿ�  AR�A���Ph'A_W���]-&Z�8T0 k� �\.�`.1d�'Qe1�t B  ��   � <�8O0aF�4>ݷ�  AR�A���P`'A_K���\-&Z�8T0 k� �X-�\-1d�'Qe1�t B  ��   � <�8O0`F�,=ݯ�  AR�A���PX'A_C���[-'Z�8T0 k� �T,�X,1d�'Qe1�t B  ��   � <�8O4_F�(<ݫ�  AR�A���PP'A_;���Z�'Z�8T0 k� �P+�T+1d�'Qe1�t B  ��   � <�8O8^F�$;ݣ�  AR�A���PH'A_7���X�(Z�8T0 k� �H*�L*1d�'Qe1�t B  ��   � <�8O8]F� :]�   AR�A���P@(A_/���W� )Z�8T0 k� �D)�H)1d�'Qe1�t B  ��   � <�8O<\F�9]�  AR�A���P8(A_'���V� )Z�8T0 k� �@(�D(1d�'Qe1�t B  ��   � <�8O<[F�8]�  AR�A���P0(A_���U�  )Z�8T0 k� �<'�@'1d�'Qe1�t B  �   � <�8O@[F�8]�  AR�A���P((A_���T� �)Z�8T0 k� =<'�@'1d�'Qe1�t B  ��   � <�8O@ZF�8]�  AR�A���P$)A_���S� �)Z�<T0 k� =<&�@&1d�'Qe1�t B  ��   � <�8ODYF�8]|  AR�A���P)A_���R� �)Z�<T0 k� =8&�<&1d�'Qe1�t B  ��   � <�8ODXF�8]t  AR�A���P)A_���P� �*Z�<T0 k� =8&�<&1d�'Qe1�t B ��   � <�8ODWF�8]p  AR�A���P)A^����O� �*Z�<T0 k� =4%�8%1d�'Qe1�t B ��   � <�8OHWF�8]h  AR|A���P)A^���N� �*Z�<T0 k� �4%�8%1d�'Qe1�t B ��   � <�8OHVF�8]d  ARxA���P *A^���M� �*Z�<T0 k� �4$�8$1d�'Qe1�t B ��   � <�8OLUF�8]`  ARtA���_�*A^���L� �*Z�<T0 k� �0$�4$1d�'Qe1�t B ��   � <�8OLTF�7]X  ARlA���_�*A^ߖ��K� �*Z�<T0 k� �0%�4%1d�'Qe1�t B ��   � <�8OPTF�7]T  ARhA���_�*A^ۖ��J� �*Z�<T0 k� �0&�4&1d�'Qe1�t B ��   � <�8OPSF�7]P  ARdA���_�*A^ӕ��I� �*Z�<T0 k� �0'�4'1d�'Qe1�t B ��   � <�8OTRF�6]H  AR`A���_�+A^ϕ��H� �*Z�<T0 k� �4'�8'1d�'Qe1�t B ��   � <�8OTQF�6]D	  AR\A���_�+A^Ǖ��G� �*Z�@T0 k� �4(�8(1d�'Qe1�t B ��   � <�8OTQF�5]@	  ARXA���_�+A^Õ��G�  �*Z�@T0 k� �4(�8(1d�'Qe1�t B ��   � <�8OXPF�5]<
  ARTA���_�+A^����F�   �+Z�@T0 k� �8)�<)1d�'Qe1�t B ��   � <�8OXOF�4]8
  ARPA���_�+A^����E� ! �+Z�@T0 k� M8)�<)1d�'Qe1�t B ��   � <�8O\OF�3]0  ARHA���_�,A^����D� ! �+Z�@T0 k� M8*�<*1d�'Qe1�t B ��   � <�8O\NF�3],  ARDA���_�,A^���|C� " �+Z�@T0 k� M8*�<*1d�'Qe1�t B ��   � <�8O\NF�2](  AR@A���_�,A^���|B�$" �+Z�@T0 k� M<*�@*1d�'Qe1�t B ��   � <�8O`MF�2]$  AR<A���_�,A^���xA�$" �+Z�@T0 k� M4%�8%1d�'Qe1�t B  ��   � <�8O`LF�2]   AR8A���_�,A^���tA�(" �+Z�@T0 k� -0 �4 1d�'Qe1�t B  ��   � <�8O`LF�2]  AR4A���_�,A^���t@�(" �+Z�@T0 k� -0�41d�'Qe1�t B  ��   � <�8OdKF�2]  AR0A���_�,A^���p?�(" �+Z�@T0 k� -,�01d�'Qe1�t B  ��   � <�8OdKF�1]  AR,A���_�-A^���l>�," �+Z�@T0 k� -,�01d�'Qe1�t B  /�   � <�8OdJF�1]  AR,A���_�-A^���l=�," �+Z�@T0 k� -0�41d�'Qe1�t B  ��   � <�8OhIF�1]  AR(A���_�-A^���h=�," �+Z�DT0 k� =0�41d�'Qe1�t B  ��   � <�8OhIF�1]  AR$A���_�-A^{��d<�0! �,Z�DT0 k� =4�81d�'Qe1�t B  ��   � <�8OhHF�1]  AR A���_�-A^w��d;�0! �,Z�DT0 k� =4�81d�'Qe1�t B  ��   � <�8OlHF�1]   ARA���_�-A^s��`:�4! �,Z�DT0 k� =8�<1d�'Qe1�t B  ��   � <�8OlGF�0\�  ARA���_�.A^o��`:�4! �,Z�DT0 k� =8�<1d�'Qe1�t B  ��   � <�8OlGF�0\�  ARA���_�.A^k��\9�8! �,Z�DT0 k� �8�<1d�'Qe1�t B  ��   � <�8OpFB�/\�  ARA���_|.A^g��X8�8  �,Z�DT0 k� �<�@1d�'Qe1�t B  ��   � <�8OpFB�/\�  ARA���_x.A^_��X8�8  �,Z�DT0 k� �<�@1d�'Qe1�t B  ��   � <�8OpEB�.\�  ARA���_t.A^[��T7�<  �,Z�DT0 k� �@�D1d�'Qe1�t B  ��   � <�8OtEB�.\�  ARA���_p.A^W��T6�<  �,Z�DT0 k� �@�D1d�'Qe1�t B  ��   � <�8OtDB�.\�  ARA���_l.A^S��T6�@ �,Z�DT0 k� �@�D1d�'Qe1�t B  ��   � <�8OtDB�.\�  AR A���_h.A^O��T6�@ �,Z�DT0 k� �D�H1d�'Qe1�t B  ��   � <�8OtCB�-\�  AR A���_d/A^K��T6�D �,Z�DT0 k� �D�H1d�'Qe1�t B  ��   � <�8OxCB�-\�  AQ�A���_`/A^G��T5�D �,Z�DT0 k� �H�L1d�'Qe1�t B  ��   � <�8OxBB�-\�  AQ�A���_\/A^C��T5�H �,Z�DT0 k� �H�L1d�'Qe1�t B  ��   � <�8OxBB�,\�  AQ�A���_X/A^?��T5�H �-Z�DT0 k� �L�P1d�'Qe1�t B  ��   � <�8O|BB�+\�  AQ�A���_T/A^;��T4�L �-Z�DT0 k� �L�P1d�'Qe1�t B  ��   � <�8O|AE�*\�  AQ�A���_P/A^7��T4�L �-Z�HT0 k� �P�T1d�'Qe1�t B  ��   � <�8O|AE�*\�  AQ�A���_L/A^3��T4�P |-Z�HT0 k� �P�T1d�'Qe1�t B  ��   � <�8O|@E� )\�  AQ�A���_H/A^/��T3�P |-Z�HT0 k� �T�X1d�'Qe1�t B  ��   � <�8O�@E� (\�  AQ�A���_D0A^/��T3 }T x-Z�HT0 k� �\�`1d�'Qe1�t B  ��   � <�8O�?E� '\�  AQ�A���_@0A^+��T3 }T x-Z�HT0 k� �d�h1d�'Qe1�t B  ��   � <�8O�?E� &\�  AQ�A���_<0A^'��P2 }X t-Z�HT0 k� �h �l 1d�'Qe1�t B  ��   � <�8O�?E� &\�  AQ�A���_<0A^#��P2 }X t-Z�HT0 k� �p$�t$1d�'Qe1�t B  ��   � <�8O�>E�$%\�  AQ�A���_80A^��P2 }\ t-Z�HT0 k� �x'�|'1d�'Qe1�t B  ��   � <�8O�>E�$$\�  AQ�A���_40A^��P1 }` p-Z�HT0 k� �|)��)1d�'Qe1�t B  ��   � <�8O�>E�$#\�  AQ�A���_00A^��P1 }` p-Z�HT0 k� ��+��+1d�'Qe1�t B  ��   � <�8O�=@�$#\�  AQ�A���_,0A^��P1 }d l-Z�HT0 k� ��,��,1d�'Qe1�t B  ��   � <�8O�=@�$"\�  AQ�A���_,0A^��P0-h l-Z�HT0 k� ��+��+1d�'Qe1�t B  ��   � <�8O�<@�$!\�  AQ�A���_(1A^��P0-l h-Z�HT0 k� ��*��*1d�'Qe1�t B  ��   � <�8O�<@�(!\�  AQ�A���_$1A^��P0-l h-Z�HT0 k� ��)��)1d�'Qe1�t B  ��   � <�8O�<@�( \�  AQ�A���_ 1A^��P0-p d-Z�HT0 k� ��)��)1d�'Qe1�t B  ��   � <�8O�;@�(\�  AQ�A���_ 1A^��P/-t d-Z�HT0 k� ��)��)1d�'Qe1�t B  ��   � <�8O�;@�(\�  AQ�A���_1A^��P/x d-Z�HT0 k� ��$��$1d�'Qe1�t B  ��   � <�8O�;@�(\�  AQ�A���_1A]���P/| `.Z�HT0 k� �� �� 1d�'Qe1�t B  ��   � <�8O�:@�(\�  AQ�A���_1A]���P.� `.Z�HT0 k� ����1d�'Qe1�t B  ��   � <�8O�:@�,\�  AQ�A���_1A]���P.� \.Z�HT0 k� ����1d�'Qe1�t B  ��   � <�8O�:@�,\�  AQ�A���_1A]���P.� \.Z�HT0 k� ����1d�'Qe1�t B  ��   � <�8O�:@�,\�  AQ�A���_1A]���P. -� \.Z�LT0 k� ����1d�'Qe1�t B  ��   � <�8O�9@�,\�  AQ�A���_1A]��P- -� X.Z�LT0 k� ����1d�'Qe1�t B  ��   � <�8O�9@�,\�  AQ�A���_2A]��P- -� X.Z�LT0 k� ����1d�'Qe1�t B  ��   � <�8O�9@�,\�  AQ�A���_2A]��P- -� X.Z�LT0 k� ����1d�'Qe1�t B  ��   � <�8O�8@�,\�  AQ�A���_2A]��P- -� T.Z�LT0 k� ����1d�'Qe1�t B  ��   � <�8O�8@�0\�  AQ�A���_ 2A]��P, -� T.Z�LT0 k� ����1d�'Qe1�t B  ��   � <�8O�8@�0\�  AQ�A���_ 2A]��P, -� T.Z�LT0 k� ��� 1d�'Qe1�t B  ��   � <�8O�8@�0\�  AQ�A���^�2A]��P, -� P.Z�LT0 k� ��1d�'Qe1�t B  ��   � <�8O�7@�0\�  AQ�A���^�2A]��P, -� P.Z�LT0 k� ��1d�'Qe1�t B  ��   � <�8O�7@�0\�  AQ�A���^�2A]ߏ�L, -� P.Z�LT0 k� ��1d�'Qe1�t B  ��   � <�8O�7@�0\�  AQ�A���^�2A]ۏ�L+ -� L.Z�LT0 k� ��1d�'Qe1�t B  ��   � <�8O�7@�0\�  AQ�A���^�2A]ۏ�L+ -� L.Z�LT0 k� � �$1d�'Qe1�t B  ��   � <�8O�6@�0\|  AQ�A���^�2A]׏�L+ =� L.Z�LT0 k� �,�01d�'Qe1�t B  ��   � <�8O�6@�4\|  AQ�A���^�2A]׏�L+ =� H.Z�LT0 k� �4�81d�'Qe1�t B  ��   � <�8O�6@�4\|  AQ�A���^�2A]ӏ�L* =� H.cLT0 k� �@�D1d�'Qe1�t B  ��   � <�8O�6@�4\x  AQ�A���^�3A]ӏ�L* =� H.cLT0 k� �L�P1d�'Qe1�t B  ��   � <�8O�5@�4\x  AQ�A���^�3A]Ϗ�L* =� D.cLT0 k� �T�X1d�'Qe1�t B  ��   � <�8O�5@�4\x  AQ�A���^�3A]Ϗ�L*�  D.cLT0 k� �D�H1d�'Qe1�t B  ��   � <�8O�5@�4\t   AQ�A���^�3A]ˏ�L*�  D.cLT0 k� �<�@1d�'Qe1�t B  �� 
  � <�8O�5@�4\t   AQ�A���^�3A]ˏ�L*  D.cLT0 k� �8�<1d�'Qe1�t B  �� 
  � <�8O�4@�4\t   AQ�A���^�3A]Ǐ�L)  @/cHT0 k� �8�<1d�'Qe1�t B  �� 
  � <�8O�4@�4\p   AQ�A���^�3A]Ǐ�L)  @/cHT0 k� �8�<1d�'Qe1�t B  �� 
  � <�8O�4@�8\p!  AQ�A���^�3A]Ï�L)  @/cHT0 k� �<�@1d�'Qe1�t B  �� 
  � <�8O�4@�8\p!  AQ�A!���^�3A]Î�L)$  @/cHT0 k� �@�D1d�'Qe1�t B  �� 
  � <�8O�4@�8\l!  AQ�A!���^�3A]���L)�,! </cHT0 k� �H�L1d�'Qe1�t B  �� 
  � <�8O�3@�8\l!  AQ�A!���^�3A]���L(�4! </Z�HT0 k� �P�T1d�'Qe1�t B  �� 
  � <�8O�3@�8\l"  AQ�A!���^�3A]���L(�<! </Z�HT0 k� �X�\1d�'Qe1�t B  �� 
  � <�8O�3@�8\l"  AQ�A!���^�3A]���L(�D! </Z�HT0 k� �`�d1d�'Qe1�t B  �� 
  � <�8O�3@�8\h"  AQ�A!���^�3A]���L(�L! 8/Z�HT0 k� �h�l1d�'Qe1�t B  �� 
  � <�8O�3@�8\h"  AQ�A!���^�3A]���L(�T  8/Z�HT0 k� �p�t1d�'Qe1�t B  �� 
  � <�8O�2@�8\h"  AQ�A!���^�3A]���L(�\  8/Z�HT0 k� �x�|1d�'Qe1�t B  �� 
  � <�8O�2@�8\h#  AQ�A!���^�4A]���L'�d  8/Z�HT0 k� ��
��
1d�'Qe1�t B  �� 
  � <�8O�2@�<\d#  AQ�A!���^�4A]���L'�l  4/Z�HT0 k� ����1d�'Qe1�t B  �� 
  � <�8O�2@�<\d#  AQ�A!���^�4A]���L'�t  4/Z�HT0 k� ����1d�'Qe1�t B  �� 
  � <�8O�2@�<\d#  AQ�A���^�4A]���L'�| 4/Z�HT0 k� ����1d�'Qe1�t B  �� 
  � <�8O�1@�<\d#  AQ�A���^�4A]���L'� 4/Z�DT0 k� ��
��
1d�'Qe1�t B  �� 	  � <�8O�1@�<\d#  AQ�A���^�4A]���L'� 0/cDT0 k� ��
��
1d�'Qe1�t B  �� 	  � <�8O�1@�<\d#  AQ�A���^�4A]���L'� 0/cDT0 k� ��
��
1d�'Qe1�t B  �� 	  � <�8O�1@�<\d#  AQ�A���^�4A]���L&ޜ 0/cDT0 k� ��
��
1d�'Qe1�t B  �� 	  � <�8O�1@�<\d#  AQ�A���^�4A]���L&ޠ 0/cDT0 k� ��
��
1d�'Qe1�t B  �� 	  � <�8O�1@�<
\d#  AQ�A���^�4A]���L&ި ,/cDT0 k� ��
��
1d�'Qe1�t B  �� 	  � <�8O�0@�<
\`#  AQ�A���^�4A]���L&ް ,/cDT0 k� ��	��	1d�'Qe1�t B  �� 	  � <�8O�0@�<
\`#  AQ�A���^�4A]���L&޸ ,0cDT0 k� ��	��	1d�'Qe1�t B  �� 	  � <�8O�0@�@	\`$  AQ�A���^�4A]���L&μ ,0cDT0 k� ��	��	1d�'Qe1�t B  �� 	  � <�8O�0@�@	\`$  AQ�A���^�4A]���L&�� ,0cDT0 k� ��	��	1d�'Qe1�t B  �� 	  � <�8O�0@�@	\`$  AQ�A!���^�4A]���L&�� (0cDT0 k� ��	��	1d�'Qe1�t B  �� 	  � <�8O�0@�@	\`$  AQ|A!���^�4A]���L%�� (0cDT0 k� ��	��	1d�'Qe1�t B  �� 	  � <�8O�0@�@\\$  AQ|A!���^�4A]���L%�� (0Z�DT0 k� ����1d�'Qe1�t B  �� 	  � <�8O�/@�@\\$  AQ|A!���^�4A]���L%�� (0Z�DT0 k� ����1d�'Qe1�t B  �� 	  � <�8O�/@�@\\$  AQ|A!���^�4A]���L%�� $0Z�DT0 k� ����1d�'Qe1�t B  �� 	  � <�8O�/@�@\\$  AQ|A!���^�4A]���L%�� $0Z�DT0 k� ��� 1d�'Qe1�t B  �� 	  � <�8O�/@�@\\$  AQxA!���^�5A]���L%�� $0Z�DT0 k� � �1d�'Qe1�t B  �� 	  � <�8O�/@�@\\%  AQxA!���^�5A]���L%�� $0Z�DT0 k� ��1d�'Qe1�t B  ��   � <�8O�/@�@\X%  AQxA!���^�5A]���L%�� $0Z�DT0 k� ��1d�'Qe1�t B  ��   � <�8O�/@�@\X%  AQxA!���^�5A]���L%�  0Z�@T0 k� ��1d�'Qe1�t B  ��   � <�8O�/@�@\X%  AQtA!���^�5A]���L$�  0Z�@T0 k� ��1d�'Qe1�t B  ��   � <�8O�.@�@\X%  AQtA���^�5A]���L$�  0Z�@T0 k� � �$1d�'Qe1�t B  ��   � <�8O�.@�D\X%  AQtA���^�5A]���L$�  0Z�@T0 k� �$�(1d�'Qe1�t B  ��   � <�8O�.@�D\X%  AQtA���^�5A]���L$�  1Z�@T0 k� �(�,1d�'Qe1�t B  ��   � <�8O�.@�D\X%  AQtA���^�5A]���L$�   1Z�@T0 k� �,�01d�'Qe1�t B  ��   � <�8O�.@�D\X%  AQtA���^�5A]���L$�$ 1Z�@T0 k� �0�41d�'Qe1�t B  ��   � <�8O�.@�D\T&  AQpA���^�5A]���L$�( 1Z�@T0 k� �8�<1d�'Qe1�t B  ��   � <�8O�.@�D\T&  AQpA���^�5A]���L$�0 1Z�@T0 k� �H�L1d�'Qe1�t B �   � <�8O�.@�D\T&  AQpA���^�5A]���L$�4 1Z�@T0 k� �X�\1d�'Qe1�t B ��   � <�8O�.@�D\T&  AQpA���^�5A]���L$�8 1Z�@T0 k� �h�l1d�'Qe1�t B ��   � <�8O�-@�D\T&  AQpA���^�5A]���L#�< 1Z�@T0 k� �{���1d�'Qe1�t B ��   � <�8O�-@�D\T&  AQlA���^�5A]���L#�@ 1Z�@T0 k� ������1d�'Qe1�t B ��   � <�8O�-@�D\T&  AQlA���^�5A]���H#�H 1Z�@T0 k� ������1d�'Qe1�t B ��   � <�8O�-@�D\T&  AQlA���^�5A]���H#	L 1Z�@T0 k� ������1d�'Qe1�t B	 ��   � <�8O�-@�D\P&  AQlA���^�5A]���H#	P 1Z�@T0 k� ������1d�'Qe1�t B
 ��   � <�8O�-@�D\P&  AQlA���^�5A]���H#	T 1Z�@T0 k� ������1d�'Qe1�t B ��   � <�8O�-@�D\P&  AQlA���^�5A]���H#	X 1Z�@T0 k� ������1d�'Qe1�t B ��   � <�8O�-@�D\P&  AQhA���^�5A]���H#	\ 1Z�@T0 k� ������1d�'Qe1�t B ��   � <�8O�-@�D\P'  AQhA���^�5A]���H#	` 1Z�@T0 k� �����1d�'Qe1�t B ��   � <�8O�-@�D\P'  AQhA���^�5A]���H#	d 1Z�@T0 k� ����1d�'Qe1�t B ��   � <�8O�,@�H\P'  AQhA���^�5A]��H#	h 1Z�@T0 k� �#��'�1d�'Qe1�t B ��   � <�8O�,@�H\P'  AQhA���^�5A]��H#	l 1Z�@T0 k� �3��7�1d�'Qe1�t B ��   � <�8O�,@�H\P'  AQhA���^�5A]��H#	p 1Z�@T0 k� �C��G�1d�'Qe1�t B ��   � <�8O�,@�H\P'  AQhA���^�6A]��H"	t 1Z�@T0 k� �S��W�1d�'Qe1�t B ��   � <�8O�,@�H\L'  AQdA���^�6A]��H"	x 2Z�@T0 k� �c��g�1d�'Qe1�t B ��   � <�8O�,@�H\L'  AQdA���^�6A]{��H"	| 2Z�@T0 k� �w��{�1d�'Qe1�t B ��   � <�8O�,@�H\L'  AQdA���^�6A]{��H"	� 2Z�@T0 k� ������1d�'Qe1�t B ��   � <�8O�,@�H\L'  AQdA���^�6A]{��H"	� 2Z�@T0 k� ������1d�'Qe1�t B ��   � <�8O�,@�H\L'  AQdA���^�6A]{��H"	� 2Z�@T0 k� ������1d�'Qe1�t B ��   � <�8O�,@�H\L'  AQdA���^�6A]{��H"	� 2Z�@T0 k� ������1d�'Qe1�t B ��   � <�8O�,@�H \L'  AQdA���^�6A]{��H"	� 2Z�@T0 k� ������1d�'Qe1�t B ��   � <�8O�,@�H \L(  AQdA���^�6A]w��H"	� 2Z�<T0 k� ������1d�'Qe1�t B ��   � <�8O�,@�H \L(  AQ`A���^�6A]w��H"	� 2Z�<T0 k� ������1d�'Qe1�t B ��   � <�8O�+@�H \L(  AQ`A���^�6A]w��H"	� 2Z�<T0 k� ������1d�'Qe1�t B ��   � <�8O�+@�H \L(  AQ`A���^�6A]w��H"O� 2Z�<T0 k� ����1d�'Qe1�t B ��   � <�8O�+@�H \H(  AQ`A���^�6A]w��H"O� 2Z�<T0 k� ����1d�'Qe1�t B ��   � <�8O�+@�H \H(  AQ`A���^�6A]w��H"O� 2Z�<T0 k� �+��/�1d�'Qe1�t B  ��   � <�8O�+@�K�\H(  AQ`A���^�6A]s��H"O� 2Z�<T0 k� �?��C�1d�'Qe1�t B  ��   � <�8O�+@�K�\H(  AQ`A���^�6A]s��H"O� 2Z�<T0 k� �O��S�1d�'Qe1�t B! ��   � <�8O�+@�K�\H(  AQ`A���^�6A]s��H"O� 2Z�<T0 k� �_��c�1d�'Qe1�t B" ��   � <�8O�+@�K�\H(  AQ`A���^�6A]s��H!O� 2Z�<T0 k� �o��s�1d�'Qe1�t B" ��   � <�8O�+@�K�\H(  AQ\A���^�6A]s��H!O� 2Z�<T0 k� �����1d�'Qe1�t B# ��   � <�8O�+@�O�\H(  AQ\A���^�6A]s��H!O� 2Z�<T0 k� ������1d�'Qe1�t B# ��   � <�8O�+@�O�\H(  AQ\A���^�6A]s��H!O� 2Z�<T0 k� ������1d�'Qe1�t B$ ��   � <�8O�+@�O�\H(  AQ\A���^�6A]o��H!O� 2Z�<T0 k� ������1d�'Qe1�t B$ ��   � <�8O�+@�O�\H(  AQ\A���^�6A]o��H!O� 2Z�<T0 k� �þ�Ǿ1d�'Qe1�t B% ��   � <�8O�+@�O�\H(  AQ\A���^�6A]o��H!O� 2Z�<T0 k� �Ӽ�׼1d�'Qe1�t B% ��   � <�8O�+@�O�\H(  AQ\A���^�6A]o��H!O� 2Z�<T0 k� ����1d�'Qe1�t B& ��   � <�8O�+@�O�\H)  AQ\A���^�6A]o��H!O� 2Z�<T0 k� �����1d�'Qe1�t B& ��   � <�8O�*@�O�\H)  AQ\A���^�6A]o��H!O� 2Z�<T0 k� ����1d�'Qe1�t B& ��   � <�8O�*@�O�\D)  AQ\A���^�6A]o��H!O� 2Z�<T0 k� ����1d�'Qe1�t B' ��   � <�8O�*@�O�\D)  AQXA���^�6A]o��H!O� 2Z�<T0 k� �'��+�1d�'Qe1�t B' ��   � <�8O�*@�O�\D)  AQXA���^�6A]k��H!O� 2Z�<T0 k� �7��;�1d�'Qe1�t B' ��   � <�8O�*@�O�\D)  AQXA���^�6A]k��H!O� 3Z�<T0 k� �G��K�1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQXA���^�6A]k��H!O� 3Z�<T0 k� �W��[�1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQXA���^�6A]k��H!O� 3Z�<T0 k� �k��o�1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQXA���^�6A]k��H!O� 3Z�<T0 k� �{���1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQXA���^�6A]k��H!O� 3Z�<T0 k� ������1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQXA���^�6A]k��H!O� 3Z�<T0 k� ������1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQXA���^�6A]k��H!O� 3Z�<T0 k� ������1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQXA���^�6A]k��H!O� 3Z�<T0 k� ������1d�'Qe1�t B) ��   � <�8O�*@�O�\D)  AQXA���^�7A]g��H!O� 3Z�<T0 k� �ˠ�Ϡ1d�'Qe1�t B) ��   � <�8O�*@�O�\D)  AQXA���^�7A]g��H!O� 3Z�<T0 k� �ߞ��1d�'Qe1�t B) ��   � <�8O�*@�O�\D)  AQXA���^�7A]g��H!O� 3Z�<T0 k� ����1d�'Qe1�t B) ��   � <�8O�*@�O�\D)  AQTA���^�7A]g��H!O� 3Z�<T0 k� �����1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQTA���^�7A]g��H O� 3Z�<T0 k� ����1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQTA���^�7A]g��H O� 3Z�<T0 k� ���#�1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQTA���^�7A]g��H O� 3Z�<T0 k� �/��3�1d�'Qe1�t B( ��   � <�8O�*@�O�\D)  AQTA���^�7A]g��H O� 3Z�<T0 k� �C��G�1d�'Qe1�t B( ��   � <�8O�*@�O�\D*  AQTA���^�7A]g��H O� 3Z�<T0 k� �S��W�1d�'Qe1�t B( ��   � <�8O�*@�O�\@*  AQTA���^�7A]g��H O� 3Z�<T0 k� �c��g�1d�'Qe1�t B( ��   � <�8O�*@�O�\@*  AQTA���^�7A]g��H O� 3Z�<T0 k� �s��w�1d�'Qe1�t B' ��   � <�8O�*@�O�\@*  AQTA���^�7A]c��H O� 3Z�<T0 k� ������1d�'Qe1�t B' ��   � <�8%S��CB�_ �#�  E���3� ��D�G�b�%!, ǊZ<8T0 k� �\�`1d�'Qe1�t B  ��/ 
  ��� �%S��CB�^ ��  E���3���D�C�b�%!- ËZ<8T0 k� �`�d1d�'Qe1�t B  ��/ 
  ��� �%S��CB�] ��  E���3���D�C�b�%!. ��Z<8T0 k� �h�l1d�'Qe1�t B  ��/ 
  ��� �%S��CR�] ��  E���3���D�?�b�%!/ ��Z<8T0 k� �l �p 1d�'Qe1�t B  ��/ 	  ��� �%S��CR�\ ��  E���3���E�;�b�%!1�Z<8T0 k� �p$�t$1d�'Qe1�t B  ��/ 	  ��� �%S��CR�[ ��  E���3���E�7�b�%2�Z<8T0 k� �t(�x(1d�'Qe1�t B  ��/ 	  ��� �%S��CR�Z ��  E���3���E�3�b�%3�Z<8T0 k� �x,�|,1d�'Qe1�t B  �_ 	  ��� �%S��CR�YC�  E���3���E�3�b�%4�Z<8T0 k� �+��+1d�'Qe1�t B  ��_ 	  ��� �%S��CR�XC�  E���3���E�+�b�%6�Z<8T0 k� �(��(1d�'Qe1�t B ��_ 	  ��� �%S��CR�WC�  E���3���F'�R�%7�Z<8T0 k� ��'��'1d�'Qe1�t B ��_ 	  ��� �%S��CR�VC�  E�� 3���F'�R�%8�Z<8T0 k� ��%��%1d�'Qe1�t B ��_ 	  ��� �%S��E2�UC�  E��3���F#�R�%9 ��Z<8T0 k� ��$��$1d�'Qe1�t B ��_ 	  ��� �%S��E2�SC�  E��3���F#�R�%: ��Z<8T0 k� �#�#1d�'Qe1�t B ��_ 	  ��� �%S��E2�RB��  DҐ3�	��F�R�%�; ��Z<8T0 k� �"�"1d�'Qe1�t B ��_ 	  ��� �%S��E2�QB��  DҐ3�	��Es�B�%�< ��Z<8T0 k� �, �0 1d�'Qe1�t B ��_ 	  ��� �C��E2�PB��  DҐ�
��Es�B�%�= ��Z<8T0 k� �@�D1d�'Qe1�t B ��_   ��� �C��E2�OB��  DҔ���Es�B�%� = ��Z<8T0 k� �P�T1d�'Qe1�t B ��_   ��� �C��E2�MB��  DҔ���Es�B�%� > ��Z<8T0 k� �d�h1d�'Qe1�t B ��_   ��� �C��E2�LR��  DҔ���Es�B�%�$? ��Z<8T0 k� �x�|1d�'Qe1�t B ��_   ��� �C��E2�KR�  DҘ	���Es�B�%�(? ��Z<8T0 k� ���1d�'Qe1�t B ��_   ��� �C��E2�IR�  DҘ
���Es�B�%�,@��Z<8T0 k� ���1d�'Qe1�t B ��_   ��� �C��CB�HR�  DҜ���Es�B�%�,@��Z<8T0 k� ���1d�'Qe1�t B $�_   ��� �C��CB�GR�  DҜ�� F�B�%�0A��Z<8T0 k� ���1d�'Qe1�t B ��_   ��� �C��CB�ER�  DҠ��F�B�%�4A��Z<8T0 k� ���1d�'Qe1�t B ��_   ��� �C��CB�DR�  DҠ��F�B�%�8B��Z<8T0 k� ���1d�'Qe1�t B ��_   ��� �ë�CB�BR�  D���F�B�%�<B���Z<8T0 k� ���1d�'Qe1�t B ��_   ��� �ë�CB�@R�  D���F�B�%�@B���Z<8T0 k� ���1d�'Qe1�t B ��_   ��� �ë�CB�=R�  D���F�B�%�HC���Z<8T0 k� Ө��1d�'Qe1�t B ��_   ��� �ç�CB�;b�  D���	F�B�%�LC���Z<8T0 k� Ө��1d�'Qe1�t B ��_   ��� �ç�CB�:bߨ  E����F�B�%�PC���Z<8T0 k� Ө��1d�'Qe1�t B ��_   ��� �ç�CB�8bߩ  E����F�B�%�TC���Z<8T0 k� Ӥ��1d�'Qe1�t B ��_   ��� �ç�CB�6b۪  E���"D��B�%�XC���Z<8T0 k� Ө��1d�'Qe1�t B ��U   ��� �ç�CR�6b۬  E��s�"D���%�\C���Z<8T0 k� ����1d�'Qe1�t B ��U   ��� �ç�CR�6�ۭ  E��s�" D���%�`C���Z<8T0 k� ����1d�'Qe1�t B ��U   ��� ����CR�5�׮  E��s�" D���$�hC���Z<8T0 k� ����1d�'Qe1�t B ��U   ��� ����CR�5�ӱ  E��s�"(D���#�pB���Z<8T0 k� ����1d�'Qe1�t B ��U   ��� ����E��4�Ӳ  E����",D��Ҍ"�tB���Z<8T0 k� Ӥ��1d�'Qe1�t B ��U   ��� ����E��4�Ӵ  I���",D��Ҍ!�|B���Z<8T0 k� Ӭ��1d�'Qe1�t B  ��U   ��� ����E��3�ϵ  I���"0D��҈!��A���Z<8T0 k� Ӵ��1d�'Qe1�t B  ��U   ��� ����E��2�Ϸ  I� ��"4D��҈ ��A���Z<8T0 k� Ӹ
��
1d�'Qe1�t B  .�U   ��� ����E2�˺  I�!��"<E��҄��@���Z<8T0 k� ���1d�'Qe1�t B  ��U   ��� ����E2�ǻ  I�"��@!E�����@���Z<8T0 k� ���1d�'Qe1�t B  ��U   ��� ����E1�ǽ  I"�"��@!E�����?���Z<8T0 k� ���1d�'Qe1�t B  ��U   ��� ����E0�þ  I"�#��@#E���|��>���Z<8T0 k� ���1d�'Qe1�t B  ��U   ��� ����E/���  I"�#��D%E���|��>���Z<8T0 k� ���1d�'Qe1�t B ��U   ��� ����EҀ-»�  I"�$s�D%E�#��xq�=���Z<8T0 k� ���1d�'Qe1�t B ��U   ��� ����EҀ-»�  I�%s�D&E�'��xq�<���Z<8T0 k� �
��
1d�'Qe1�t B ��U   ��� ���EҀ,���  I %s�@&E�+��tq�;���Z<8T0 k� ���1d�'Qe1�t B ��U   ��� �3�EҀ,���  I&s�@'F/��tq�:���Z<8T0 k� ���1d�'Qe1�t B ��U   ��� �3w�EҀ+���  I's��@)F3��l�8���Z<8T0 k� Ø��1d�'Qe1�t B  ��U   ��� �3s�EҀ*���  E�'s��@)F7��l�8���Z<8T0 k� Ô��1d�'Qe1�t B  ��U   ��� �3s�EҀ*���  E�(s��@)F8�h�7���Z<8T0 k� Ð��1d�'Qe1�t B  ��U   ��� �3o�EҀ*���  E�(s��@)F<�d�6���Z<8T0 k� Ð��1d�'Qe1�t B  ��U   ��� �3k�EҀ*���  E�)s��@)F@�`�4���Z<8T0 k� Ì��1d�'Qe1�t B  ��U   ��� �3g�C�*���  Es+���@+FH	�Xq�2���Z<8T0 k� ���1d�'Qe1�t B  ��U   ��� �Cc�C�)���  Es +���@,FL�Tq�1���Z<8T0 k� ���1d�'Qe1�t B  ��U   ��� �C_�C�)���  Es$,���@-FP�Pr 0���Z<8T0 k� ���1d�'Qe1�t B  ��U   ��� �C_�C�(���  Es(-���@-E�T�Hr 0���Z<8T0 k� |��1d�'Qe1�t B  ��U   ��� �CW�C�'���  Es,/���D/E�\�@r.���Z<8T0 k� �x�|1d�'Qe1�t B  ��U   ��� ��S�C�|'���  Es0/��D/E�`�<r-���Z<8T0 k� �t�x1d�'Qe1�t B  ��U   ��� ��O�C�|&��  Es00��H0E�d4r,���Z<8T0 k� �p
�t
1d�'Qe1�t B  ��U   ��� ��O�C�|&�{�  Es40��H1E�h0r+���Z<8T0 k� �p
�t
1d�'Qe1�t B  ��U   ��� ��G�C�x%�s�  Es82��P2E�p$
b)���Z<8T0 k� �h
�l
1d�'Qe1�t B  ��U   ��� ��C�C�x$�o�  Es82��T3E�t	b'���Z<8T0 k� �`�d1d�'Qe1�t B  ��U   ��� ��?�C�x#�k�  Es<3��T3E�xb&���Z<8T0 k� �X�\1d�'Qe1�t B  ��U   ��� ��;�C�t#�g�  Es<3��
X4E�� b%���Z<8T0 k� �P�T1d�'Qe1�t B  ��U   ��� ��3�C�p"�_�  Es@4��
�`5E��#b"���Z<8T0 k� �H�L1d�'Qe1�t B  ��U   ��� ��/�C�l!�[�  Es@4Ӏ
�d6E��$�b!���Z<8T0 k� �O��S�1d�'Qe1�t B  ��U   ��� ��+�E�l!�W�  Es@4�x
�h6E��%�b  ���Z<8T0 k� �O��S�1d�'Qe1�t B  ��U   ��� ��'�E�h �S�  EsD5�t	�p7E��&�b ���Z<8T0 k� �K��O�1d�'Qe1�t B  ��U   ��� ���E�`�K�  EsD5�l	�x7E��(�b ���Z<8T0 k� �3��7�1d�'Qe1�t B  �U   ��� ���E�`�G�  EsD5�h�|7E��)�b 	���Z<8T0 k� ���#�1d�'Qe1�t B  ��    ��� ���E�`�C�  EsD5�dҀ8E��)�b 	���Z<8T0 k� ����1d�'Qe1�t B  ��    ��� ���E�X�?�  EsD5�\Ҍ8E��+�b 	���Z<8T0 k� ����1d�'Qe1�t B  ��    ��� ���E�X�8   EsD5�XҐ8E��+�R	���Z<8T0 k� �����1d�'Qe1�t B  ��    ��� ���E�T�4  EsD5�TҘ8E��,� R	���Z<8T0 k� ������1d�'Qe1�t B  ��    ��� �                                                                                                                                                                            � � �  �  �  c A�  �J����  �     6 \���� ]�&x&x   � **   $ N     ����     *
���ٺ    �| }             	 
   X           ��     ��    0

         ����          ��S��    �����S�    �� l   	                        �      ��   0           *'          ��     *���P     ��e   
          
  �         ?0     ��    8
	          ���         qs    ���  qs           
    ��       		 ���          �       ��   0	          A\s          . Ul�     A\s U|�      �              
 A c          <�     ��    8	
'	           ����  ��	      B ��    ���� ��                            ��]             �  ��     		 5             78�          V����     73�����     H��               3 �         �     ���   0

          ��"�  T     j�X�5    ��#*�Y	�    ����                � ��        ��     ���   (
            ��         ~�R�+      ��R�+    ��               �          �     ���   8�		          �q  $ �       �����     �V��L�    �k�               �n         	 ��      ���   (
            3�c           ��o     3��*P     `�/              
   �$         
  �`     ���   PB           `���
     ��hE     `��j�      ��                    ���8             �  ���    8		 1 	                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         ����  ��        � ��" '����iT ܜ� '�@��>��                x                j  �  �	   �                         ��    ��       � �      ��   �           "                                                 �                          *�� *� A�� 7��    3     ����          
 	      
       � �\ ���O       �� �e� �� f�  s����  ����. ����< ����J ����X � GD ``� H 0a� Hd a� H� b ���� ���� ���� ����  ����. ����< ����J ����X � 
� W� 
�< W� 
�\ W� �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  
�\ U� 
�� V  
�| V ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����8�� <      ������  
�fD
��L���"����D" � j  "  B   J jF�"     
�j,
 ��
��
��"    B�j l �  B �
� �  �  
�  ��  ��     ���  �   ��    ��     ��S       ��  ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �      ��" �  ���        � � �  ��        �        ��        �        ��        � 	 	  �    �z 
����        ��                         T�) , � ���                                     �                ����          
  	 ��	���%��   <�8�� F��            6BUF  Housley v      0:55                                                                        4  4     �icVX� c^`_K. � K6 �BS �" � �!� � � *8# 	C � �
c~ � � c� � �J� � � J� � scV � � c^ � �"� � � "� � �"� � �*� � �*l � *Fd �*8d �)�d *Fd*l0*
lP  *CT [� � [
� � �*l � *Fd � *8d �!)�d "*Fd#*l0$*
lP  *CTP  *CTP  *CTP  *CT8 )*DLX  *K<8 +*ILX  *H<Y  *H<A  *IL z /"�> j0�( j 
�7 � 
�8 � 
�7 s  "O u �5
�4 w  "O u |  "O u �8*4= �  *N] �  *N]P ;"R �X  "K � z="4 � >*T �  *Nl                                                                                                                                                                                                                           � p       �     @ 
        j     Y P E ^  ��        	            �������������������������������������� ���������	�
��������                                                                                          �� 
 ��� � ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   ��, 1  * ��� :� A� �� ��@�� �@��                                                                                                                                                                                                                                                                                                                               @�                                                                                                                                                                                                                                             	       �        ��   K
�J     �b  	                           ���������������������������������� 7����������������"�                                                                                                                                         C  Y                 Y      Y   A          	 	 
  	 
 
 ����������� ����� ���� ������������� ���������������� ������������������������� �� �����������������������  � ���������� ������ �� ��� ����������������� ������������ �����������������������������������������������                                    �          �  L�J      Q                             �����������������������������������������������������                                                                       	                                                                     Y    YY              Y          YY                 	 	  ��������������������������� ����������� ������ ���� ����������� ������ � �������� ������������� �� �� ��� ������������ � ��� ������� ���������������� ����������������������  ����� �� �������� ������������������ � ��             A                                                                                                                                                                                                                                       	                                                                    �             


             �   }�         �#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" > D 6                                 � �?�E �e�                                                                                                                                                                                                                                                                                    E)n1n  �                c            `            d                                                                                                                                                                                                                                                                                                                                                                                                                            � � �  � ��  � ��  � 2��  � 2��  � ��  �����}������������������������������������&                       �          �   & AG� �  x   
              �                                                                                                                                                                                                                                                                                                                                        F I   �                     !��                                                                                                                                                                                                                            Y    �� �~ ��      �� Z      ����������� ����� ���� ������������� ���������������� ������������������������� �� �����������������������  � ���������� ������ �� ��� ����������������� ������������ ����������������������������������������������� ��������������������������� ����������� ������ ���� ����������� ������ � �������� ������������� �� �� ��� ������������ � ��� ������� ���������������� ����������������������  ����� �� �������� ������������������ � ��             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    '      &     ��                       f     � ' �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$ ^h  ��  p    �f ��    �f �$ ^$ �@      �       �     �  v 
� � v                   x       �  �   �      7        �   ��    �   �$ ^$         �      � ��     � �$ ^$  &x   x x        �  �            �   ���          H     }PS   yL  ��������������������������������GvdDGw6wGwcfGwsfGwv6Gww6GwwcGwwcDDDDwwwwffffffffffffffffUUUUttttDDDDwwwwffffffffffffffffUUUUtttwN���t���wN��wt��wwN�wwt�wwwNwwwtGwweGwwU�tvf�wff�Fff�Fff��df��ffwwwwUUUUffffftDDft33gt5egt6Vgt5gwwwwUUUUffffDDDD3333eeeeVVVVwwwwwwwwUUUUffffDDFF35FfefDDVVFUufGfwwwwGwwwGwwwUUUUffffDDDDUUUUffffwwwwwwwuwwwuUUUUffffDDDDUUUUffffwwwwUUUUffffddDDfd33DD6VUd5eft6WwwwwUUUUffffDDGf35GfVVGvefGv6VGvwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwN�Fft�FfwN�dwt�fwwNGwwtGwwwDwwwtwt6Wwt5gwt6Wwt5gwt6Wwt5gtt6Wwt5gDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD6VGd5fGd6VGd5fGd6VGd5fGd6VGd5fGdFt5gFt6WFt5gFt6WFt5gFt6WFt5gFt6W5fGw6VGw5fGw6VGw5fGw6VGw5fGG6VGwgwwwvwwwwgwwwvwwwwgwwwvwwwwgwwwvGt6WGt5gDt6WDt5gND6WNt5gNt6WNt5g6VGd5fGf6VGw5fDD6VGU5fGf6VGf5fGfDDDDffffwwwwDDDDUUUUffffffffffffFt5gft6Wwt5gDD6WUt5gft6Wft5gft6W5fGt6VGt5fGD6VGD5fD�6VG�5fG�6VG�GwwwDwww�Gww�Dww~�Gww�Dww�DGw~�DNt6SNt5fNt6VNteeNwFVNwteNwwFfffd3333ffffVVVVeeeeVVVVeeeeffffDDDD333DffcDVVSDeecDVVSDeecDfVSDFecDUUUUDDDDDDDDDDDDDDDDDDDDDDDDDDDDD333D6ffD6VVD5fdD6VDD5fDD6VDD5fD3333ffffVVVVDDDD33335UUU5Vff5VDD3333ffffVVVVDDDD3333UUUUffffDDDD6VGfefGfVVGwDDDD3333UUUUffffDDDDffffffffwwwwDDDD3333UUUUffffDDDDft5cft6Vwt5eDDDD3333UUUUffffDDDD3333ffffeeeeDDDD3333UUUVffeVDD5V333DffcDeecDF6SDD5cDD6SDD5cDD6SDD333D6ffD5eeD6VVD5eeD6VVD5ffD6Vd5fG�fVG�efG�VVG�edw�VGw�dww�Ffffffffwwwwwwww����DDDDNNDD��������gwwwwwwwwwww��wwDDGwDDDw��DG���Dwwwwwwwwwwwww~��wwn�wwvwwwwgwwwvFfffFfffCeeeCVVVCeeeCVVVCeeeCVVVfDDDfDDDfDDDVDDDfDDDVDDDfDDDVDDDDfSDD5cDD6SDD5cDD6SDD5cDD6SDD5cDD6VDD5fDD6VDD5fDD6VDD5fDD6VDD5fD5VDD5VDD5VDD5VDD5VDD5VDD5VDD5VDDDDDDDDDADDDADDDDDDDDDDDADDDADDDDDDDDDDDDDDwDDDDDDDDDDDDDwDDDDD5VDD5VDD5VDD5VDD5VDD5VDD5VDD5VD5cDD6SDD5cDD6SDD5cDD6SDD5cDD6SDDDDfDDDfDDD5DDD6DDD5DDD6DDD5DDD6fffdfffdeeedVVVdeeedVVVdeeedVVVdCeeeCVVVCeeeCVVVCeeeCVVVCeeeCVVVfDDDVDDDfDDDVDDDfDDDVDDDfDDDVDDDD6SDD5c3D6VfD5eeD6VVDVffDDDDDDDDDDDD3333ffffeeeeVVVVffffDDDDDDDDD6VD35fDffVDeefDVVVDfffDDDDDDDDD5VDD5VDD5V335UUU5UUU5UUUVfffDDDDDDDDDDDD3333UUUUUUUUUUUUffffDDDDDD5VDD5V335VUUUVUUUVUUUVffffDDDDD5cDD6S3D5ffD6VVD5eeD6ffDDDDDDDDD5fD36VDfefDVVVDeefDfffDDDDDDDDDDDD5DDD6DDD5DDD6DDD5DDD6DDD5DDD6eeedVVVdeeedVVVdeeedVVVdeeedVVVdwwww�twwww~ww�w�wtwwtwwww~w�wwwwDDDDDDDDDADDDDDADDDDDDDDDDDtDD4DDqt4DDDD4DDsDDDDDDDDDDDD7AtCADADDADADDDDDDDADDDADDADqDADqDDDDDADDDADDDAADAADqADDAGADDDDwwwywww�www�www�www�www�www�www�������������������������www�www�www�www�www�www�www�www����������������������!�����!�-����������!-�����������!�����wwwwwwwtwwwOwww�wwt�ww�wwOGww�D��������������-��������������������������!����������-������NNNNNNNNNNNNN���FfwfDDDDDDDDDDDDNNNDNNNDNNND����gvftDDDDDDDDDDDDwts"wwB2ww22ws#Cws#4ww2twws�www�www�www�www�www�www�www�wwwywwww��������wwww������!��������wwwwww��w��w2��w���w��t���(�wy���������y���w�����y��Gwwwwt33Dt343CeeeCVVVEeeetVVVvEee�DVVzDFf�DDDfDDDVDDDe333VfffeeeeVVVVffffDDDDDDDDDDDD3333ffffeeeeVVVVffffDDDDDDD5DDD6333efffVeeeeVVVVffffDDDDeeedVVVdeeedVVVGeedgVVDzfdD�DDD�Df��NvDGN�DNN�DND~DGD��NDNt�DDDN#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFw"GC42wsDCwt�Cwt��ws�DGt�T7DfEGt{�Gwz��w���wt�Gw��wt�Gw�wtw�{�Gww��w��w2��w���w��w���x�wy����wwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wt3Gwt4wCGGttwG4�twO�wGt�GwE��wTfNw~D�����������������DD��ww�N��D�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wfuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGy�wwy�wtw�wOw�w�w�D�w2?�wCOGww�Dwwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGww23ws""wr22w244w#tD�t3~�}�ww}O3#�w""7w##'wCC#wDG2w3G~������wwwwVtwwUvwwenwwvWwwv�wwtwwtGww�3#�w""7w##'wCC#wDG2w3G~��7���wwww}�ww}�ww}�www�www}www}wwwwwwwr��ww��ww���w4��w��ww��www}ww'r'ww"GCw2wswCwtwCwtw�wswDGtwB'tww"w#w�2w�3w�3wG4wtGDwww"wr!r'wrwuUUG4wwD4wwCtwwCtww7tww7twwGtww8�3�3�3�8�3�3�33333"2#333"33UUUUwwwtwwwtwwwtwwwtwwwtwwwtwwwt��33�?33�?33�?333333#23323#3UUUUwwwwwwwwwwwwwfgvwwwwwwwwwwwwUUUUwwwtwwwtwwwtfwfdwwwtwwwtwwwtUUUUwwwwwwwwwwwwwwwwwwuwwwWwwwwwUUUUwwwWwwwWwwwWwwuwwwuwwUuwwwUwC�38C838C�38C833C332C"33C2#3UUUUwww~www~www~www~www~www~www~UUUUwfwnwvw~wfw~wvw~www~wfw~wgw~UUUUuwwwuwwwuwwwwWwwwWwwwWuwWUwwUUUUwwwwwwwwwwwwwwwwWwwwwwwwwwwwUUUUwwwdwwwdwwwdwwwdwwwdwwwdwwwdUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwUUUVwwwvwwwvwwwvwwwvwwwvwwwvwwwvGtwwGtwwGtwwGtwwGtwwGtwwGtwwGtwwwwwtwwwtwwwtwwwtwwwtwwwtwwwtwwwtww�www�www�www�www�www�www�www�w�www�www�www�www�www�www�www�wwwwwwdwwwdwwwdwwwdwwwdwwwdwwwdwwwdwwwvwwwvwwwvwwwvwwwvwwwvwwwvwwwvGtUUGTffGTffEdffEdffFdffFdffFdffUUUUfffffffffffffffffffffffff���UUUUffffffffffffffffffffffff����UU�Uff�eff�Vff�Vff�fff�fff�fʦ�f�UUU�fff�fff�fff�fff�fff�fff�fffUUUUffffffffffffffffffffffffffffwwwdwwwdd333d333d333d333d333dwwwwwwww33333333333333333333wwwvwwwv33363336333633363336FdffFdffAC333C333C333C333C333��������33333333333333333333�f�f�fFf�33�333�333�333�333�3�fff�fff33333333333333333333ffffffff33333333333333333333333d333d333d333d333d3333����wwww333333333333333333333333����wwww333633363336333633363333����wwwwC333C333C333C333C3333333����wwww33�333�333�333�333�33333����wwww�����<��5UUU5UUSU553SS2#33"532 5�����<��5UUU5UUUU555SSSS33333��������UUUUUUUU5555SSSS3333��������UUU�UU_�55=�SS]�33;������l���eUUUUUUSU552SS2#S3"3S2 0�����<��5UUU5UUSU552SS2#33"332 0����ȩ��S�UUU��US:�U59��38��009������<��UUUUUUUU5555SSSS33333������ÓUUX�UUS�SSX�553�338�003�����3���UUUU5UUUU555SSSS33333�����̚�Ue�5UX�U5Y�5X��S9��3����������UUUUUUUSU5523S2#"302 0�����<��5UUU5UUSU552SS2#33"302 0�����<��5UUV5UUUU555SSSU33353��������UUUUUUUUU5553SSS33330����l���eUUSUUU3SSS%U3"5S2#3S" "#  %                     200            "          "                         0;�  ��  �� ��  ۰  ۰  ��  ��                          #                         P"R                         "#                       "#  "                    0"                                                    �  9                     �#�� ��� ��� ��  �       02(�" �  � ��0(�������� �����   �                    "                         205            "         R 20R                                                                                    ��  ��  �� �� �  �  �  �   �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��  �S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                                  �  � y� ���         ���i���}���������������    �������������������            {  �y�  ˙` ̹� ��i`                                                           	���}���l|���̛��̜�ww�����������qqA}����}q���̙��w���w}w���������w��͝��yq�|�qk}�����ww�    �   {   �     � qy� ��     	   	     �     s�ww���͜���}���}��ww����t��twwwww}q�q|����qwqw}ww���q|����{��wiyww|��{  ِ  y`  ��  �   �   �        ww                            wy�� ��  ��   y              ������������{��̙v��י�  �y    �������������������i���v�w�     �̹p�͙ �ٛ ٗ  ��                   �      �                   wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            "! "   "      ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "                "            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       "! "   "      ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        wݪ 
�� 
�� ��� ��� �̼ �� 	�� 
�� ���"��8�+ӊ"#H�  �E  �T  X�  �   �          "   "   �   ��  ��� ��� �ت �͈ ��� �ː ��� ��@ �U@ �U@ ET  TD  C0  C0  �0  ��  �   �   "/  " � !/  � ���                 �  �˰ ̻� {�ڠ        �  �   �� ��  �      �   �� ��  �"  �            �   �"  ""  !� �� ��  �               �   ������  ��   "   "   "  �� ��                   ����������                �����                      �  �  �   �   ��  �                            �   ���                            �   �                                                                                                                 �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                 �� �̽���ݪ۽w�}�֪�vv���p���      ���� ��                             �    �                    �   �   �                                   ��  ��  ���                    � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                        �          �   � � �  ��� ��  �                    �                        ���� ��� ����                            ��  ��  ���              �  �˰ ��� �wp ���                    �   ���                            �   �    ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r`��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                       � ��                  �  �˰ ��� �wp ���                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                  �   �  "������"    /   �  �   ��                             �                        ���� ��� ����                                    � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                    �  ��  ̽  ��  �w 
�� ���̹����	��̚���ȭ�̻������  ��  H� EU 4E C3  D;  ��  ��  ��  �  �  �   �  "  ��               �   �   �   �   ��  ��� ��� ��� ͻ���ة��ڌ�̽��˽����虚�DD��UT�"DUJ�3ET��DD��4M��ً�������۰��ـ+���+�ۿ��ۏ����"� �    �   �   �   ɀ  ��  ��         �    �  �       �                � ��� ��� ��  �                �   �     �   �           �  ��  ��  ��  ��� ��� ��� ��˰ɜ˰��˻�̻���������3���DDD�                                                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  �   �"  ""  !� �� ��  �               �   ������  ��               �    �                    �   �   �                                   ��  ��  ���   ���� �                                                                                                                                                                                         �� ���
�������˽������̽�]��+I۲"T�""T32.T33>@4C CDT �E@ ��  ʐ  �       "   "�� � ��� �wp ��� �vz �w� �����˻���˰�̰� ��  ��  ��� � �+ �+ �  .   "�   �   �   �    � ��  �                     �  �˰ ���                 ��  ��  ���           U   U  U  U  	T  ,� ,� "  " "  ��  �              �   � � �  ��� ��  �                    �                        ���� ��� ����         �EU �E  
�   �               �"�!/"�  �                                                                                                                                                                                 �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �   �   "   "   "  !�    ��                                 �   �                      �������  ���    �                    ��  ��  ���     ��   �  ��  �  �  �         � �������������  �                                �   �                                                                                                     �  �  �  �  �   �   �  
�  
�  ��  ��  �� 	�� ��� ��������Y� U�  �  �  �  �  ��� �  ��  
   �   "   "     �    �   �   �   �   �   ת� ��� ����������ڀ�̽��̽������̻ �˸ ��� ��C UUC DT3 ES3 ES3 UB� [B"�������� " ��"/�" � "/� � ��                �   �                          ���� ���  ��    �     �  �  ��  �   �                 "��" �"  �"     ��   �          ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                   �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �   �   �   ˰  ˙  ɪ  ��� ټ� �̰ �̰ ��� ��  ��  �   �   ��  �   �   �   �                       �                        ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                             �  ��� ��� ��� �ݪ�                       �   �    �z� 
�� ������������ ˍ� ��� ���������ˉ����� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��                    ˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                                         �  ��  �� ��  �� ���                              �������  �                     �  �   �  �  ��  �  ��  �                                                                                                                                                                                                                �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""���������������������""""������II������""""������IIII""""������DI�I�""""������DI�I�""""�����IIDIIIA""""��������DD""""������IADD�A��""""��������I���I�������I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��                                 � � �� � � � � ����l(�(a(�""""��������AA�A                	 
   ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD   ������� ������� �� ������������   � � � � � � � �����((�l(=LL����������D����3333DDDD   ��	�
��������    ��������������������   ��� � � � � �����((�(( """"����������A������        ����     ! " # # $! % &  ����  ' (����� � � �����(-(5(Xx""""�������I�I������ ) * + , - .  �ڤ�  / 0 � 1 2�� 3 4  �ؤ� / 5 6+*) � � � ��� � �����(�xww""""�������I��D���I�������     7 8 9 : : : : : ; < = = = = = = > ?::::: @ A B     � � � � ��� �����ww�(�D�M�D���M������3333DDDD C CC 7 8 DD  E F G H         DD  E F G H A B CCC �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD    7 8               ��!���%� �  A B   �� � � ��� � ����(W(�m(`""""�����AMAD������   Q 7 8                       A B(Q   � � � � ��� ���	B�(a((M""""������������������ V W X 7 8                       A B(XWV � � � ��� � ���	C�(-(� 
(�fFfFDfFFfFffdFffff3333DDDD V W \ 7 8                       A B(\WV� ���� � � ��	E	D�(( (-(�DDFFDfFFfdFffff3333DDDD V W ] ^ _ ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` a b(]WV��� � � � � ��	F ��(X((6(5""""wwwwwwwGGD V W c d e f g h i j V W  k h i d e f l V W(j m(h(g(f(e(dcWV � � � � � � � ��	G ��l((�x""""wwwwwwqwAqwAwA V W n o p q ] r s t V Wn ] r u o p q v V W(t(s(r(](q(p(onWV���������H������yxww""""wwwwqwqAwAqAqAq V W w f g h i d e f V W x i d e f k h y V W(f(e(d(i(h(g(f(QWV � ��O�N�M�L�K�J�I������w(+�(A�A�A�A��LD�����3333DDDD V W z { ] r u o p q V W | u o p q ] r u V W(q(p(o(u(r(](q }WV�A�A�V�U�T�S�R�Q���P(�((5(U(,�A�LDL�L�D�L�����3333DDDD V W ~  � � � � � � � � � � � � � � � ���(��(��(�(�((~WV�]�]�\�[�Z�Y�X���P(N(,(U((=((+""""wwwwwwDGAD � � � � � � �  �   �  � �� �� �  � �� � � � ���U�U�b�a�`�_���P(U(V(=((( ((5""""wwwwqqDAAq �     � � � � � � � � � � � �����������    ��i�h�g�f�e���P)d((( ((,(U((=""""wwwwwwwGGwGGwGwGw � � � � � � � � � � � � � � � � ����������� � � � ���u�t�s�r�p�p�-(,(N(,(U((=((( UQUUQUUQUUQUUUDUUUUU3333DDDD � � � � � � � � � � � � � � � � � �� � � � � � ��� � � � ��!x!y!z!{!|!}!y!~ � � � � � � � �DEQQUUDUTEUUUU3333DDDD � � � ��� � � � � ��� � � �� � ���� � � � � ���� � �!!�!�!�!�!�!�!� � � � � � � � �""""������������������������ � � � � � � � � � � � � � � � ��� � � � � � � � � � �� � � ��� � � � � � �����(W(�m(`""""�������DAADAI � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqicVX� c^`_K. � K6 �BS �" � �!� � � *8# 	C � �
c~ � � c� � �J� � � J� � scV � � c^ � �"� � � "� � �"� � �*� � �*l � *Fd �*8d �)�d *Fd*l0*
lP  *CT [� � [
� � �*l � *Fd � *8d �!)�d "*Fd#*l0$*
lP  *CTP  *CTP  *CTP  *CT8 )*DLX  *K<8 +*ILX  *H<Y  *H<A  *IL z /"�> j0�( j 
�7 � 
�8 � 
�7 s  "O u �5
�4 w  "O u |  "O u �8*4= �  *N] �  *N]P ;"R �X  "K � z="4 � >*T �  *Nl3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E���������������������������������������������������������������������������������������������������������������������������������������9�K�X�O�U�J���\�K�X����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������,�>�0�	�
�������������������� � � � � � �����������������������������������������%� � ������������������@�9�1� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                