GST@�                                                            \     �                                               �   �                        ����e r�	 J���������������z���        �h     #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    "�j* ,  �����
�"     �j@ �    ��
  �                                                                               ����������������������������������       ��    =b= 0Q0 44 111  4            	 
                    ��� �� � � ��                 nh 	)
         8�����������������������������������������������������������������������������������������������������������������������������?o  0  5o  8    +     '            �  
     
            �	  47  V  �	                  Y            :: �����������������������������������������������������������������������������                                  '       �   @  &   �   �                                                                                 '    	n)h
  Y    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E ' �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    �`A���A�K�L�
���;�C�{�E��l��������3�T0 k� �� �� U8D"!U2d   ��? 
   ����B�aA���A�G�L�	����;�Ds�E��k��������3�T0 k� �p�tU8D"!U2d   ��? 
   ����B�bA���A�C�L�	����;�Do�C��j�������3�T0 k� �\	�`	U8D"!U2d   ��? 
   ����B�cA���A�?�L�	����;�Dg�C��i�������3�T0 k� �H�LU8D"!U2d   ��? 
   ����B�cA���A�;�L�	����;�D_�C��i�������3�T0 k� �4�8U8D"!U2d   ��? 
   ����B�dA���A�7�L�	���;�D[�C��h�������3�T0 k� � �$U8D"!U2d   ��? 
   ����B�eA���A�7�L�	���;�DS�C��g�������3�T0 k� ��U8D"!U2d   ��? 
   ����B�fA���A�3�L�	���;�DK�C��f]� ����3�T0 k� ��!� !U8D"!U2d   ��? 
   ����B�fA��A�/�L����;�DC�C��e]ߘ �� ��3�T0 k� ��%��%U8D"!U2d   ��? 
   ����B�gA��A�+�L����;�D?�C��d]ۘ �� ��3�T0 k� ��*��*U8D"!U2d   ��? 
   ����B|hA�{�A�'�L����;�D7�C��c]ט �� ��3�T0 k� ��/��/U8D"!U2d   ��? 
   ����BxiA�w�A�'�L����;�D/�C��c]ט �� ��3�T0 k� ��3��3U8D"!U2d   ��? 
   ����BpiA�w�A�#�L����;�D'�C��b]Ә �� ��3�T0 k� ��8��8U8D"!U2d   ��? 
   ����BljA�s�A��L����;�D�C��a]Ϙ �� ��3�T0 k� ��=��=U8D"!U2d   ��? 
   ����BhkA�s�A��L����;�D�C��`]Ϙ �� ��3�T0 k� �tA�xAU8D"!U2d   ��? 
   ����B`kA�o�A��L����;�D�C��_]˘ �� ��3�T0 k� �`F�dFU8D"!U2d   (�? 
   ����B\lA�k�A��L����;�D�C��]]ǘ �� ��3�T0 k� +dJ�hJU8D"!U2d   ��?    ����BXmA�k�A��L��#��;�D��C��\]Ø �� ��3�T0 k� +lO�pOU8D"!U2d   ��?    ����BTmA�g�A��L��'��;�D��C��[]Ø�� ��3�T0 k� +pS�tSU8D"!U2d   ��?    ����BLnA�c�A��L��'��;�D�C��Z]���� ��3�T0 k� +tW�xWU8D"!U2d   ��?    ����BHoA�c�A��L��+��;�D�C��Y]���� ��3�T0 k� +|[��[U8D"!U2d   ��?    ����BDoA�_�A��L��+��;�DߧC��X]���� ��3�T0 k� +�`��`U8D"!U2d   ��?    ����B@pA�_�A��L��/��;�DקC��W]���� ��3�T0 k� ��d��dU8D"!U2d   ��?    ����B<qA�[�A��L��3��;�C�ϨC�|V]���� ��3�T0 k� ��g��gU8D"!U2d   ��?    ����B4qA�W�A��L��3��;�C�èC�tT]���� ��3�T0 k� ��k��kU8D"!U2d   ��?    ����B0rA�W�A���L��7��;�C�C�pS]���� ��3�T0 k� ��n��nU8D"!U2d   ��?    ����B,rA�S�A���L��7��;�C�C�lR]��� ��3�T0 k� ��q��qU8D"!U2d   ��?    ����B(sA�S�A���L��;��;�C�C�dQ]��{� ��3�T0 k� ;�t��tU8D"!U2d   ��?    ����B$sA�O�A���L��;��;�C�C�`O]��s� ��3�T0 k� ;�w��wU8D"!U2d   ��?    ����B tA�K�A���L��?��;�I���C�XN]���o� ��3�T0 k� ;�y��yU8D"!U2d   ��?    ����BuA�K�A��L��?��;�I���E>TM]���g� ��3�T0 k� ;�{��{U8D"!U2d   ��?    ����BuA�G�A��L��C��;�I���E>PK]���c� ��3�T0 k� ;�}��}U8D"!U2d   ��?    ����BvA�G�A��L��C��;�I���E>HJ]���[� ��3�T0 k� � �U8D"!U2d   ��?    ����BvA�C�A��L��G��;�I�{�E>DI]���S� ��3�T0 k� ����U8D"!U2d  
 ��?    ����BwA�C�A��L��G��;�I�s�E>@G]���O� ��3�T0 k� ��� �U8D"!U2d  
 ��?    ����BwA�?�A��L��K��;�I�k�E><F]���G� ��3�T0 k� �(��,�U8D"!U2d  	 ��?    ����BxA�?�A��L��K��;�I�g�E>4D]���?� ��3�T0 k� �4��8�U8D"!U2d  	 ��?    ����B xA�;�A��L��O��;�I�_�E>0C]���;� ��3�T0 k� ,D��H�U8D"!U2d   ��?    ����B�yA�;�A��L��O��;�I�[�E>,A]���3� ��3�T0 k� ,P��T�U8D"!U2d   ��?    ����B�xA�7�A��L��S��;�I�S�K�(@]���+� ��3�T0 k� ,`��d�U8D"!U2d   ��?    ����B�xA�7�A�ߏL��S��;�I�O�K�$>]���#� ��3�T0 k� ,l��p�U8D"!U2d   ��?    ����B�xA�3�A�ߏL��W��;�I�G�K� =]���� ��3�T0 k� ,x��|�U8D"!U2d   ��?    ����B�xA�3�A�ۏL��W��;�I�C�K�<]���� ��3�T0 k� ������U8D"!U2d   ��?    ����B�wA�/�A�ۏL��W��;�I�?�K�:]���� ��3�T0 k� ������U8D"!U2d   ��?    ����B�wA�/�A�׏L��[��;�I�;�K�9]���� ��3�T0 k� ������U8D"!U2d   ��?    ����B�wA�+�A�׏L��[��;�I�7�K�7]����� ��3�T0 k� ������U8D"!U2d   ��    ����B�wA�+�A�ӏL��[��;�I�3�K�6]����� ��3�T0 k� ������U8D"!U2d   ��     ����B�vA�+�A�ӏL��[��;�I�/�K�5]����� ��3�T0 k� L�����U8D"!U2d    ��     ����B�vA�'�A�ϏL��_��;�I�+�K� 4]���� ��3�T0 k� L�����U8D"!U2d    ,�     ����B�vA�'�A�ϏL��_��;�I�'�K��2]���߿��3�T0 k� L�����U8D"!U2d    ��     ����B�vA�#�A�ϏL��_��;�I�#�K��1]���׾��3�T0 k� L�����U8D"!U2d    ��     ����B�vA�#�A�ˏL��_��;�I��K��0]���Ͼ��3�T0 k� L�����U8D"!U2d   ��     ����B�uA��A�ˏL��c��;�I��K��/]��ǽ��3�T0 k� ������U8D"!U2d   ��     ����B�uA��A�ǏL��c��8 I��K��.]������3�T0 k� ������U8D"!U2d   ��     ����B�uA��A�ǏL��c��8 I��K��,]������3�T0 k� ������U8D"!U2d   ��     ����B�uA��A�ǏL��c��8 I��K��+]�������3�T0 k� ������U8D"!U2d   ��     ����B�uA��A�ÏL��g��8 I��K��*]�������3�T0 k� ������U8D"!U2d   ��     ����B�tA��A�ÏL��g��8 I��K��)]�������3�T0 k� ,�����U8D"!U2d   ��     ����B�tA��A�ÏL��g��8 I��K��(]�������3�T0 k� ,�����U8D"!U2d   ��     ����B�tA��A���L��g��8 I��K��']�������3�T0 k� ,�����U8D"!U2d   ��     ����B�tA��A���L��k��8 L�K��&]�������3�T0 k� ,�����U8D"!U2d   ��     ����B�tA��A���L��k��8L�K��%]������3�T0 k� ,�����U8D"!U2d   ��     ����B�sA��A���L��k��8L�K��$]�{����3�T0 k� ������U8D"!U2d   ��     ����B�sA��A���L��k��8L�K��#]�s����3�T0 k� ������U8D"!U2d   ��     ����B�sA��A���L��k��8L�K��"]�k����3�T0 k� ������U8D"!U2d   ��     ����B�sA��A���L��o��8L�K��!]�c����3�T0 k� ������U8D"!U2d   ��     ����B�sA��A���L��o��8L�K�� ]�[����3�T0 k� ������U8D"!U2d   ��     ����B�sA��A���L��o��8L�K��]�S����3�T0 k� <�����U8D"!U2d   ��     ����B�rA��A���L��o��8L��K�]�K���3�T0 k� <�����U8D"!U2d   ��     ����B�rA��A���L��o��8L��K�]{�C��{�3�T0 k� <���U8D"!U2d   ��     ����B�rA��A���L��o��8L��K�]{�;��w�3�T0 k� <���U8D"!U2d   ��     ����B�rA��A���L��o��8L��K�]{�3��s�3�T0 k� <���U8D"!U2d   ��     ����B�rA��A���L��s��8L��K�]{�+��o�3�T0 k� �|��U8D"!U2d   ��     ����B�rA��A���L��s��8L,��K�]{�#��k�3�T0 k� �|��U8D"!U2d   ��    ����B�rA��A���L��s��8L,��K�]{����g�3�T0 k� �x�|U8D"!U2d   ��     ����B�qA��A���L��s��8L,��K�]{����c�3�T0 k� �x�|U8D"!U2d   ��     ����B�qA��A���L��s��8L,�K�]{����_�3�T0 k� �t~�x~U8D"!U2d   ��     ����B�qA���A���L��s��8L,�K�]{����[�3�T0 k� ,t~�x~U8D"!U2d   ��     ����B�qA���A���L��s��8L,�K�]{���� W�3�T0 k� ,p~�t~U8D"!U2d   ��     ����B�qA���A���L��s��8L,�K�]w���� S�3�T0 k� ,p~�t~U8D"!U2d   ��     ����B�qA���A���L��s��8L,�K�]w��� K�3�T0 k� ,l~�p~U8D"!U2d    ��     ����B�qA���A���L��s��8L,�K�]w��� G�3�T0 k� ,l~�p~U8D"!U2d    ��     ����B�pA���A���L��s��8L,�K�]w�߳ C�3�T0 k� �h~�l~U8D"!U2d    ��     ����B�pA���A���L��s��8L,�K�]w�׳?�3�T0 k� �h}�l}U8D"!U2d    .�     ����B�pA���A���L��s��8L,�K�]w�ϳ;�3�T0 k� �d}�h}U8D"!U2d    ��     ����B�pA���A���L��s��8L,�K�]w�ǲ7�3�T0 k� �d}�h}U8D"!U2d    ��    ����B�pA���A���L��s��8L,�K�]w���3�3�T0 k� �d}�h}U8D"!U2d    ��     ����B�pA���A���L��s��8L,�K�]w���/�3�T0 k� L`}�d}U8D"!U2d    ��     ����B�pA���A���L��s��8L,�K�]w���/�3�T0 k� L`}�d}U8D"!U2d    ��     ����B�pA���A���L��o��8L,�K�]w���+�3�T0 k� L\}�`}U8D"!U2d    ��     ����B|pA���A���L��o��8L,�K�]w���'�3�T0 k� L\}�`}U8D"!U2d    ��     ����B|oA���A���L��o��8L,�K�]w���'�3�T0 k� LX}�\}U8D"!U2d    ��     ����B|oA���A���L��o��8L,�K�]s���#�3�T0 k� �X|�\|U8D"!U2d    ��     ����BxoA���A���L��o��8L,�K�]s��� �3�T0 k� �X|�\|U8D"!U2d    ��     ����BxoA���A���L��o��8L,߫K�|]s��� �3�T0 k� �T|�X|U8D"!U2d    ��     ����BtoA���A���L��o��8L,߫K�|
]s��� �3�T0 k� �T|�X|U8D"!U2d    ��     ����BtoA���A���L��o��8L,߫K�x
s�.� �3�T0 k� �T|�X|U8D"!U2d    ��     ����BtoA���A���L��o��8L,߫K�x	s�.w� �3�T0 k� �P|�T|U8D"!U2d    ��     ����BpoA���A���L��o��8L,۫K�ts�.s� �3�T0 k� �P|�T|U8D"!U2d    ��     ����BpoA���A���L��o��8L,۫K�ts�.k� �3�T0 k� �P|�T|U8D"!U2d    ��     ����BpoA���A���L��o��8L,۫CMps�.g� �3�T0 k� �L|�P|U8D"!U2d    ��     ����BlnA���A���L��o��8L,۫CMps�._� �3�T0 k� �L|�P|U8D"!U2d    ��     ����BlnA���A���L��o��8L,׫CMps�.[� �3�T0 k� �L{�P{U8D"!U2d    ��     ����BlnA���A���L��o��8L,׫CMls�.S� �3�T0 k� �H{�L{U8D"!U2d    ��     ����BhnA���A���L��o��8L,׫CMls�.O� �3�T0 k� �H{�L{U8D"!U2d    ��     ����BhnA���A���L��o��8L,׫K�hs�.K� �3�T0 k� �H{�L{U8D"!U2d    ��     ����BhnA���A���L��o��8L,׫K�h-s�.C� �3�T0 k� �D{�H{U8D"!U2d    ��     ����BdnA���A���L��o�#,8L,ӫK�d-s�.?�/��3�T0 k� �D{�H{U8D"!U2d    ��     ����BdnA���A���L��o�#,8L,ӫK�d-o�.;�/��3�T0 k� �D{�H{U8D"!U2d    ��     ����BdnA���A���L��o�#,8L,ӫK�d-o�.3�/��3�T0 k� �@{�D{U8D"!U2d    ��     ����BdnA���A���L��o�#,8L,ӫK�`-o�./�/��3�T0 k� �@{�D{U8D"!U2d    ��     ����B`nA���A���L��o�#,8L,ӫK�` -o�.+�/��3�T0 k� �@{�D{U8D"!U2d    ��     ����B`nA���A���L��o�#,8L,ӫK�` -o�.'�/��3�T0 k� �<{�@{U8D"!U2d    ��    ����B`mA���A���L��o�#,8L,ϫK�_�-o�.#�/��3�T0 k� �<{�@{U8D"!U2d    ��     ����B`mA���A���L��o�#,8LϫK�_�-o�.�/��3�T0 k� �<z�@zU8D"!U2d    ��     ����B\mA���A���L��o�#,8LϫK�[�o�.�/��3�T0 k� �<z�@zU8D"!U2d    ��     ����B\mA���A���L��o�#,8LϫK�[�o�.�/��3�T0 k� �8z�<zU8D"!U2d    ��     ����B\mA���A���L��o�#,8LϫK�[�o�.�/��3�T0 k� �8z�<zU8D"!U2d    ��     ����BXmA���A���L��o��8L˫K�W�o�.�/��3�T0 k� �8z�<zU8D"!U2d    ��     ����BXmA���A���L��o��8L˫K�W�o�.�/��3�T0 k� �8z�<zU8D"!U2d    ��     ����BXmA���A���L��o��8L˫K�W�o�.�/��3�T0 k� �4z�8zU8D"!U2d    ��     ����BXmA���A���L��o��8L˫K�W�o�-��/��3�T0 k� �4z�8zU8D"!U2d    ��     ����BXmA���A���L��o��8L˫K�S�o�-��/��3�T0 k� �4z�8zU8D"!U2d    ��     ����BTmA���A���L��o��8L˫K�S�o�-��/��3�T0 k� �4z�8zU8D"!U2d    ��     ����BTmA���A���L��o��8L˫K�S�]o�-�/��3�T0 k� �0z�4zU8D"!U2d    ��     ����BTmA���A���L��o��8A\˫K�O�]o�-�/��3�T0 k� �0z�4zU8D"!U2d    ��     ����BTmA���A���L��o��8A\˫K�O�]o�-�/��3�T0 k� �0z�4zU8D"!U2d    ��     ����BPmA���A���L��o��8A\˫K�O�]o�-�/��3�T0 k� �0z�4zU8D"!U2d    ��     ����BPmA���A���L��o��8A\˫K�K�]o�-�/��3�T0 k� �0z�4zU8D"!U2d    ��     ����BPlA���A���L��o�#8A\˫K�K�o�-ߪ/��3�T0 k� �,y�0yU8D"!U2d    ��     ����BPlA���A���L��o�#8A�˫K�K�o�-۪/��3�T0 k� �,y�0yU8D"!U2d    ��     ����BPlA���A���L��o�#8A�˫K�K�k�-ת/��3�T0 k� �,y�0yU8D"!U2d    ��     ����BLlA���A���L��o�#8A�˫K�G�k�-Ӫ/��3�T0 k� �,y�0yU8D"!U2d    ��     ����BLlA���A���L��o�#8A�˫K�G�k�-Ϫ/��3�T0 k� �,y�0yU8D"!U2d    ��     ����BLlA���A���L��o�#8A�˫K�G�k�-Ϫ��3�T0 k� �(y�,yU8D"!U2d    ��     ����BLlA���A���L��o�#8L\˫K�G�-k�-˪��3�T0 k� �(y�,yU8D"!U2d    ��     ����BLlA���A���L��o�#8L\˫K�C�-k�-Ǫ��3�T0 k� �(y�,yU8D"!U2d    ��     ����BHlA���A���L��o�#8L\˫K�C�-k�é��3�T0 k� �(y�,yU8D"!U2d    ��     ����BHlA���A���L��o�#8L\˫K�C�-k�����3�T0 k� �$y�(yU8D"!U2d    ��     ����BHlA���A���L��o��8L\˫K�?�-k������3�T0 k� �$y�(yU8D"!U2d    ��     ����BHlA���A���L��o��8L\˫K�?�-k������"s�T0 k� �$y�(yU8D"!U2d    ��     ����BHlA���A���L��o��8L\˫K�?�-k������"s�T0 k� �$y�(yU8D"!U2d    ��     ����BDlA���A���L��o��8L\˫K�?�-k�����"s�T0 k� �$y�(yU8D"!U2d    ��     ����BDlA���A���L��o��8L\˫K�;�k�����"s�T0 k� � y�$yU8D"!U2d    ��     ����BDlA���A���L��o��8L\˫K�;�k�����"s�T0 k� � y�$yU8D"!U2d    ��     ����BDlA���A���L��o��8Ll˫K�;�k����"s�T0 k� � y�$yU8D"!U2d    ��     ����BDlA���A���L��o��8Ll˫K�;�k����"s�T0 k� � y�$yU8D"!U2d    ��     ����BDlA���A���L��o��8Ll˫K�;�k����"s�T0 k� � y�$yU8D"!U2d    ��     ����B@lA���A���L��o��8Ll˫K�7�g�ퟪ��"s�T0 k� � y�$yU8D"!U2d    ��     ����B@kA���A���L��o��8Ll˫K�7�g�ퟪ��"s�T0 k� � y�$yU8D"!U2d    ��     ����B@kA���A���L��o��8Ll˫K�7�c�훪��"s�T0 k� �x� xU8D"!U2d    ��     ����B@kA���A���L��o��8Ll˫K�7�c������3�T0 k� �x� xU8D"!U2d    ��     ����B@kA���A���L��o��8Ll˫K�7�]_������3�T0 k� �x� xU8D"!U2d    ��     ����B@kA���A���L��o��8Ll˫K�3�]_������3�T0 k� �x� xU8D"!U2d    ��     ����B<kA���A���L��o��8Ll˫K�3�]_������3�T0 k� �x� xU8D"!U2d    ��     ����B<kA���A���L��o��8Ll˫K�3�][������3�T0 k� �x� xU8D"!U2d    ��     ����B<kA���A���L��o��8Ll˫K�3�][������3�T0 k� �x� xU8D"!U2d    ��     ����B<kA���A���L��o��8Ll˫K�3�]W������3�T0 k� �x�xU8D"!U2d    ��     ����B<kA���A���L��o��8Ll˫K�3�]W������3�T0 k� �x�xU8D"!U2d    ��     ����B<kA���A���L��o��8Ll˫K�/�]W������3�T0 k� �x�xU8D"!U2d    ��     ����B<kA���A���L��o��8Ll˫K�/�]S�����3�T0 k� �x�xU8D"!U2d    ��     ����B<kA���A���L��o��8Ll˫K�/�]S����{�3�T0 k� �x�xU8D"!U2d    ��     ����B8kA���A���L��o��8Ll˫K�/�]S��w�"��T0 k� �x�xU8D"!U2d    ��     ����B8kA���A���L��o��8Ll˫CM/�]O��o�"��T0 k� �x�xU8D"!U2d    ��     ����B8kA���A���L��o��8Ll˫CM/�]O�{�k�"��T0 k� �x�xU8D"!U2d    ��     ����B8kA���A���L��o��8Ll˫CM+�]K�-{�c�"��T0 k� �x�xU8D"!U2d    ��     ����B8kA���A���L��o��8Ll˫CM+�]K�-w�_�"��T0 k� �x�xU8D"!U2d    ��     ����B8kA���A���L��o��8Ll˫CM+�]K�-w�W�"��T0 k� �x�xU8D"!U2d    ��     ����B8kA���A���L��o��8Ll˫CM+�]G�-s�S�"��T0 k� �x�xU8D"!U2d    ��     ����B8kA���A���L��o��8Ll˫CM+�]G�-s�K�"��T0 k� �x�xU8D"!U2d    ��     ����B8kA���A���L��o��8Ll˫CM+�]G�-o�C�"��T0 k� �x�xU8D"!U2d    ��     ����B4kA���A���L��o��8Ll˫CM+�]C�-o�?�"��T0 k� �x�xU8D"!U2d    ��     ����B4kA���A���L��o��8Ll˫CM'�]C�-k�7�"��T0 k� �x�xU8D"!U2d    ��     ����B4kA���A���L��o��8Ll˫CM'�]C�-k��/�3�T0 k� �x�xU8D"!U2d    ��     ����B4kA���A���L��o��8Ll˫CM'�]C�-g��+�3�T0 k� �x�xU8D"!U2d    ��     ����B4kA���A���L��o��8Ll˫C]'�]?�-g��#�3�T0 k� �x�xU8D"!U2d    ��     ����B4kA���A���L��o��8Ll˫C]'�]?�-c���3�T0 k� �x�xU8D"!U2d    ��     ����B4kA���A���L��o��8Ll˫C]'�]?�-c���3�T0 k� �x�xU8D"!U2d    ��     ����B4kA���A���L��o��8Ll˫C]'�];�-c���3�T0 k� �x�xU8D"!U2d    ��     ����B4kA���A���L��o��8Ll˫C]'�];�-_���3�T0 k� �x�xU8D"!U2d    ��     ����B4kA���A���L��o��8Ll˫C]#�];�-_����3�T0 k� �x�xU8D"!U2d    ��     ����B0kA���A���L��o��8Ll˫C]#�];�-[����3�T0 k� �x�xU8D"!U2d    ��     ����B0kA���A���L��o��8Ll˫C]#�]7�-[����3�T0 k� �x�xU8D"!U2d    ��     ����B0kA���A���L��o��8Ll˫C]#�]7�-W�>��3�T0 k� �x�xU8D"!U2d    ��     ����B0kA���A���L��o��8Ll˫C]#�]7�-W�>��3�T0 k� �x�xU8D"!U2d    ��     ����B0kA���A���L��o��8Ll˫C]#�]7�-W�>��3�T0 k� �x�xU8D"!U2d    ��     ����B0jA���A���L��o��8L\˫Cm#�]3�-S�>��3�T0 k� �w�wU8D"!U2d    ��     ����B0jA���A���L��o��8L\˫Cm#�]3�-S�>��3�T0 k� �w�wU8D"!U2d    ��     ����B0jA���A���L��o��8L\˫Cm�]3�-S�>��3�T0 k� �w�wU8D"!U2d    ��    ����B0jA���A���L��o��8L\˫Cm�]3�-O�>��3�T0 k� �w�wU8D"!U2d    ��     ����B0jA���A���L��o��8L\˫Cm�]/�-O�>��3�T0 k� �w�wU8D"!U2d    ��     ����B0jA���A���L��o��8L\˫Cm�]/�-K�>��3�T0 k� �w�wU8D"!U2d    ��     ����B0jA���A���L��o��8BL˫Cm�]/�-K�>��3�T0 k� �w�wU8D"!U2d    ��     ����B0jA���A���L��o��8BL˫Cm�]/�-K�>��3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8BL˫Cm�]+�-G�>��3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8BL˫Cm�]+�-G�N��3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8BL˫Cm�]+�-G�N��3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8BL˫C}�]+�-C�N�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8@˫C}�]+�-C�Nw�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8@˫C}�]'�-C�No�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8@˫C}�]'�-?�Ng�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8@˫C}�]'�-?�N_�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8@ϫI]�]'�-?�NW�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8K�ϫI]�]'�-?�NO�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8K�ϫI]�]#�-;�NG�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8K�ϫI]�]#�-;�N?�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8K�ϫI]�]#�;�^;�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8K�ϫIm�]#�;�^3�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8K�ϫIm�]#�;�^+�3�T0 k� �w�wU8D"!U2d    ��     ����B,jA���A���L��o��8K�ӫIm�]#�;�^#�3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�ӫIm�]�;�^�3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�ӫIm�]�;�>�3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�ӫCM�]��;�>�3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�ӫCM�]��7�>�3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�ӫCM�]��7�=��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�ӫCM�]��7�=��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�׫CM�]��7�=��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�׫CM�]��7�=��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�׫CM�]��7�=��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�׫CM�]��7�=��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�׫CM�]��3�=��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�׫CM�]��3�=��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�׫C]�]��3�=��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�׫C]�]��3�M��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�׫C]�]��3�M��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�۫C]�]��3�M��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�۫C]�]��3�M��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8K�۫C]�]��3�M��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8	K�۫C]�]��3�M��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8	K�۫C]�]��3�M��3�T0 k� �w�wU8D"!U2d    ��     ����B(jA���A���L��o��8	K�۫C]�]��3�M��3�T0 k� �w�wU8D"!U2d    ��     ����B�C�D�P'�dp|C�E�C�E�W��v��2B�
T0 k� ��f��fU8D"!U2d    ��    � 8 �C�D�P( ft|C�E�G�Eo�X��v��2B�
T0 k� ��d��dU8D"!U2d    ��    � 9 �C�D�P*h||C�E�K�Eo�Y��v��2C�
T0 k� ��c��cU8D"!U2d    ��    � : 	PC�D�P+j�|C�E�O�Eo�[��u��B C�
T0 k� ��b��bU8D"!U2d    ��    � ; PC��D�P,�k�|C�E�O�Eo�\��u��B C�
T0 k� �b��bU8D"!U2d    ��    � < P C��D�P-�m��|C�E�S�E` ]��u��B$D�
T0 k� �c��cU8D"!U2d    ��    � < _�C��EP0�p��|C�E�[�E``��t��B(D�
T0 k� �c��cU8D"!U2d    ��    � < _�C��EP1� r��|C�E�[�E`b��s��R,D�
T0 k� �c��cU8D"!U2d    ��    � <  _�C��EP2�$s��|C�E�_�E`c��s��R0D3�
T0 k� �c��cU8D"!U2d    ��    � <��_�C��EP4�(t��|C�E�c�E`d��r��R0D3�
T0 k� �c��cU8D"!U2d    ��    � <��_�C��EP5�0v��|C�E�c�E`f��r��R4E3�
T0 k� �b��bU8D"!U2d    ��    � <��O�AP�EoP6�4w��|C�E�g�EPg��q��R8E3�
T0 k� �a��aU8D"!U2d    ��    � <��O�AP�EoP8�8x��|C�E�g�EPi��q��R<E3�
T0 k� �_��_U8D"!U2d    ��    � <��O�AP�EoP9�<y��|C�E�k�EPj�p��
�@E3�
T0 k� �]��]U8D"!U2d    ��    � <��O�AP�EoP;�Dz��|C�E�k�EP l�o��
�DE3�
T0 k� �[��[U8D"!U2d    ��    � <��O�E��"EoL>�P|�� |C�E�o�EP$n�n��
�LF3�
T0 k� ��Y��YU8D"!U2d    ��    � <��O�E��#EoL?�T}�� |C�E�o�EP$p�m��
�PF3�
T0 k� ��W��WU8D"!U2d    ��    � <��O�E��$EoLA}X~}�!|C�E�o�C�(q�l��
�XF3�
T0 k� ��V��VU8D"!U2d    ��    � <��O�E�%EoHB}`}�!|C�E�s�C�(r�k��
�\F3�
T0 k� �|U��UU8D"!U2d    ��    � <��ϸE�'EoHD}d�~ !|C�E�s�C�(t��j��
�`F3�
T0 k� �xT�|TU8D"!U2d    ��    � <��ϰE�(EoHE}h~!|C�E�s�C�(u��i��
�dF3�
T0 k� �pS�tSU8D"!U2d    ��    � <��ϬE�)EoDG}p~!|C�E�s�C�,v��h��
�lF3�
T0 k� �lR�pRU8D"!U2d    ��    � <��ϠE�,E_@J}x~~!|C�E�s�C�,y��f��
�tG3�
T0 k� �lP�pPU8D"!U2d    ��    � <��ϜE��-E_@L}�~~ !|C�E�s�C�,z��e��
�|G3�
T0 k� �tN�xNU8D"!U2d    ��    � <��ϔE�/E_<M}�}~(!|C�E�o�EP({�|d��
�G3�
T0 k� �xM�|MU8D"!U2d    ��    � <��ϐE�0E_8N}�}~,!|C�E�o�EP(|�tc��
�G3�
T0 k� �xL�|LU8D"!U2d    ��    � <��ψE�2E_8P}�|~4 |C�E�o�EP(}�pb��
�G3�
T0 k� �tK�xKU8D"!U2d    ��    � <��τE��4E_4Q}�{n8 |C�E�o�EP(~�la��
�G3�
T0 k� �tI�xIU8D"!U2d    ��    � <��πE��5E_0Sm�{n@ |C�E�k�EP(��h_��
�G3�
T0 k� �tH�xHU8D"!U2d    ��    � <���|E��7E_0Tm�znD|C�E�k�EP$�d^��
�H3�
T0 k� �pG�tGU8D"!U2d    ��    � <���p
Dpx=E_(Wm�ynP|C�E�g�EP �X[��
�H3�
T0 k� �hD�lDU8D"!U2d    ��    � <���l
DptAE_$Xm�xnT|C�E�c�E@ ~�TZ��
�H3�
T0 k� �`B�dBU8D"!U2d    ��    � <���h
DplDE_ Y=�wnX|C�E�c�E@~ PX��
�H3�
T0 k� �dC�hCU8D"!U2d    ��    � <���h	DphGEO[=�vn\|C�E�_�E@~ LW��
��H3�
T0 k� �hC�lCU8D"!U2d    $�    � <���d	DphGEO\=�und|C�E�_�E@} HW��
��H3�
T0 k� �lE�pEU8D"!U2d    �    � <���`OphHEO]=�tnh|C�E�[�E@} @W��
��H3�
T0 k� �lF�pFU8D"!U2d    �� 	   � <���\OphHEO^=�tnl|C�E�W�E�| 8V��
��I3�
T0 k� �dF�hFU8D"!U2d    �� 	   � <���XOpdIEO_=�s^l|C�E�W�E�| 4V��
��I3�
T0 k� �`F�dFU8D"!U2d    �� 	   � <���POpdJEOa=�q^t|C�E�O�E�{ (V����I3�
T0 k� �TF�XFU8D"!U2d    �� 	   � <���LOp`JEN�bm�p^x|C�E�K�E�{ $V����I3�
T0 k� �PF�TFU8D"!U2d    �� 	   � <��?HOp`KEN�cm�o^x|C�E�G�E�z  V��� I3�
T0 k� �LE�PEU8D"!U2d    �� 	   � <��?HOp`LEN�dm�n�||C�E�G�E� z U���I3�
T0 k� �HE�LEU8D"!U2d    �� 	   � <��?DOp\LEN�dm�l�||C�E�C�E� z UR���I3�
T0 k� �DE�HEU8D"!U2d    �� 	   � <��?@Op\ME>�em�k�|C�E�?�E��y�TR���I3�
T0 k� �8H�<HU8D"!U2d    �� 	   � <��?<Op\ME>�fm�j�|C�E�;�E��y�TR���I3�
T0 k� �0K�4KU8D"!U2d    �� 	   � <��/<OpXNE>�fm�i�|C�E�;�E��y�TR���J3�
T0 k� �(M�,MU8D"!U2d    �� 	   � <��/8OpXNE>�g]�h�|C�D�7�Eo�y�SR��� J3�
T0 k� �$N�(NU8D"!U2d    �� 	   � <��/8OpXOE>�g]�g�|C�D�3�Eo�x�S����$J3�
T0 k� � O�$OU8D"!U2d    �� 
   � <��/4OpTPE>�h]�e�|C�D�/�Eo�x� R����,J3�
T0 k� �O�OU8D"!U2d    �� 
   � <���0OpTPCN�h]�d�|C�D�+�Eo�x��R����0J3�
T0 k� �P�PU8D"!U2d    �� 
   � <���0OpTQCN�i��b�|C�D�'�E_�w��R����0J3�
T0 k� �T�TU8D"!U2d    �� 
   � <���,OpPQCN�i��a�|C�D�'�E_�w��R����4J3�
T0 k� �V�VU8D"!U2d    �� 
   � <���,OpPRCN�i��`��|C�D�#�E_�w��Q����8J3�
T0 k� �X�XU8D"!U2d    �� 
   � <���(OpPRCN�i��_��|C�D��E_�w��Q����8J3�
T0 k� �Z�ZU8D"!U2d    �� 
   � <���(OpPSCN�i��^��|C�D��E_�v��Q����<J3�
T0 k� �[�[U8D"!U2d    �� 
   � <���$OpLSCN�i��]��|C�D��C��v��Q����<K3�
T0 k� �\�\U8D"!U2d    �� 
   � <���$OpLTCN�i��\��|C�D��C�v��Q����@K3�
T0 k� �]�]U8D"!U2d    �� 
   � <��� OpLTCN�i��[~�|C�D��C�v �Q����@K3�
T0 k� �Y�YU8D"!U2d    �� 
   � <��� OpLTCN�i�[~�|C�D��C�u �Q����DK3�
T0 k� � V�$VU8D"!U2d    �� 
   � <���E`HUCN�h�Z~�|C�D��C�u �Q����DK3�
T0 k� �(S�,SU8D"!U2d    �� 
   � <���E`HUE>�h�Y~�|C�D��E�u �Q��DK3�
T0 k� �,Q�0QU8D"!U2d    �� 
   � <���E`HVE>�h�X~||C�D��E�u �Q��DK3�
T0 k� �0P�4PU8D"!U2d    �� 
   � <���E`DWE>�g�Wn||C�D��E�u �Q��DK3�
T0 k� �4O�8OU8D"!U2d    �� 
   � <���E`DWE>�g�Wn||C�D��E�u �Q��DK3�
T0 k� �8N�<NU8D"!U2d    �� 
   � <���E`@XE>�g}�Vnx|C�E��E�tO�Q��DK3�
T0 k� �,K�0KU8D"!U2d    �� 
   � <��?	EP<YE>�e}�Unx|C�E��E�tO�Q��DK3�
T0 k� �$I�(IU8D"!U2d    �� 
   � <��?	EP<ZE>�e}�U�t|C�E���D?|tO�Q��DL3�
T0 k� � G�$GU8D"!U2d    �� 
   � <��?
EP8ZE.�d}�T�t|C�E���D?xsO�Q��@L3�
T0 k� �F� FU8D"!U2d    �� 
   � <��?EP4[E.�d��T�p|C�E���D?psO�Q��@L3�
T0 k� �E�EU8D"!U2d    �� 
   � <��?EP0\E.�c��S�p|C�E���D?lsO�Q��@L3�
T0 k� �D�DU8D"!U2d    �� 
   � <���EP0\E.|b��S�l|C�F��D?ds��Q��<L3�
T0 k� �D�DU8D"!U2d    ��    � <���EP,]E.xa��Sl|C�F��I�`s��Q��<L3�
T0 k� � D�DU8D"!U2d    ��    � <��� E@(]B�xa��Sh!�C�F�I�\s��Q{�8L3�
T0 k� ��D��DU8D"!U2d    ��    � <��� E@$^B�t`�Sd!�C�F�I�Xs��Qw�8L3�
T0 k� ��D��DU8D"!U2d    ��    � <��� E@ ^B�t_�R`!�C�F�I�Ps��Qo�4L3�
T0 k� ��D��DU8D"!U2d    ��    � <��� E@_B�t^�R`!�C�D��I�Ls��Qk�0L3�
T0 k� ��E��EU8D"!U2d    ��    � <��� E@_B�p]�R
\!�C�D��I�Hs��Qc�0L3�
T0 k� ��F��FU8D"!U2d    ��    � <����P�`B�p\�R
X!�C�D��I�Ds��Q_�,L3�
T0 k� ��F��FU8D"!U2d    ��    � <����P�`B�p\�R
T!�C�D��I�@s��QW�(L3�	T0 k� ��F��FU8D"!U2d    ��    � <����P�aB�l[
�R
P!�C�D��I�@s��QO�$L3�	T0 k� ��F��FU8D"!U2d    ��    � <����P�aB�lZ
�Q
L!�@ D��I�<s��QK� L3�	T0 k� ��D��DU8D"!U2d    ��    � <��� P�bClY
|Q
H!�@ D��I�8s��PC��L3�T0 k� ��C��CU8D"!U2d    ��    � <�� P� bClX
xQ
D!�@ D��I�4s��P;��M3�T0 k� ��C��CU8D"!U2d    ��    � <�� P��cClV
pQ
<|<D��I�0s��O+��M3�T0 k� ��B��BU8D"!U2d    ��    � <�� P��cClU
lQ
8|<D��I�,s��O#��M3�T0 k� ��B��BU8D"!U2d    ��    � <�� P��dClS
dQ
0|<D��I�,s��O���M3�T0 k� ��A��AU8D"!U2d    ��    � <��/P��dClR
`P
.,|<D��I�(s��N���M3�T0 k� ��A��AU8D"!U2d    ��    � <��/!P��eClQ
\P
.(|<D��I�(s��N��� M3�T0 k� ��@��@U8D"!U2d    ��    � <��/"P��eClP
TP
. |<D��I�(s��M����M3�T0 k� ��?��?U8D"!U2d    ��    � <��/#P��eClO
PP
.|<I��I�$s��L�����M3�T0 k� ��>��>U8D"!U2d    ��    � <��/%P��fClN
-LP
.|<I��I�$s��L�����M3�T0 k� ��>��>U8D"!U2d    ��    � <���&P��fCpL
-DP
.|<I��I�$s��K�����M3�T0 k� ��=��=U8D"!U2d    ��    � <���'P��gCpK
-@P
.|<I��I� s��K�����M3�T0 k� ��<��<U8D"!U2d    ��    � <���)P��gCpJ
-8O
.!�<I��I� s��J�����M3�T0 k� ��;��;U8D"!U2d    ��    � <���*P��gCtI
-4O
. !�<J�I� s��I�����M3�T0 k� ��;��;U8D"!U2d    ��    � <���,EO�hCtG,O
-�!�<J�I� s��H�����M3�T0 k� ��:��:U8D"!U2d    ��    � <���-EO�hCtF$O
-�!�<J�I� s��G�����M3�T0 k� ��7��7U8D"!U2d    ��    � <���/EO�hCxE O
�!�<J�I� s��G����M3�T0 k� ��4��4U8D"!U2d    ��    � <���2EO�iC|BO
�!�<F�I� s��E���M3�T0 k� ��1��1U8D"!U2d    ��    � <��� 3EO�iC|AO
�!�<F�A� s��D���N3�T0 k� ��/��/U8D"!U2d    ��    � <��� 5EO�iC�?O
�!�<F�A� s��C���N3�T0 k� ��-��-U8D"!U2d    ��    � <��?$6EO�iC.�>�N��!�<F�A� s��B	����N3�T0 k� ��,��,U8D"!U2d    ��    � <��?$8E?�iC.�<�N��!�<F�A� s��@	����N3�T0 k� ��*��*U8D"!U2d    ��    � <��?(:E?�iC.�;�N��|<E���A� s��?	����N3�T0 k� ��)��)U8D"!U2d    ��    � <��?(;E?�hC.�9,�N��|<E���A_ s��>	����N3�T0 k� ��'��'U8D"!U2d    ��    � <��?,=E?�hC.�8,�N��|<E���A_ s��=	���N3�T0 k� ��&��&U8D"!U2d    ��    � <��/,?E?�hC.�6,�N��|<E���A_ s��;	�w��N3�T0 k� ��%��%U8D"!U2d    ��    � <��/0@E?�gC.�5,�N��|<E���A_ s��:	�s��xN3�T0 k� ��#��#U8D"!U2d    ��    � <��/4BE?�gC.�3,�N��|<E���A_ s��9	�o��pN3�T0 k� ��"��"U8D"!U2d    ��    � <��/4DE?�gC.�2 l�N��|<E���A_ s��7	�g��hN3�T0 k� ��!��!U8D"!U2d    ��    � <��/8FE/�fC.�0 l�N��|<E��A_ s��6	�c��`N3�T0 k� ����U8D"!U2d    ��    � <��/@IE/�eE��- l�N
�|<E��A_ s��3	�[��PN3�T0 k� ����U8D"!U2d    ��    � <��/DKE/�dE��, l�N
�|<E��A_ s�1	�W��HN3�T0 k� ����U8D"!U2d    ��(    � <��/DME/�dE��* l�N
�|<E��A s�/	�S��@N3�T0 k� ����U8D"!U2d    ��(    � <��HNE/�cE��( l�N
�|<E��A s�.	�O��8N3�T0 k� ����U8D"!U2d    ��(    � <��LPE��bE��' l�N
�|<E��A s�,	�K��0N3�T0 k� ����U8D"!U2d    ��(    � <��PRE�|bE��% l�N
�|<E��A s�*	�G��(N3�T0 k� ����U8D"!U2d    ��(    � <��TTE�|aE��#�N
�|<E��A s�(	�C�� N3�T0 k� ����U8D"!U2d    ��(    � <��TTE�|aE��!�N
�|<E��A s�'	�?��N3�T0 k� ����U8D"!U2d    ��(    � <��TTE�|aE�� �N
�|<E��A s�%	�;��N3�T0 k� ����U8D"!U2d    ��(    � <�� TTE�|aE���N
x|<CO#�A s�!	�7���M3�T0 k� ����U8D"!U2d    ��(    � <�� TTE�|aE���N
t|<CO'�A s�	�3���M3�T0 k� ����U8D"!U2d    ��(    � <�� TTE��aE��|N
-p|<CO'�A so�	�3���M3�T0 k� ����U8D"!U2d    ��(    � <�� TTCO�aE��|N
-h|<CO+�A so�	�/���M3�T0 k� �t�xU8D"!U2d    ��(    � <�� TTCO�aE���xN
-d|<CO+�@� so�	�/���L3�T0 k� �h�lU8D"!U2d    ��(    � <��OXTCO�aE���xM
-\|<CO/�@� so|	�+���L3�T0 k� �\�`U8D"!U2d    ��(    � <��OXTCO�aE���tM
-X|<CO/�@� so|	�+���L3�T0 k� �X�\U8D"!U2d    ��(    � <��OXTCO�aE���tM
-T|<CO/�@� sox	�'���K3�T0 k� �P �T U8D"!U2d    ��(    � ;��O\SCO�aE���pM
-L|<C_3�@� sot	�'��K3�T0 k� �K��O�U8D"!U2d    ��(    � :��O\SCO�`E���pM
-H|<C_3�@� sop	�'��J3�T0 k� �G��K�U8D"!U2d    ��(    � 9��\SCO�`E��	�lM
-@|<C_3�@� sop	�'��I3�T0 k� �C��G�U8D"!U2d    ��(    � 8��\RCO�_E���lL
-8|<C_3�@� sol	�#��I3�T0 k� �C��G�U8D"!U2d    ��(    � 7��`RCO�_E���lL
-4|<C_3�@� soh		�#��H3�T0 k� �?��C�U8D"!U2d    ��(    � 6��`QCO�^E���lL,|<C_3�@� s_d	�#��H3�T0 k� �?��C�U8D"!U2d    ��(    � 5��`QCO�^E���lK$|<C_3�@� s_`	�#��G3�T0 k� �?��C�U8D"!U2d    ��(    � 4��`PC_�]P^� �lK |<C_3�@� s_\	�#��G3�T0 k� �8 �< U8D"!U2d    ��(    � 3��`PC_�\P^���hJ|<C_3�@� s_X	�#��F3�T0 k� �4�8U8D"!U2d    ��(    � 2��`PC_�\P^���hJ|<@�3�@� s_W�	�#��|F3�T0 k� �0�4U8D"!U2d    ��(    � 1��`OC_�\P^���hI|<@�3�@� s_S�	�#��tE3�T0 k� �,�0U8D"!U2d    ��(    � 0��`OC_�[P^���hI|<@�3�@� s�O�	�#��pE3�T0 k� �+��/�U8D"!U2d    ��(    � /��`OC_�ZP_��lH�|<@�3�@� s�K�	���hD3�T0 k� �'��+�U8D"!U2d    ��(    � .��`NC_�YPo��lH�|<@�3�@� s�G�	���`D3�T0 k� �#��'�U8D"!U2d    ��(    � -��`NC_�XPo��lG,�|<@�3�@� s�G�	���\D3�T0 k� �#��'�U8D"!U2d    �(    � ,��`NC_�XPo��lF,�|<CO3�@� s�G�	���TC3�T0 k� �#��'�U8D"!U2d    ��(    � +��`NC_�XPo��lF,�|<CO3�@� s�G�	���PC3�T0 k� �#��'�U8D"!U2d    ��(    � *��`MC_�VPo��pD,�|<CO3�@� s�G�Q��DB3�T0 k� �#��'�U8D"!U2d    ��(    � (���`MCo�UPo��pC�|< CO3�@� s�G�Q��<A3�T0 k� �#��'�U8D"!U2d    ��(    � &���`MCo�TPo�|pB�|< CO3�@� s�G�Q��8@3�T0 k� �#��'�U8D"!U2d    ��(    � %���`LCo�SPo�|pB�|< CO3�@� s�G�Q��4?3�T0 k� ���#�U8D"!U2d    ��(    � $���\LCo�RP_�|pA�|< CO3�@� s�G�Q�,?3�T0 k� ����U8D"!U2d    ��(    � "���\KCo�QP_�|t@�|< CO3�@� s�G���(>3�T0 k� ����U8D"!U2d    ��(    �  ��o\KCo�PP_�|t?�|< CO3�@� s�G���$=3�T0 k� ����U8D"!U2d    ��(    � ��o\JCo�NP_��t=�|< CO3�@� s�C��� <3�T0 k� ����U8D"!U2d    ��(    � ��oXICo�KP^���t;�|?�CO3�@� s�C����:3�T0 k� ����U8D"!U2d    ��(    � ��oXHCo�JCN���x:�|?�C_3�@� s�?����:3�T0 k� ����U8D"!U2d    ��(    � ��oXHCo�ICN���x9��|?�C_3�@� s�?����93�T0 k� ����U8D"!U2d    ��(    � ��_TGC�GCN���x8��|?�C_3�@� s�;����83�T0 k� ����U8D"!U2d    ��(    � ��_TFC�ECN���x6��|?�C_3�@� s�;����73�T0 k� ����U8D"!U2d    ��(    � ��_PFC�DCN���x5��|?�C_3�@� s�;����63�T0 k� ����U8D"!U2d    ��(    � ��_LDC�AN>���|2��|?�C_3�@� s�7�A���3"��T0 k� ����U8D"!U2d    ��(    � ��_LDC�?N>���|1��|?�C_3�@� s�3�A���2"��T0 k� ����U8D"!U2d    ��(    � ��_HCC�=N>���|/��|?�C_3�@� s�3�A���1"��T0 k� ����U8D"!U2d    ��(    � 
��_DBC�;N>���|.|�|?�C_3�@� s�/�A���0"��T0 k� ����U8D"!U2d    ��(    � ��O@BC�9N>���|,|||?�C_3�@� s�/�A���/"��T0 k� �����U8D"!U2d    ��(    � ��O<AC�7N>���+|x|;�Co3�@� so+�����."��T0 k� �����U8D"!U2d    ��(    � ��O8@C�4N>���'|t|;�Co3�@� so#�����+"��T0 k� ������U8D"!U2d    ��(    � ��O4@CO�2N>���&t|;�Co3�@� so#�����*"��T0 k� �����U8D"!U2d    ��    �  ��O0@CO�0N>���$p|;�Co3�@� so�����)"��T0 k� ����U8D"!U2d    ��    �����O,?CO�.N>���"p|;�Co3�@� s_�����'3�T0 k� �����U8D"!U2d    ��    �����O(?CO�,N>��� l|;�Co3�@� s_�����&3�T0 k� �����U8D"!U2d    ��    �����?$?CO�)N>���l|;�Co3�@� s_�����%3�T0 k� ����U8D"!U2d    ��    �����? ?E/�'N>���l|;�Co3�@� s_�����$3�T0 k� ����U8D"!U2d    ��    �����??E/�#N>���h
|;�Co3�@� so�����!3�T0 k� �Ӹ�׸U8D"!U2d    ��    �����??E/�!N>���h|;�C3�@� so����� 3�T0 k� �Ƕ�˶U8D"!U2d    ��    �����O?E/�N>�	܄h|;�C3�@� sn���#���3�T0 k� ������U8D"!U2d    ��    �����O?E/�N>�	܄�d|;�C3�@� sn���#���3�T0 k� ������U8D"!U2d    ��    �����O?E/�N>�	܄�d|;�C3�@� sn��#���3�T0 k� ������U8D"!U2d    ��    �����O?E�N>�	܄�d|7�C3�@� s���#���3�T0 k� ������U8D"!U2d    ��    ����O@E�N>�	܄�h|7�I_3�@� s���#���"s�T0 k� ������U8D"!U2d    ��    ����~��@E�E��	��h|7�I_3�@� s���#���"s�T0 k� ������U8D"!U2d    ��    ����}��AE�E�ߐ	��h|;�I_3�@� s�ߧ�#���"s�T0 k� ������U8D"!U2d    ��    ����|��AE�E�ߎ	��l|;�I_3�@� s�ۦ�#���"s�T0 k� ������U8D"!U2d    ��    ����{��AE�E�ߏ	��l|;�A3�@� s�פ�'���"s�T0 k� ������U8D"!U2d    ��    ����z��BE�
E�ߏ	��l �;�A3�@� s�ӣ�'� �"s�T0 k� ������U8D"!U2d    ��    ����y��BE�E�ې	܄�s��;�A3�@� s�ϡ�'� �"s�T0 k� ������U8D"!U2d    ��    ����x��CE�E�ې	܄�s��;�A/�@� s�ˠ�'� �"s�T0 k� ������U8D"!U2d    ��    ����w��CE�E�ې	܄�w��;�A/�@� s�ß�'� �"s�T0 k� ������U8D"!U2d    �    ����u��DEE�׏	܄�{��;�E�+�@� s����'� �"s�T0 k� ������U8D"!U2d    ��    ����s��EE��E�׎	����;�E�+�@� s����'� �3�T0 k� �{���U8D"!U2d    ��    ����q��EE��E�׎	����;�E�'�@� s����'�p�3�T0 k� �w��{�U8D"!U2d    ��    ����p��FE��E�Ӎ	�|���;�E�'�@� s����'�p�3�T0 k� �s��w�U8D"!U2d    ��    ����o�FE��E�Ӎ	�|���;�E�#�@� s����'�p�3�T0 k� �o��s�U8D"!U2d    ��    ����n�FE�#�E�ύ	�|���;�E��@� s����+�p�
3�T0 k� �k��o�U8D"!U2d    ��    ����m�GE�'�E�ό	܄|���;�E��@� s����+�p�	3�T0 k� �g��k�U8D"!U2d    ��    ����l�GE�/�E�ˌ	܄|���;�E��A s���q+�p�3�T0 k� �c��g�U8D"!U2d    ��    ����k�HE�3�E�ˌ	܄|���;�E��A s���q+�p�3�T0 k� �_��c�U8D"!U2d    �    ����i�HE�;�E�ǌ	܄|���;�E��A s���q+�p�3�T0 k� �W��[�U8D"!U2d    ��    ����g��HE�?�E�Ì	܄����;�Eo�A s���q+�`�3�T0 k� �S��W�U8D"!U2d    ��    ����e��IE�G�E	�����;�Eo�A s���q+�`�3�T0 k� �K��O�U8D"!U2d    ��    ����c��JEpS�On��	�����;�Eo�A_ s�{�a'�`� 3�T0 k� �C��G�U8D"!U2d    ��    ����a�|JEpW�On��	�����;�Eo�A_ s�s�a'�`��3�T0 k� �;��?�U8D"!U2d    ��    ����_NxKEp_�On��	����;�Eo�A_ s�o�a'�`��3�T0 k� �7��;�U8D"!U2d    ��    ����]NpKEpc�On�������;�E^��A_s�k�a'�`��3�T0 k� �/��3�U8D"!U2d    ��    ����[NhLEpk�On�������;�E^��A_s�c�a#�`��3�T0 k� �+��/�U8D"!U2d    ��    ����YN`LEpo�On�������;�E^��C�s�_�Q#�`��3�T0 k� �'��+�U8D"!U2d    ��    ����WN\MEps�On�������;�E^�C�s�[�Q�`��3�T0 k� �#��'�U8D"!U2d    ��    ����VNTNEp{�On�������;�E^�C�s�S�Q�`��3�T0 k� ���#�U8D"!U2d    ��    ����TNLNEp�On��L����;�C��C�s�O�Q�`��3�T0 k� ����U8D"!U2d    �    ����RNDOEp��On��L����;�C��C�s�K�Q�P��3�T0 k� ������U8D"!U2d   ��    ����P�<PEp��On��L����;�C�ߖEOs�G�Q�P��3�T0 k� ����U8D"!U2d   ��    ����N�4QEp��On��L�����;�C�ۖEOs�?�Q�P��3�T0 k� �ӱ�ױU8D"!U2d   ��    ����L�0QEp��On�L�����;�C�חEOr�;���P��3�T0 k� ����öU8D"!U2d   ��    ����J�(REp��On�܈����;�C�ϗEOr�7���P��3�T0 k� ������U8D"!U2d   ��    ����H� SA���On{�܈����;�C�˘EOr�3������3�T0 k� ������U8D"!U2d   ��    ����G�TA���Onw�܈����;�C�ǘEOr�/������3�T0 k� ������U8D"!U2d   ��?    ����F�UA���Ons�܈����;�CE?r�+������3�T0 k� �o��s�U8D"!U2d   ��?    ����E�VA���Ono�܈����;�CE? q�'�������3�T0 k� �[��_�U8D"!U2d   ��?    ����D� WA���Onk�L�����;�C���E? q�#�������3�T0 k� �G��K�U8D"!U2d   ��?    ����C��XE`��Ong�L�����;�C���E>�q��������3�T0 k� �7��;�U8D"!U2d  	 ��? 
   ����B��YE`��Onc�L�|���;�C���E>�p��������3�T0 k� �#��'�U8D"!U2d  	 �? 
   ����B�ZE`��On_�L�|���;�C���E��p��������3�T0 k� ����U8D"!U2d  
 �? 
   ����B�[E`��A�[�L�
|���;�C���E��o�������3�T0 k� ������U8D"!U2d  
 ��? 
   ����B�\E`��A�[�L�
|���;�C���E��o�������3�T0 k� ������U8D"!U2d   ��? 
   ����B�]E`��A�W�L�
|���;�C���E��n�������3�T0 k� ������U8D"!U2d   ��?
   ����B�]E`��A�S�L�
����;�C���E��m�������3�T0 k� ������U8D"!U2d   ��? 
   ����B�^A���A�O�L�
����;�C��E��m�������3�T0 k� ������U8D"!U2d   ��? 
   ����B�_A���A�O�L�
���;�C�{�E��l��������3�T0 k� ������U8D"!U2d   ��? 
   ����B                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��X ]� � �� j~Z    9     ��
	     j��
#f    ���s   
                 6          �      ���   (
	         ��ו   Q       ���>,    ��ۑ��J     ���L   
                 7�        ��     ���   8
�           ���-         �g�4    �����g�4     &                     D         �      ���   	@	
           R   $ $      �/�     R�/:                         �$          ��     ���   H
$
         ���]         .�[%J    ���]�[%J                          ���$          �       ���   H
	!          		�  ��
     B���     	6���     4                      ���7              X  ���    0          ��9 � �
    V�6�W    ��9�6��      �                d ���B          ���    ��`   8	          ��� 5 5	     j�C	�    �����C	�    ��                	���B         ��    ��@   0
%           ���s    	   ~�Do�    ��&�D�+    �}�'                 ���B�        �      ��H   0	          ��Z(  ? ? 
	   ��LMA    ��c�LMA                        O	���B         	 ���    ��@   8         ���  � �	   ��gZ    ���^�h`"    �$�                 ���B         
 p�     ��`   P
		          B ��     � �?�     B �?�                             ���q             �  ��@    P                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          w}'  ��        ��Q�     w~��[X    ���s "                  x                j  �        �                          w    ��        ��       w  �                                                               �                         �
���g�/�[��6�C�D�L�g �����     
     	        
    j �5  ���N       $� �r@ %� s@ �d  u� ɤ  v  �� v` $d s ���J ����X � d n� �D s� �d s����< ����J ����X � �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0� ���� ����� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����B������ �  ������  
�fD
��L���"����D" � j  "  B   J jF�"    "�j * , ����
��"     �j @�    �
� �  �  
�  j    ��     ��
       j    ��     ��
      ����  ��     ��D          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �       ��t(  ��        �T ���        �        ��        �        ��        �   f�     ��� v �        ��                         ���    ����                                     �                 ����              j�
 ���%��  ���B��                18 Craig Simpson n y   4:58                                                                        2  2      �
"�b$�$$�;CB=CD< CL4 �C5 � C"- �	kV � �
k\ � �k` � �kj � � kr � �ks � �c~ � � c� � �c� � � c� � �C. � � C6 � �K � � K � �c� � � c� � �c� � �c� � � c� � �"� � � "� � �� � �
� � z "* | �!"2 | � ""@ | �#": � � $"P � �%!� �&"* |'"< �"("2 |:)"6 |:*"
 �B +"L �Z  "R �Z  "C �:."6 |B /" �B  "D �B  "D �B 2" �B  "D �:4"6 |B 5" �B  "D �I  "D �]  "R �A 9"D �Y  "R �U  " �=<"< �E="2 |]>"6 |] "
 �                                                                                                                                                                                                                         �� P         �     @ 
        _     U P E X  ��                     	�������������������������������������� ���������	�
��������                                                                                          ��    ��a�� ��������������������������������������������������������   �4, ,    m�� �	�A ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	        `    (     �  H�J                                     ������������������������������������������������������                                                                                                                                               �        �      �        �    ��              
 	  
	 
 	 	 � ��� �� �����������  �������� ���� �������� ��������������������������� ������������������� �������������� �������������������������� ����������   � ������� ������������ �������������������  ��������������������������� �������������                                     *    *    ��  D�J    	 �9  	                           ������������������������������������������������������                                                                       	                                                                    �      �      �        �        �  �          	  
 	 
 	 	 ��������� ������ � ���� �������� � ���� �������������� ��������������������������������������������������������������� ��������������������������������������������� ��  �������������� �������� �������� �������� ������������ ������ ��� ��������                                                                                                                                                                                                                                                                                                                   
        �             


           �   }�         ������������������������������������    ����������������  '���������������������������������������������                                                                                �ww�ww333wwwwwwww�ww�ww�ww�ww333wwww I @ 5 
               	                 � o<�Q �\                                                                                                                                                                                                                                                                                         	n)h
  Y        c      c                  `      m      k                       ��                                                                                                                                                                                                                                                                                                                                                                                       �  � ��  � @��  � ��  � (��  � ��  ��8�n����������������J�����F�����y�����������          .   �� ����	       	  	�   & AG� �   X   
           �f�                                                                                                                                                                                                                                                                                                                                      p C B   �      ��        "         !��                                                                                                                                                                                                                        Y��   �� � Ѱ��      �� @      � ��� �� �����������  �������� ���� �������� ��������������������������� ������������������� �������������� �������������������������� ����������   � ������� ������������ �������������������  ��������������������������� ���������������������� ������ � ���� �������� � ���� �������������� ��������������������������������������������������������������� ��������������������������������������������� ��  �������������� �������� �������� �������� ������������ ������ ��� ��������   �� �     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    8      5      w                       e     �   �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$     �      �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@      
h> ��   
h> �$ ^$  �� � ��� �� � ��� �$  � �  �� �  �      �       ���� e�����  g���        f ^�         �� v��            ��Xn���2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �   3       �  �3 3�=������<��̼��� �3 33==ƙ�<ə�ƙ�3ƙ��ƙ���i� 3= ��3=�l�ә��<��l<��l<��l<���<    �   3=  �30 ��� ���=��������                        +   3     0  �<  3� 3� =� =� 0� 0������������������3�33033�0�3�0��;f��;��̽�������3��3��<���<�f���̳=�=�������3303<�<00�<30�3����������������=��=��3�3�=�3�0  �=  �3  �3� ��0 ̳0 �0 �0  0� =� =� 3�  3�  �<  0  33�0�3�0�3�0�3303�303�303�303303��<���0<��0<033<033003300330033030�30�<00�<0330333033303330333033�0��<���0�03303303=03=03��0 ̳0 ��0 �3� �3� �=  0  3�     �                           <�03=��3=�� 3��  �=  �        033003300330�330��303= ��33    330333033303330333<��333ݰ    0=�0<3���;�3 �=  3�             �                           wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                                    �����   �   �   �   ����                                     	�  		  	 � 	 	 	   	   	   	   	  ��                  ��   	   	   	   	   	   	 	 	 � 		  	�                 �   	    �   	    �   	    �   	   	   �  	   �  	   �  	   �                                      
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           " """ "!   " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             " """ "!   " ""  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                        "! ""! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                                 ��	����ɪ�ܙ����ݼ "-� "� J.��#��C>Z�C U�D �Z�#�U"�C"�� ���                �  �˰ ̻� �wp ׶� �vp �w� ɪ� ��� ��� �ۙ ��� �
� �" 0�" 0.�@ "�            ����˰ + �"  "" "  � �     �  �  ��  �   �                 U   U  U  U  	T  ,� ,� "  " "  ��  �              �   � � �  ��� ��  �                    �                        ���� ��� ����                            ��  ��  ��� ���                                                                                                                                                                                             �U  EU  U  3  ��  ��  �   �   �   �                   U�  U�@ EZ� 4Z� 3ZS U� E����" ��� 
��  �" ""�"" �"!  �  �                        "  "/  "��� "  !��  ���  �       �  ��  ̽  ��  �w  �� 
�� ��� ��� ��� ��� ��� ��� ��� �� ���    �   �   �   �   �   ˰  ˙  ɪ  ��� ټ� �̰ �̰ ��� ��  ��                              ��    
�  ��  ��  ��  �����  �   �          ��                           � ��                    ���� �                                                                                                                                                                                        �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ��������  ��                            �   ���  ���  �                    �    ��                 � �  �  �                      �  �  �  �               ���                                                        ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                         �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �                     �    � �� �  �� 	  
  �  ",  ""  �"   "                      ��  ��  �          ���� ��� ����                            ��  ��  ���   ���� �                                                                                                                                                                                       �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                             �  ��� ��� ��� �ݪ�                       �   �    �z� 
�� ������������ ˍ� ��� ���������ˉ����� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��                    ˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                                         �  ��  �� ��  ��       �  � � �� ��     �         �   �                     �     �                                      � ����ݼ� ����                                                                                                                                                                ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                        "  .���"    �     �                                       �   ���                            �   �                                                                                                                �   �  �  �  ��  ��  C�  U=  UJ  DZ  D  E  �4 
�: ���+��"��""� """ ""   �   �                        ɪ��ɪw̚�p�������������˻��۽��ݸ�̲-ۻ"""�""�2"�@  �C  �D  �T  D@  �   �   �   "�  "     �� �  �                                        ܰ ˻ �ݚ��w{`  g`  w                      �  �  ��"� ��� "               ����   �       �                                   �    ���  ��                    ��  ��  ���  �   ��  ��  ��  �  �   ��  ��                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  �   �   �   �   �       �     �"  "  �   "                                    �   �   �            �� �� �� g} �� vw                     �    � �  ��                  ���                � �������������  �                                                                                                                                          	��ˋ����۪��ۚ{Ƚ�g˽˖�-��"�� .� 
�8 
�� 
D> DC �D0 �D 
�C U@ �� 	�� ��" , " "/ "/� �� �   �                    �   ��  ��  w�  k�� g�� w�� ��� �۹ ��� ��� 3̰ �  >�" 2� 2"�DC �3  ��  ��  +   "   "   "/� ��     �                               �  �� �  �  �   �     ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                     ��  ��  ���                   ���                                                                                                                                                                             �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                                 ���                                                                                                                                                                                                   �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    DD@DD@                        �� ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(����������������� � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(����������������� 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5���������������� x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x���������������� w w x y�������H���������������������������������H������yxww����������������  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(���������������� , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,���������������� +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+���������������� 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5���������������� =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=����������������     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( ���������������� � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � ����������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq
"�b$�$$�;CB=CD< CL4 �C5 � C"- �	kV � �
k\ � �k` � �kj � � kr � �ks � �c~ � � c� � �c� � � c� � �C. � � C6 � �K � � K � �c� � � c� � �c� � �c� � � c� � �"� � � "� � �� � �
� � z "* | �!"2 | � ""@ | �#": � � $"P � �%!� �&"* |'"< �"("2 |:)"6 |:*"
 �B +"L �Z  "R �Z  "C �:."6 |B /" �B  "D �B  "D �B 2" �B  "D �:4"6 |B 5" �B  "D �I  "D �]  "R �A 9"D �Y  "R �U  " �=<"< �E="2 |]>"6 |] "
 �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.����������������������������������������� ��=�K�X�X�_��B�G�Q�K� � � � � � � � � � �2�0�.�����������������������������������������#��-�X�G�O�M��<�O�S�V�Y�U�T� � � � � � � �/�.�7�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������2�0�.� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������/�.�7� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                