GST@�                                                            \     �                                               �����      �      "         �������J���ʰ������������������         i     #    ����                                d8<n    �  ?     �����  �
fD�
�L���"����D"� j   " B   J  jF�"     "�j  " ���
��
�"    B�jl �   B ��
   �                                                                              ����������������������������������      ��    bb= QQ0 4 111 44              		 

                     ��� �   � �                 nn ))
         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                ��  �       �   @  #   �   �                                                                                '     )n)n
  �    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE * �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    C�8s3���<E�$�S��+����B��c����3�<Z��T0 k� �ǜ�˜'$2(u e1�t A  ��    ��� �C�4s?���<E#W��+����B��c����2�<Z��T0 k� �˝�ϝ'$2(u e1�t A  ��    ��� �E�0sO���<E!c��+��ϔB��c����/�@Z��T0 k� �מ�۞'$2(u e1�t A  ��    ��� �E�,sW���<E g�+��הB��c��	��-�DZ��T0 k� �۟�ߟ'$2(u e1�t A  ��    ��� �E�(	s_���<E o�+��ۓB��c����,�DZ��T0 k� ����'$2(u e1�t A  ��    ��� �E�$sg���<E(s�+���I�c��� +�HZ��T0 k� ����'$2(u e1�t A  ��    ��� �E� sk���<B�0{�+�q�I�c���)�LZ��T0 k� ����'$2(u e1�t A  ��    ��� �E�ss���<B�8��+�q�I�c�� �(�LZ��T0 k� �����'$2(u e1�t A  ��    ��� �E��s����=B�H���+�q��I�c�� � %�PZ��T0 k� ������'$2(u e1�t A  ��    ��� �E��c����=B�P���+�r�I" c	����($�TZ��T0 k� �����'$2(u e1�t A  ��    ��� �E��c����=B�T����+r�I"c	����($�TZ��T0 k� ����'$2(u e1�t A  ��    ��� �E��c��� =B�\����+r�I"c	����,#�XZ��T0 k� ����'$2(u e1�t A  ��    ��� �E��c���=B�l����+~r#�I"c	����8!�`Z��T0 k� ����'$2(u e1�t A  ��    ��� �E��c���=B�t����+}�'�I c	����@!�dZ��T0 k� ����'$2(u e1�t A  ��    ��� �E��c��� =B�|����+}�/�I(c	����H �dZ��T0 k� ���#�'$2(u e1�t A  ��    ��� �E��c���(=B������+|�7�I,c	����L�hZ��T0 k� �#��'�'$2(u e1�t A  ��    ��� �E��c���0=B������+|�;�I0c	����T�lZ��T0 k� �+��/�'$2(u e1�t A  ��    ��� �E��cÒ�@=B������+{�G�I<c	����`�pZ��T0 k� �3��7�'$2(u e1�t A  ��    ��� �C��cǑ�H=B������+{�O�I"@c���hstZ��T0 k� �7��;�'$2(u e1�t A  ��    ��� �C��cː�P=B������+z�S�I"Dc���psxZ��T0 k� �?��C�'$2(u e1�t A  ��    ��� �C��SϏ�X=B������+z�[�I"Hc���tsxZ��T0 k� �C��G�'$2(u e1�t A  ��    ��� �C��SӍ�`=B������+y�_�I"Lc��s|s|Z��T0 k� �G��K�'$2(u e1�t A  ��    ��� �C��S׌�h=B������+y�c�I"Pc��s�s�Z��T0 k� �K��O�'$2(u e1�t A  ��    ��� �C��Sۋ�p=B�����+x�k�ITc��s�s��Z��T0 k� �S��W�'$2(u e1�t A  ��    ��� �C���S߉��=B�����+x�s�I\c��s�s��Z��T0 k� �[��_�'$2(u e1�t A  ��    ��� �C���S���=B�����+w�{�I\c��s�s��Z��T0 k� �_��c�'$2(u e1�t A  ��    ��� �C���S���=B���#��+w��I`c��s�s��Z��T0 k� �g��k�'$2(u e1�t A  ��    ��� �C���S���=B���+��+v҃�I"dc��s�s��Z��T0 k� �k��o�'$2(u e1�t A  ��    ��� �C���S���=B��
�3��+vҋ�I"hc���s�c��Z��T0 k� �o��s�'$2(u e1�t A  ��    ��� �C���C���=B� 
�;��+vҏ�I"hc���s�c��Z��T0 k� �s��w�'$2(u e1�t A  ��    ��� �C���C���=I	�C��+uғ�I"lc���s�
c��Z��T0 k� �{���'$2(u e1�t A  ��    ��� C���C���=I	�G��+ur��I"lc���s�	c��Z��T0 k� �����'$2(u e1�t A  ��    ��� C���C���=I�O��+tr��Ipc���c�c��Z��T0 k� ������'$2(u e1�t A  ��    ��� E���C���=I �_��+tr��Ipc���c�c��Z��T0 k� ������'$2(u e1�t A  ��    ��� E���C���=I $�g��+sr��Itc���c�c��Z��T0 k� ������'$2(u e1�t A  ��    ��� E���3���=I ,�o��+sr��Itc���c�c��Z��T0 k� ������'$2(u e1�t A  ��    ��� E���3���=I 0�w��+s�I"tc���c��c��Z��T0 k� ������'$2(u e1�t A  ��    ��� E���3���=I 4���+r�I"xc���c��c��Y���T0 k� ������'$2(u e1�t A  ��    ��� E�þ3߈�>I@Ϗ��+r�ØI"xc���c��c��Y���T0 k� ������'$2(u e1�t A  ��    ��� Eѻ�3߈�>IDϗ��+q�ǗI"xc���c��c��Y���T0 k� ������'$2(u e1�t A  ��    ��� Eѷ�3߉�>ILϟ��+q�˗Ixc���c��c��Y���T0 k� ������'$2(u e1�t A  ��    ��� E᯹#ߊ�>IPϧ�@+q�ϗIxc������c��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� E᣶#ߋ�,>I \Ϸ�@�xrזIxc������c��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� E៵#ߌ�4>I dϿ�W��xrەIxc������S��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� Eᗳ#ۍ�<>I h���W��xrߔ@xc������S��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� Eᓲ�ߎ�D>I p���W��xr�@xc������S��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� Eዱ�ߏ�L>I x���W��xr�@xc������S��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� E���ߑ�\>B�����W��xr�@xc�����S��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� D1w��ߒ�d>B�����W��xr�@bxc�����S��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� D1o��ߓ�l>B�����W��xb��@bxc�����S��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� D1k��ߔ�t>B����W��xb��@bxc�����S��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� D1[��ߖ��>B����W��xb��@bxc�����S��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� E�S��ߘ��>B����W��xc�@bxc�����S��Y���T0 k� ������'$2(u !ae1�t A  ��    ��� E�K��ߙє>B���#�W��xc�@bxcB#����C��Y���T0 k� �����'$2(u !ae1�t A  ��    ��� E�G��ߚѠ>B���+�W��xc�@bxcB'����C��Y���T0 k� ����'$2(u !ae1�t A  ��    ��� E�?�ߜѨ>B���3�W��xc�@bxcB+����C��Y���T0 k� ����'$2(u !ae1�t A  ��    ��� E�7�ߝѰ>B���;�W��xc�@bxcB/����C��^���T0 k� ����'$2(u !ae1�t A  �    ��� E�/�ߞѸ>B���C�W��xc�@bxcB3����C��^���T0 k� ����'$2(u !ae1�t A  �    ��� E�'�ߠ��>B���K�W��xc�@bxc �7����C��^���T0 k� ����'$2(u !ae1�t A  ��    ��� E��ߢ��>E���_�W��xc�@bxc �?����C��^���T0 k� ����'$2(u !ae1�t A  ��    ��� E��ߣ��>E���g�W��xc�@bxc �C����C�_���T0 k� ����'$2(u !ae1�t A  ��    ��� E��ߥ��>E��o�W��xc�@bxc �C����{�_���T0 k� ����'$2(u !ae1�t A  ��    ��� E���ߦ��=E��w�W��x��@bxc �G����{�_���T0 k� ����'$2(u !ae1�t A  ��    ��� E���ߧ��=E���W��x��@bxc �K����w�_���T0 k� ����'$2(u !ae1�t A  ��    ��� E��ߨ��=E����W��x��@bxc �O���w�_���T0 k� ����'$2(u !ae1�t A  ��    ��� E��#ߩ� =E�$���W��x��@bxc �S���s�_���T0 k� ������'$2(u !ae1�t A  ��    ��� E��#ߪ�=B�,���W��x��@bxc �W���o�_���T0 k� ������'$2(u !ae1�t A  ��    ��� E�ۧ#߬�<B�4���W��x��@bxc �W���o�_���T0 k� ������'$2(u !ae1�t A  �    ��� E�ק#߭�<B�< ���W��x��@bxc �[���k�_���T0 k� ������'$2(u !ae1�t A  ��    ��� E�ק#߮� <B�D ���W��x��@�xc �_���k�_���T0 k� ������'$2(u !ae1�t A ��    ��� E�צ#߯�(;B�O����W��x��@�xc �c���g�[���T0 k� ������'$2(u !ae1�t A ��    ��� F ӥ#߰�0;B�W����W��x�#�@�xc �g���g�[���T0 k� ������'$2(u !ae1�t A ��    ��� F Ϥ#߱�8;B�_����W��x�#�@�xc �g���c�[���T0 k� ������'$2(u !ae1�t A ��    ��� F Ϥ#߲�@:B�g��ǷW��x�#�@�xc �k���c�[��T0 k� ������'$2(u !ae1�t A ��    ��� F ϣ#߳�H:B�o��˸W��x�#�Axc �o���_�[��T0 k� ������'$2(u !ae1�t A ��    ��� F ˢ#ߴrP9B�w��ӸW��x�'�Axb �o���_�[��T0 k� ������'$2(u !ae1�t A ��   ��� F ˢ#ߵrX9B���۹W��x�'�Axb �s���[�[��T0 k� ������'$2(u !ae1�t A ��    ��� F ˡ#߶r`8B���߹W��x�'�Axb �w���[�[��T0 k� ����'$2(u !ae1�t A ��    ��� E�ˡ#߷rh8C����BO�x�+�Axb �w���W�[��T0 k� ����'$2(u !ae1�t A ��    ��� E�ˠ#߸rp8C����BO�x�+�C�xb �{���W�[��T0 k� ����'$2(u !ae1�t A ��    ��� E�ˠ߸rx7C����BO�x�+�C�xb ����S�[��T0 k� �|
��
'$2(u !ae1�t A ��    ��� E�ˠ߹r|7C�����BO�x�+�C�ta ����S�[��T0 k� �t�x'$2(u !ae1�t A ��    ��� E�˟ߺr�6C�����BO�x�/�C�ta �����O�[��T0 k� �l�p'$2(u !ae1�t A ��    ��� B�˟߻r�6C����@�x�/�C�ta �����O�[��T0 k� �d�h'$2(u !ae1�t A ��    ��� B�˞߼r�6C����@�x�/�C�p` �����O�[��T0 k� �\�`'$2(u !ae1�t A ��    ��� B�˞߽r�5C����@�x�3�Ap` �����K�[��T0 k� �T�X'$2(u !ae1�t A ��    ��� B�ϝ߾r�5C����@�x�3�Al_ �����K�[��T0 k� �L�P'$2(u !ae1�t A ��    ��� B�ϝ߾r�4C����@�x�3�Al_ �����K�[��T0 k� �D�H'$2(u !ae1�t A ��    ��� B�ӝ߿r�4C����B��x�3�Al_ �����G�[��T0 k� �<�@'$2(u !ae1�t A ��    ��� B�Ӝ����4C���'�B��x�3�Ah^ �����G�[��T0 k� �4!�8!'$2(u !ae1�t A ��    ��� B�ל�����3C���+�B��x�3�Ah^ �����G�[��T0 k� �,#�0#'$2(u !ae1�t A ��    ��� B�ۛ�����3C���/�B��x�3�Ad] �����G�[��T0 k� �$&�(&'$2(u !ae1�t A ��    ��� B�ۛ�����3C���3�B��x�3�Ad] �����G�[��T0 k� �(� ('$2(u !ae1�t A ��    ��� B�ߛ�����2C��;�B��x�3�Ad] �����C�[��T0 k� �+�+'$2(u !ae1�t A  ��    ��� B�������2C��?�B��x�3�A`\ �����C�[��T0 k� �-�-'$2(u !ae1�t A  ��    ��� B�������2C��C�B��x�3�A`\ �����C�[��T0 k� �0�0'$2(u !ae1�t A  ��    ��� B�������1C��G�B��x�7�A`\ �����C�[��T0 k� ��2� 2'$2(u !ae1�t A  /�    ��� B�������1C#��K�B��x�7�A\[ �����C�[��T0 k� ��5��5'$2(u !ae1�t A  $�    ��� B�������1C+��S�B��x�7�A\[ �����C�[��T0 k� 2�5��5'$2(u !ae1�t A  ��    ��� B��������0C3��W�B��x�7�A\[ �����?�[��T0 k� 2�6��6'$2(u !ae1�t A  ��    ��� B��������0C"7��[�B��x�7�AXZ �����?�[��T0 k� 2�6��6'$2(u !ae1�t A  ��    ��� B��������0C"?��_�B��x�7�AXZ �����?�Zd�T0 k� 2�6��6'$2(u !ae1�t A  ��    ��� B�������/C"G��c�B��x�7�AXZ �����?�Zd�T0 k� 2�6� 6'$2(u !ae1�t A  ��    ��� B������/C"O��g�B��x�7�ATY �����?�Zd�T0 k� ��7� 7'$2(u !ae1�t A  ��    ��� B������/C"W��k�B��x�7�ATY �����?�Zd�T0 k� ��7� 7'$2(u !ae1�t A  ��    ��� B������/C"_��o�B��x�7�ATY �����?�Zd�T0 k� � 7�7'$2(u !ae1�t A  ��    ��� B������.C"g��s�B��x�7�APX �����;�Zd�T0 k� �5�5'$2(u !ae1�t A  ��"    ��� B������.C"k��w�B�x�7�APX �����;�Zd�T0 k� �2�2'$2(u !ae1�t A  ��"    ��� B�'�����.C"s��{�B�x�7�APX �����;�Zd�T0 k� �1�1'$2(u !ae1�t A  ��"   ��� B�+����� .C"{���B�x�7�APX �����;�Zd�T0 k� �0�0'$2(u !ae1�t A  ��"    ��� B�3�����$-C"�����B�x�7�ALW �����;�Zc��T0 k� �.� .'$2(u !ae1�t A  ��"    ��� B�;�����(-B�����B�x�;�ALW �����;�Zc��T0 k� � -�$-'$2(u !ae1�t A  ��"   ��� B�?�����,-B�����B�x�;�ALW �����;�Zc��T0 k� �$-�(-'$2(u !ae1�t A  ��"    ��� B�G�����4-B�����B�#x�;�AHW �����;�Zc��T0 k� �(-�,-'$2(u !ae1�t A  ��"    ��� B�O�����8,B�����B�'x�;�AHV �����7�Zc��T0 k� �,,�0,'$2(u !ae1�t A  ��"    ��� B�W�����<,B�����B�+x�;�AHV �����7�Zc��T0 k� �0,�4,'$2(u !ae1�t A  ��"    ��� B�_�����@,B�����B�3x�;�AHV �����7�Zc��T0 k� �4,�8,'$2(u !ae1�t A  ��"    ��� B�c�����D,B�����B�7x�;�ADU �����7�Zc��T0 k� �8,�<,'$2(u !ae1�t A  ��"    ��� B�k�����H+B�����B�?x�;�ADU �����7�Zc��T0 k� �<+�@+'$2(u !ae1�t A  ��"    ��� B�s�����L+B�����B�Cx�;�ADU �����7�Zc��T0 k� �@*�D*'$2(u !ae1�t A  ��"    ��� B�{�����P+B������B�Kx�;�ADU �����7�Zc��T0 k� �D*�H*'$2(u !ae1�t A  ��"    ��� Bу�����T+B������B�Ox�;�A@U �����7�Zc��T0 k� �H*�L*'$2(u !ae1�t A  ��"    ��� Bы�����X+B������B�Wx�;�A@T �����7�Zc��T0 k� �L*�P*'$2(u !ae1�t A  ��"    ��� Bї�����\*C�����B�_x�;�A@T �����3�Z���T0 k� �P)�T)'$2(u !ae1�t A  ��"    ��� Bџ����\*C�����B�cx�;�A@T �����3�Z���T0 k� �T)�X)'$2(u !ae1�t A  ��"    ��� B������`*C�����B�kx�;�A@T �����3�Z���T0 k� �X)�\)'$2(u !ae1�t A  ��"    ��� B������d*C�����B�sx�;�A<S �����3�Z���T0 k� �\)�`)'$2(u !ae1�t A  ��"    ��� B������h*C�����B�wx�;�A<S �����3�Z���T0 k� �`)�d)'$2(u !ae1�t A  ��"    ��� B�Ñ���l)C�����B�x�;�A<S �����3�Z���T0 k� �d(�h('$2(u !ae1�t A  ��"    ��� B�ːS���p)C�����B��x�;�A<S �����3�Z���T0 k� �h(�l('$2(u !ae1�t A  ��"    ��� B�ӐS��st)C�����B��x�?�A<S �����3�Z���T0 k� �l(�p('$2(u !ae1�t A  ��"    ��� B�ߐS��sx)C�����B��x�?�A8R �����3�Z���T0 k� �l(�p('$2(u !ae1�t A  ��"    ��� B��S��sx)C����B��x�?�A8R �����3�Z���T0 k� �p(�t('$2(u !ae1�t A  ��"    ��� B��S��s|(C����B��x�?�A8R �����/�Z���T0 k� �t(�x('$2(u !ae1�t A  ��"    ��� B������s�(C����B��x�?�A8R �����/�Z���T0 k� �x'�|''$2(u !ae1�t A  ��"    ��� B�����s�(C����B��x�?�A8R �����/�Z���T0 k� �|'��''$2(u !ae1�t A  ��"    ��� B�����C�(C����B��x�?�A4Q �����/�Z���T0 k� ��#��#'$2(u !ae1�t A  ��"    ��� B�����C�(C'����B��x�?�A4Q �����/�Z���T0 k� �� �� '$2(u !ae1�t A  ��"    ��� B�����C�(C+����B��x�?�A4Q ����/�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B�'����C�'C3����B��x�?�A4Q ����/�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B�3����C�'C;����B��x�?�A4Q ����/�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B�;����C�'CC����B��x�?�A4Q ����/�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B�C����C�'CK����B��x�?�A0P ����/�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B�O����C�'CS����B��x�?�A0P ����/�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B�W����C�'CW����B��x�?�A0P ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B�_����C�'C#_����B��x�?�A0P ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B�k����C�&C#g����B��x�C�A0P ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B�s����C�&C#o����B�x�C�A0P ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B�{����C�&C#w����B�x�C�A,P ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B����C�&C#{����B�x�C�A,O ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B����C�&C#����B�x�C�A,O ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B����C�&C#����B�#x�C�A,O ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� B£����C�&K�����B�+x�C�A,O ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� E������C�&K�����B�/x�C�A,O ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"   ��� E������C�%K�����B�7x�C�A,O ����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� E������C�%K�����B�?x�C�A,O �����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� E�ǌ���C�%K����#�B�Gx�C�A(N �����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� E�Ӎ���C�%K����'�B�Kx�C�A(N �����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� E�ۍ���C�%K����/�B�Sx�C�A(N �����'�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� E�����C�%K����3�B�[x�C�A(N �����'�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� E�����C�%K����7�B�cx�C�A(N �����+�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Lr����C�%K����?�B�gx�C�A(N �����/�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Lr����C�$K����C�B�ox�C�A(N �����3�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Lr����C�$K�ò�K�B�wx�C�A(N �����7�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Lr����C�$K�Ǳ�O�B�x�C�A$M �����7�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Lr����C�$K�˰�W�Bуx�C�A$M �����;�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Lr����C�$K�Ϯ�_�Bыx�G�A$M �����?�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Ls���C�$K�ӭ�c�Bѓx�G�A$M �����C�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Ls���C�$K�׬�k�K��x�G�A$M �����C�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Ls���C�$K�۫�s�K��x�G�A$M �����G�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Ls���C�$K�ߪ�w�K��x�K�A$M ����K�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Ls���C�$K����K��x�K�A$M ����K�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Ls���C�#K��҇�K��x�O�A$M ����O�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Ls���C�#K��ҋ�K��x�O�A M ����S�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� Ls���C�#K��ғ�K��x�S�A L ����S�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� L����C�#K��қ�K��x�S�A L ����W�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� L����C�#K��ң�K��x�S�A L ����[�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� L����C�#K������K��x�W�A L ����[�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� L����C�#K������K��x�W�A L ����_�Z���T0 k� ����'$2(u !ae1�t A  ��"    ��� L����C�#K������K��x�[�A L ����_�Z���T0 k� ��� '$2(u !ae1�t A  ��"    ��� L����C�#K������K��x�[�A L ����c�Z���T0 k� ��� '$2(u !ae1�t A  ��"    ��� L����C�#K�����K��x�_�A L ����g�Z���T0 k� ��� '$2(u !ae1�t A  ��"    ��� L����C�#K�����K��x�_�A L ����g�Z���T0 k� � �'$2(u !ae1�t A  ��"   ��� L����C�#K�����K��x�_�A L ����k�Z���T0 k� � �'$2(u !ae1�t A  ��"    ��� L�#���C�#K�����K��x�c�A L ����k�Z���T0 k� � �'$2(u !ae1�t A  ��"    ��� L�#���C�"K�����K��x�c�AK ����o�Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�'���C�#K�����K�x�g�AK ����o�Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�'���C�#K�����K�x�g�AK ����s�Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�'���C�#K�����K�x�g�AK ����s�Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�+���C�$K����K�x�k�AK ����w�Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�+���C�$K����K�x�k�AK ����w�Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�+���C�$K����K�x�k�AK ����{�Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�/���C�%K����K�x�o�AK ����{�Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�/���C�%K�#��#�K�#x�o�AK �����Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�/���C�%K�#��+�K�'x�s�AK �����Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�3���C�&K�'��3�K�/x�s�AK ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�3���C�&K�+��;�K�3x�s�AK ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�7���C�&K�+��C�K�7x�w�AK ������Z���T0 k� ��'$2(u !ae1�t A  ��"   ��� L�7���C�&K�/��K�K�;x�w�AK ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�7���C�'K�/��S�K�?x�w�AK ������Z���T0 k� ��'$2(u !ae1�t A  ��"   ��� L�7���C�'K�3��[�K�Cx�{�AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�;���C�'K�7��k�K�Kx�{�AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�;���C�(K�7��s�K�Ox�{�AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�;���C�(K�7��{�K�Sx��AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�;���C�(K�3���K�Wx��AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�;���C�)K�3���K�[x��AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�;���C�)K�3���K�_x���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�?���C�)K�3���K�cx���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�?���C�)K�3���K�gx���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�?���C�*K�3���K�gx���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�?���C�*K�3���K�kx���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�C���C�*K�3��K�ox���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�C���C�*@/��þK�sx���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�C���C�+@/��˽K�wx���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� L�C�C�C�+@/�	�ӽK�{x���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� LsG�C�C�+@/�	�ۼK�x���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� LsG�C�C�+@/�	�ۼK�x���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� LsG�C�C�+E�/�	��K��x���AJ ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� LsG�C�C�,E�/�	��K��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� LsG�C�C�,E�/�
�K��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� LsK�C�C�,E�/�
�K��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�K�C�C�,E�/�
��K��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�K�C�C�,E�/�
��K��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�K�s�C�-Et/�
��K��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�O�s�C�-Et/���K��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�O�s�C�-Et/���K��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�S�s�C�-Et/���B��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�S�s�C�-Et/���B��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�W�s�C�.Et/���B��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�W�s�C�.Et/���B��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�[�s�C�.LT/���B��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�[�s�C�.LT/�t#�B��x���AI ������Z���T0 k� ��'$2(u !ae1�t A  ��"    ��� D�[�s�C�.LT/�t'�B��x���AI ������Z���T0 k� � � '$2(u !ae1�t A  ��"    ��� D�[�s�C�/LT/�t+�B��x���AI ������Z���T0 k� � � '$2(u !ae1�t A  ��"    ��� D�_�s�C�/LT/�t/�E��x���AI ������Z���T0 k� � � '$2(u !ae1�t A  ��"    ��� D�_�s�D /LT/�t3�E��x���AI ������Z���T0 k� � � '$2(u !ae1�t A  ��"    ��� D�c�s��D /LT/�t7�E��x���AI ������Z���T0 k� � � '$2(u !ae1�t A  ��"    ��� D�g����D /LT/�t?�E��x���AI ������Z���T0 k� � � '$2(u !ae1�t A  ��"    ��� D�g����D /LT/�tC�E��y���AI ������Z���T0 k� �!�!'$2(u !ae1�t A  ��"    ��� D�g����D 0LT/�tG�E��y���AI ������Z���T0 k� �!�!'$2(u !ae1�t A  ��"    ��� D�k����D 0LT/�tK�E��y���AI �#�����Z���T0 k� �!�!'$2(u !ae1�t A  ��"    ��� D�k����D 0LT/�tO�E��y���AI �#�����Z���T0 k� �!�!'$2(u !ae1�t A  ��"   ��� D�o����D 0LT/�tS�E��z���AI �#�����Z���T0 k� �!�!'$2(u !ae1�t A  ��"    ��� D�s����D 0Ld/�tW�E��z���AI �#�����Z���T0 k� �!�!'$2(u !ae1�t A  ��"    ��� D�w����D 0Ld/�t[�D��z���AI �#�����Z���T0 k� �!�!'$2(u !ae1�t A  ��"    ��� D�{����D 0Ld/��[�D��{���AI �#�����Z���T0 k� �"�"'$2(u !ae1�t A  ��"    ��� D�{����D 1Ld/��_�D��{���AI �#�����Z���T0 k� �"�"'$2(u !ae1�t A  ��"    ��� D�����D 1Ld/��c�D��|���AH �#�����Z���T0 k� �"�"'$2(u !ae1�t A  ��"    ��� D����D 1Ld/��g�D��|���AH �#�����Z���T0 k� �"�"'$2(u !ae1�t A  ��"    ��� E������t 1Ld/��k�D�}���AH �#�����Z���T0 k� �%�%'$2(u !ae1�t A  ��"    ��� E� o�	� QCL�d�;�����E;�O	��%O����bs� T0 k� ��%� %'$2(u e1�t A  ��U    � 	�8E� s�	�PCL�d� =�����E;�N	��%O����
bs� T0 k� ��%� %'$2(u e1�t A  ��U    � 	�8E�$w�	�OCL�b�(?�����E;pL	��%O����bs� T0 k� ��%� %'$2(u e1�t A ��U    � 	�8B�$w�	�NE<�a	\(?�����E;hK	��%O����bs� T0 k� ��%� %'$2(u e1�t A ��U    � 	�8B�({�	�NE<�`	\,@�����E;lI	��%O����bs� T0 k� ��%��%'$2(u e1�t A  ��U    � 	�8B�(�	��ME<x_	\0@�����E+lH	��%O����bs� T0 k� ��&��&'$2(u e1�t A  ��U    � 	�8B�,�	��ME<t^	\0A�����E+lF	��%O����bs� T0 k� ��%� %'$2(u e1�t A  ��U    � 	�8B�0"��	��LE<h\	\4B�����E+lC	��%O�����bs� T0 k� ��$� $'$2(u e1�t A  ��U    � 	�8E�4$��	��LE<dZ	l8C�����E+pA	��%?�����Z3� T0 k� ��#� #'$2(u e1�t A  ��U    � 	�8E�8&��	��LE<`Y	l8D�����E+p?	��%?����Z3� T0 k� ��#� #'$2(u e1�t A  ��U    � 	�8E�<'���	��LE<XX	l8D{����E+p=	��%?����Z3� T0 k� ��'$2(u e1�t A  ��U    � 	�8E�@)���	��LE<TW	l<E{����E+t<	��%?����Z3� T0 k� ��'$2(u e1�t A  ��U    � 	�8E�H,���	��LE<TW	l<D| ۋ�E+x8	��%?s���Z3� T0 k� ��'$2(u e1�t A  ��U    � 	�8E�L.���	��LI\PWL<D| ۏ�E+x6	��%?k���Z3� T0 k� ��'$2(u e1�t A  ��U    � 	�8E�T/���	��LI\LWL<C|ۏ�E+|4	��%?g���Z3� T0 k� ��'$2(u e1�t A  ��U    � 	�8E�X1���	��LI\HWL<C|ۏ�E+�3	��%?_���Z3� T0 k� �� '$2(u e1�t A  ��U    � 	�8E�`4���	��LI\DWL<C�ۓ�E�/	��%?O���Z3� T0 k� � �$'$2(u e1�t A  ��U    � 	�8E�h6ܻ���LI\@VL<C�ۗ�E�-	��%?G���Z3� T0 k� �,�0'$2(u e1�t A  �U    � 	�<E�l7ܿ���KIl@VL<C�ۗ�E�+	��%?C���Z3� T0 k� �4�8'$2(u e1�t A ��    � 	�@E�t8�����KIl<VL<C�ۛ�E�*	��%/;���Z3� T0 k� �@�D'$2(u e1�t A ��    � 	�DE��;�����KIl8VL<C�۟�E�&	��%//���Z3� T0 k� �X�\'$2(u e1�t A ��    � 	�HE��<����JIl8VL<C�ۣ�E�$��%/'���Z3� T0 k� �d �h '$2(u e1�t A ��    � 	�LE�>����JE,8V<C�맶E�#��%/#���Z3� T0 k� �p!�t!'$2(u e1�t A ��    � 	�PE�?����JE,4V<C�뫵E�!��%/���Z3� T0 k� �x#�|#'$2(u e1�t A ��    � 	�TE�@����IE,4V<C�뫴E���%/���Z3� T0 k� ��%��%'$2(u e1�t A ��    � 	�WE�B����IE,4V<C믲E���%/����Z3� T0 k� ��'��''$2(u e1�t A ��    � 	�ZE�C�����HE,0V<C볱E���%/����Z3� T0 k� ��)��)'$2(u e1�t A ��    � 	�]E�D�����HE,0V\<C 뷰E���%/����Z3� T0 k� ��+��+'$2(u e1�t A ��    � 	�`B��G����GE,0U\<C$뿭E����%.����Z3� T0 k� ��/��/'$2(u e1�t A ��    � 	�dB��H����GE,0U\<C$ëE���%����Z3� T0 k� ��1��1'$2(u e1�t A ��    � 	�hB��I����GE,0T\<C(ǪE���%����Z3� T0 k� ��3��3'$2(u e1�t A ��    � 
�kB��J����FB�0T\<C(˨E���%����Z3� T0 k� ��5��5'$2(u e1�t A ��    � �nB��K����FB�0T\<C�(ϧE����%����Z3� T0 k� ��7��7'$2(u e1�t A ��    � �qB��M�'���FB�0S�<C�,ӥD����%����Z3� T0 k� ��9��9'$2(u e1�t A ��    � �tB��N�+���EB�0S�<C�,ۤD�� ��%�����Z3� T0 k� � ;�;'$2(u e1�t A ��    � �wB��O�3���EB�0S�<C�0ߢD��"��%�����Z3� T0 k� �<�<'$2(u e1�t A ��    � �zB�Q�C���DB�0S�<B�0�D�%��%���#�Z3� T0 k� � @�$@'$2(u e1�t A ��    � �~B�R�K���DB�0R�<B�4�D�&��%���'�Z3� T0 k� �,B�0B'$2(u e1�t A ��    � ��B�S�S���DB�0R�<B�4��D�(��%���+�Z3� T0 k� �8D�<D'$2(u e1�t A ��    � ��B�$T�[���CB�4R�<A�4���D�$)��%���/�Z3� T0 k� �DF�HF'$2(u e1�t A ��    � ��B�,U�c���CB�4Q�<A�8���D�,*��%���3�Z3� T0 k� �PH�TH'$2(u e1�t A ��    � ��B�4V�k���CB�4Q�<@�8��D�4,��%���;�Z3� T0 k� �XJ�\J'$2(u e1�t A ��    � ��B�<W�s���BC8P�<@�<��D�<-�%���?�Z3� T0 k� �dL�hL'$2(u e1�t A ��    � ��B�DX�{���BC8P�<?�<��D�D/|%��	�C�Z3� T0 k� �pN�tN'$2(u e1�t A ��    � ��EXZ�����AC<O�<?�@��O�P/p%���K�Z3� T0 k� ��R��R'$2(u e1�t A �    � ��E`[�����AC<O�<?�@�#�O�X0l%���O�Z3� T0 k� ��T��T'$2(u e1�t A ��   � ��Eh\�����AE,<O�<?�@�'�O�`0d%���W�Z3� T0 k� ��V��V'$2(u e1�t A ��    � ��Ep]�����AE,@O�<?�@�/�O�h1O\%���[�Z3� T0 k� ��W��W'$2(u e1�t A ��    � ��Ex^�� ��@E,@O�<?�D�3�O�p1OX%���_�Z3� T0 k� ��Y��Y'$2(u e1�t A ��    � ��E�_�� ��@E,HO�<?�D�C�O��2OH&���k�Z3� T0 k� ��]��]'$2(u e1�t A ��    � ��E�`�� ��?EHO�<>�D�G�O��3OD&���o�Z3� T0 k� ��_��_'$2(u e1�t A ��    � ��E��a�� ��?ELN�<>�D�O�O��3O<&�� s�Z3� T0 k� ��a��a'$2(u e1�t A ��    � ��E��b����?EPN�<>�@�W�O��4O4&�� {�Z3� T0 k� ��c��c'$2(u e1�t A ��    �  ��E��c����?EPN�<>�@�_�O��4O,'�� �Z3� T0 k� ��e��e'$2(u e1�t A ��    � !��E��d����>ETN�<>�@�c�O��4O('�� ��Z3� T0 k� �g�g'$2(u e1�t A ��    � "��E��e����>B�XN�<=�@�k�O��5O '�� ��Z3� T0 k� �i�i'$2(u e1�t A ��    � #��E��f����>B�\N�@=�<�sO��5O(�  ��Z3� T0 k� �k�k'$2(u e1�t A ��    � $��E��g���>B�\N�@=�<�{�O��6O(� ��Z3� T0 k� �$m�(m'$2(u e1�t A ��    � %��E��h���>B�`N�D=�<��O��6?)� ��Z3� T0 k� �0o�4o'$2(u e1�t A  ��    � &��E��i���=B�`N�D=�<���O��6? *� ��Z3� T0 k� �<q�@q'$2(u e1�t A  -�    � '��BN�j�� =B�dN�H<�<���O��7>�*� ��Z3� T0 k� �Dr�Hr'$2(u e1�t A  ��    � (��BN�k�$�=B�dN�H<�<���O��7>�+� ��Z3� T0 k� �Pt�Tt'$2(u e1�t A  ��    � )��BN�k�0 �=B�hN�L<�<���O��8>�,���Z3� T0 k� �\v�`v'$2(u e1�t A  ��    � *��BO l�8 �=B�hN�L<�<���O��8>�-���Z3� T0 k� �hx�lx'$2(u e1�t A  ��    � +��BOm�@ �=B�hN�P<�<���O��8>�.���Z3� T0 k� �pz�tz'$2(u e1�t A ��    � ,��BOn�H �=B�hN�T;�<��O��9>�/�$õZ3� T0 k� �||��|'$2(u e1�t A ��    � -��BOo�S��=B�lM�T;�<��O��9>�0�(˵Z3� T0 k� ��~��~'$2(u e1�t A ��    � .��BOp�[��=B�lM�X;�<ǃO��9>�1�,ӵZ3� T0 k� ������'$2(u e1�t A ��    � /��BO$p�g��=B�lM�\;�<σO��:.�2�0׵Z3� T0 k� ������'$2(u e1�t A ��    � 0��BO(q�o��=B�pM�\;�8׃D��:.�3�8ߵZ3� T0 k� ������'$2(u e1�t A *�    � 1��BO0r�w��=B�pM�`;�8߄D� :.�5�<�Z3� T0 k� .�����'$2(u e1�t A ��    � 2��BO8s��� <B�tM�`:�8��D�;.�6�D �Z3� T0 k� .���ă'$2(u e1�t A  ��    � 3��BO<tއ�� <B�tL�d:�8��D�;.�7�H!�Z3� T0 k� .Ȃ�̂'$2(u e1�t A  ��    � 4��BOLuޛ��$<B�xL�l:�8��D�=.�:�T" ��Z3� T0 k� .����'$2(u e1�t A  .�    � 5��BOPv���(<B�|K�l:�8��D� =.�;�\"!�Z3� T0 k� .����'$2(u e1�t A  ��    � 6��BOXv���,<B�|K�p:�8��D�$>��<�d#!�Z3� T0 k� �����'$2(u e1�t A  ��    � 7��BO\w���0<B��K�t9�8��D�,>��>�h$!�Z3� T0 k� � ���'$2(u e1�t A  ��    � 8��BOdx���4<B��J�x9�8�#�D�0?��?�p$!�Z3� T0 k� ��'$2(u e1�t A  ��    � 9��BOhy����8<C�J�x9�8�/�D�8@��A�x%!�Z3� T0 k� ��'$2(u e1�t A  ��    � :��BOpx����8<C�J�|9�8�7�D�@A��B�|&!#�Z3� T0 k� � ~�$~'$2(u e1�t A  ��    � ; BOtx����<<C�I��9�8�?�D�DB.�C��&!+�Z3� T0 k� �,~�0~'$2(u e1�t A  ��    � < BO|x����@<C�I��9�8�G�D�LB.�E��'!3�Z3� T0 k� �4}�8}'$2(u e1�t A  ��    � < BO�x����D<C�I��8�8�O�D�TC.�F��(!7�Z3� T0 k� �@}�D}'$2(u e1�t A  ��    � < BO�w����H<C�I��8�8�W�D�XD.�H��)�?�Z3� T0 k� �L}�P}'$2(u e1�t A  ��    � < BO�w����H<C�I��8�8�_�D�`E.�J��*�G�Z3� T0 k� �T|�X|'$2(u e1�t A  ��    � < BO�w����L<C�I��8�8�k�D�hF.�K��*�K�Z3� T0 k� �`|�d|'$2(u e1�t A  ��    � < BO�w���P<C�I��8�8�s�D�pG.�M��+�S�Z3� T0 k� �h{�l{'$2(u e1�t A  ��    � < BO�v���T<C�I��7�8�{�D�tH�N��,�[�Z3� T0 k� �t{�x{'$2(u e1�t A  ��    � < BO�v���X<C�I��7�8���D�|I�P��-�c�Z3� T0 k� ��z��z'$2(u e1�t A  ��    � < BO�v���\<C�I��7�8���D�J�Q��/�g�Z3� T0 k� ��z��z'$2(u e1�t A  ��    � <  BO�v�'��\<C�I��7�8���D�K�S��0�o�Z3� T0 k� ��y��y'$2(u e1�t A  ��    � < #F�v�/��`<C�I��7�8���D��M�T��1�w�Z3� T0 k� ��y��y'$2(u e1�t A  ��   � < &F�u�7��d<C�I��6�8���D��N�V��2�{�Z3� T0 k� ��x��x'$2(u e1�t A  ��    � < )F�u�?��h<C�I��6�8ͯ�D��O�W��3��Z3� T0 k� ��x��x'$2(u e1�t A  ��    � < ,F�u�G��h<@l�I��6�8ͷ�D��P�Y��5��Z3� T0 k� ��x��x'$2(u e1�t A  ��    � < .F�u�O��l;@l�I��6�8Ϳ�D��Q��Z��6��Z3� T0 k� ��w��w'$2(u e1�t A  ��    � < 0E��uW��p;@l�I��6|8�ǊE��R��\��7��Z3� T0 k� ��w��w'$2(u e1�t A  ��    � < 1E��u_��t;@l�I��5|8�ϊE��S��]��9��Z3� T0 k� ��u��u'$2(u e1�t A  ��     � < 2E��ug��t;@l�J��5|8�׊E��T��^��:��Z3� T0 k� ��t��t'$2(u e1�t A  ��     � < 3E��uw��|:@l�J��5|8��E��V�a�=��Z3� T0 k� ��t��t'$2(u e1�t A  ��     � < 5E��u�܀:@l�J��5|8��E��W�c0?��Z3� T0 k� ��t� t'$2(u e1�t A  ��     � < 7E��t��܄9@l�J��4|8���B��X�d0@��Z3� T0 k� �s�s'$2(u e1�t A  ��     � < 9E��t��܈9@l�J��4 <8��B��Y�e0B��Z3� T0 k� �s�s'$2(u e1�t A  ��     � < ;E� t��܈9@l�K��4 <8��B��Y�g0C��Z3� T0 k� �r�r'$2(u e1�t A  ��     � < =E�t��܌9@l�K��4 <8��B��Z�h0 E��Z3� T0 k� �r� r'$2(u e1�t A  ��     � < ?E�t��܌9@l�K��4 <8��B�[�i0$G��Z3�T0 k� �$r�(r'$2(u e1�t A  ��     � < AE�t߯�ܔ8@l�K��3 <<�'�B�\��j@(I��Z3�T0 k� �,r�0r'$2(u e1�t A  ��     � < CE� t߷�ܘ8@l�K��3 <<�/�B�]��l@,J��Z3�T0 k� �4r�8r'$2(u e1�t A  ��     � < EE�(t߿�ܜ8@l�K��3 <@�7�B�^��m@0L��Z3�T0 k� �<r�@r'$2(u e1�t A  ��     � < GE�0t���ܠ8@l�L��3 <@�?�B�$_��n@8N��Z3�T0 k� �Hn�Ln'$2(u e1�t A  ��     � < IE�8t���ܤ8@l�L��3 <D
�G�B�,_��o@<P��Z3�T0 k� �Pk�Tk'$2(u e1�t A  ��     � < KE�@s�����7@l�L��2 <D	�O�B�4`�p0@Q��Z3�T0 k� �Xh�\h'$2(u e1�t A  ��     � < ME�Hs�����7@l�L��2 <H�W�B�<a�q0DS�Z3�T0 k� �`g�dg'$2(u e1�t A  ��     � < OE�Ts�����7@l�L��2 <L�_�B�Db�s0HU�Z3�T0 k� �lf�pf'$2(u e1�t A  ��     � < Q@p\r�����7@l�L��2 LP�k�B�Lc�t0LW�Z3�T0 k� �xc�|c'$2(u e1�t A  ��     � < S@pdr�����7@l�M��1 LT�s�B�Tc�u0PZ�Z3�T0 k� ��`��`'$2(u e1�t A  ��     � < U@plr�����7@l�M� 1 LX�{�B�\d�v0T^"�Z3�T0 k� ��^��^'$2(u e1�t A  ��     � < W@ptq����7@l�M�1 L\���B�de�w0Xa"#�Z3�T0 k� ��Z��Z'$2(u e1�t A  �     � < YF��p����7@�M�0 Ld ���B�tf��y0Xa"/�Z3�T0 k� ��S��S'$2(u e1�t A ��    � < [F��p����7@�M�0 Lk����B�|g��z0\b"7�Z3�T0 k� ��P��P'$2(u e1�t A ��    � < ]F��p�#���7@�M�0 Ls����B��h��{0dc";�Z3�T0 k� ��L��L'$2(u e1�t A ��    � < ^F��p�+���7@�N�0 Lw����B��h��{0he�C�Z3�T0 k� ��H��H'$2(u e1�t A ��    � < `F��p�3���7@�N�/ L{����B��i��|0lf�K�Z3�T0 k� ��E��E'$2(u e1�t A ��    � < aF��p�;���7B��N� / L�����BΜj��}0pg�O�Z3�T0 k� ��A��A'$2(u e1�t A ��    � < cF��p�?���7B��N�$/ \���ǏBΤj��}0th�W�Z3�T0 k� ��>��>'$2(u e1�t A ��    � < dF��p�G���7B��N�$. \���ϏBάk�~0xj�[�Z3�T0 k� ��:��:'$2(u e1�t A ��    � < fF��p�O���7B��N�(. \���׏Bδl�~0|i�c�Z3�T0 k� ��7��7'$2(u e1�t A ��    � < gF��o�W���7B��N�,. \����Bμl�0�i�g�Z3�T0 k� ��3��3'$2(u e1�t A ��    � < hF��o�_���7B��N�0. \����E��m�0�i�o�Z3�T0 k� ��0��0'$2(u e1�t A ��    � < jF��o�g���7B��N�4- \����E��n�0�h�s�Z3�T0 k� ��,��,'$2(u e1�t A ��    � < kF��o�o���7B��O�8- \�����E��n�$�0�h�{�Z3�T0 k� ��)��)'$2(u e1�t A ��    � < mF��o�w��7B��O�<- \����E��o�(�0�h��Z3�T0 k� ��%��%'$2(u e1�t A ��    � < nF� o���7B��O�@- \����E��o�00�h���Z3�T0 k� ��!��!'$2(u e1�t A ��    � < pF�o����7B��O�D, \����E��p�80�g���Z3�T0 k� ����'$2(u e1�t A ��    � < qF�o����7B��O�H, \����E��p�@0�g���Z3�T0 k� ����'$2(u e1�t A ��    � < sF�o����8B��O�L+ l���'�E� q�D~0�g���Z3�T0 k� ��� '$2(u e1�t A ��    � < tF�o����8B��O�P+ l���/�E�q�L~0�f���Z3�T0 k� � �'$2(u e1�t A ��    � ; uF�$o����8B��O�T+ l���7�E�r�T}0�f���Z3�T0 k� ��'$2(u e1�t A ��    � : wF�,o����$8B��O�X+ l���?�E�r�\}0�f���Z3�T0 k� ��'$2(u e1�t A ��   � 9 xF�4o����(8B��P�X* l���G�E� s�d|0�f���Z3�T0 k� �	�	'$2(u e1�t A ��    � 8 zF�8n����08B��P�\* l���O�E�(s�l{0�e���Z3�T0 k� ��'$2(u e1�t A ��    � 7 {F�@n����48B��P�`* l���[�E�4s�p{0�e·�Z3�T0 k� � �$'$2(u e1�t A ��    � 6 }F�Hn�ǽ�<8B��P�d) l���c�E�4s�|z0�e»�Z3�T0 k� �'��+�'$2(u e1�t A ��    � 5 ~F�Ln�ϼ�D8B��P�h) l���k�E�<s�z0�e¿�Z3� T0 k� �/��3�'$2(u e1�t A ��    � 3 �F�Tn�׻�H8B��P�l) l���s�E�@s�y0�e���Z3� T0 k� �3��7�'$2(u e1�t A ��    � 1 �F�Xn�ߺ�P8B��P�p( l���{�E�Hs��x0�d���Z3� T0 k� �7��;�'$2(u e1�t A ��    � / �F�hn ��\9B� P�t( m�ϋ�B�Xs��w0�d���Z3� T0 k� �C��G�'$2(u e1�t A ��    � - �F�ln ��d9B�P�x( m�ߗ�B�`r��v0�d���Z3��T0 k� �K��O�'$2(u e1�t A ��    � + �F�tn ���l9B�Q�|' m�ߟ�B�hr��v0�d	r��Z3��T0 k� �O��S�'$2(u e1�t A ��    � ) �E�xn��t9B�Q�|' m�ߧ�B�pr��u �d	r��Z3��T0 k� �W��[�'$2(u e1�t A ��    � ' �E��n��|9B�Q��' =#�߯�B�xq��t �d	r��Z3��T0 k� �[��_�'$2(u e1�t A ��    � $ �E��m��݄9B�Q��' ='�߷�E�q��s �e	r��Z3��T0 k� �_��c�'$2(u e1�t A ��    � ! �E��m��݌9E�$Q��& =/����E�q�r �e	r��Z3��T0 k� �g��k�'$2(u e1�t A ��    �  �E��m�#�ݔ9E�,Q��& =3��ǓE�p�q �e	r��Z3��T0 k� �k��o�'$2(u e1�t A ��    �  �E��m�+���9E�0Q��& =;��ϓE�p�p�e	���Z3��T0 k� �s��w�'$2(u e1�t A ��    �  �E��l�7���9E�@Q��% =G���E�op n�f	��Z3��T0 k� �����'$2(u e1�t A ��    �  �E��l�?���9E�DQ͔% =K���E�o m�f	��Z3��T0 k� ������'$2(u e1�t A  ��    �  �E��k�G���9E�LQ͘% =S��E�o l�f	��Z3��T0 k� ������'$2(u e1�t A  ��    �  �E��k�O���9E�TP͜% =W���B��n k�f	r�Z3��T0 k� ������'$2(u e1�t A  -�    �  �E��j�W���:E�\P͜$ =_��B��n $j�f	r�Z3��T0 k� ������'$2(u e1�t A  ��    � 	 �E��j�_���:E�`P͠$ =c��B��n ,i g	r�Z3��T0 k� ������'$2(u e1�t A  ��   �  �E��i�g���:B�hP͠$ Mk��B��n 4hg	r�Z3��T0 k� ������'$2(u e1�t A  ��    �  �E��i�o���:B�pOͤ$ Mo��B��m <gg	r�Z3��T0 k� ������'$2(u e1�t A  ��    �   �E��h�w���:B�xOͨ# Ms�'�B��m�Df�g	��Z3��T0 k� ������'$2(u e1�t A ��    ��� �E��g����:B��Oͨ# M{�/�B��m�Ld�g	��Z3��T0 k� ������'$2(u e1�t A ��    ��� �E��e����:B��N}�# M��?�B�l�`b�$g	��Z��T0 k� ������'$2(u e1�t A ��    ��� �E��e��:B��M}�# M��G�B�l�ha�(g	��Z��T0 k� �ß�ǟ'$2(u e1�t A ��    ��� �E��d��:B��M}�" M��O�B�l�p`�0g	r�Z��T0 k� �Ǜ�˛'$2(u e1�t A ��    ��� �E�c��:B��L}�" M���W�B�$l�x_�4g	r�Z��T0 k� �Ϙ�Ә'$2(u e1�t A ��    ��� �E�a��$:B��K}�" M���_�B�,kЀ^�<g	r�Z��T0 k� �Ӕ�ה'$2(u e1�t A ��    ��� �E�`��,:B��K}�" M���k�B�4kЈ\�@g	r�	Z��T0 k� �ۑ�ߑ'$2(u e1�t A ��    ��� �E�_��4:B��J}�" ]���s�B�<kА[�Hg	r�	Z��T0 k� �ߍ��'$2(u e1�t A ��    ��� �E�^�ˡ�<:C�I}�" ]���{�B�DkМZ�Pf ��	Z��T0 k� ����'$2(u e1�t A ��   ��� �E�$[�۠�L:C�H}�! ]�����B�TjЬW�\f ��
Z��T0 k� ����'$2(u e1�t A  ��    ��� �E�(Z���T;C�G��! ]ä���B�`j�V�de ��
Z��T0 k� ����'$2(u e1�t A  ��    ��� �E�,Y���`;C�G��! ]Ǣ���B�hj�U�he ��bC��T0 k� ��|��|'$2(u e1�t A  (�    ��� �C�0W���h;C�F��  ]ˡ���B�pi��T�pe2�bC��T0 k� 2}�}'$2(u e1�t A  ��    ��� �C�4V���p;C�E��  ]ӟ���B�xi��R�xd2�bC��T0 k� 2~�~'$2(u e1�t A  /�    ��� �C�<S�΀;C D�� ]ߜp��B��ip�Pфc2�bC��T0 k� 2�'$2(u e1�t A  ��    ��� �C�@R�Έ;CC� ]�pǘB��ip�Nьc2�bC��T0 k� 2���'$2(u e1�t A  ��    ��� �C�DP�ΐ;CB� m�pϘB��hp�Mєb"�bC��T0 k� ����'$2(u e1�t A  ��    ��� �C�DO'�Θ;CA� m�pחB��hp�Kќa"�bC��T0 k� �#��'�'$2(u e1�t A  ��    ��� �C�HL7�Ψ;C(?� m��@�B��hq H�`"�bC��T0 k� �+��/�'$2(u e1�t A  ��    ��� �C�LJC�ް;C,?�� n�@�B��h�F�_"�bC��T0 k� �3��7�'$2(u e1�t A  ��    ��� �C�LHK�޸;C4>�� n�@��B��g�E�^�Z��T0 k� �7��;�'$2(u e1�t A  ��    ��� �C�PGS���;C<=�� n�A�B��g�C��]�Z��T0 k� �?��C�'$2(u e1�t A  ��    ��� �C�PE[���;CD<�� n�A�B��g�A��] Z��T0 k� �C��G�'$2(u e1�t A  ��    ��� �C�TBo���;CT:�� n���B��g�,>��[ Z��T0 k� �O��S�'$2(u e1�t A  ��    ��� �C�T@w���;C\9�� n#��#�B��f�0<��ZZ��T0 k� �S��W�'$2(u e1�t A  ��    ��� �C�T>���;Cd8�� n+��+�B��f�8:��XZ��T0 k� �W��[�'$2(u e1�t A  ��    ��� �C�T<����;C.l7��~+��/�B� f�@9��VZ��T0 k� �_��c�'$2(u e1�t A  ��    ��� �C�T:����;C.p7��~+��7�B�f�D7�T�Z��T0 k� �c��g�'$2(u e1�t A  ��    ��� �C�T9��� <C.x6��~+�?�B�f�L5�R�Z��T0 k� �g��k�'$2(u e1�t A  ��    ��� �C�T7���<C.�5� ~+�G�B�f�P3�P�Z��T0 k� �o��s�'$2(u e1�t A  ��    ��� �C�T5���<C.�4�~+�O�B�$e�X1�(N�bS��T0 k� �s��w�'$2(u e1�t A  ��    ��� �C�T3���<C.�3�~+�W�B�,e�\/�4L�bS��T0 k� �w��{�'$2(u e1�t A  ��    ��� �C�T/�ã�(<C.�1�~+�c�B�<e�h+�HI�bS��T0 k� ������'$2(u e1�t A  ��    ��� �C�P-�ˣ�4<C.�0��+�k�B�De�p*�TGsbS��T0 k� ������'$2(u e1�t A  ��    ��� �C�P+�ף�<<C.�/��+�s�B�Le�t(�`Es bS��T0 k� ������'$2(u e1�t A  ��    ��� �C�P)�ߣ�D<C.�.� �+��w�B�Te�|&�hCs$bS��T0 k� ������'$2(u e1�t A  ��    ��� �C�L'���L<B��-�$
�+���B�`d��$�tBs$bS��T0 k� ������'$2(u e1�t A  ��    ��� �C�L%���T<B��,�(	�+��B�hd��"�|@s(bS��T0 k� ������'$2(u e1�t A  ��    ��� �C�H#����\<B��+�,�+��B�pd�� >�(bS��T0 k� ������'$2(u e1�t A  ��    ��� �C�H!���d<B��*�0�+��B�xd��=�,bS��T0 k� ������'$2(u e1�t A  ��    ��� �C�D���t<B��(�<�+����B��d��¤9�0Z��T0 k� ������'$2(u e1�t A  ��    ��� �C�@���|<E�'�@�+����B��d��°8�4Z��T0 k� ������'$2(u e1�t A  ��    ��� �C�<�#���<E�&�D�+����B��c��¸6�8Z��T0 k� ����Ú'$2(u e1�t A  ��    ��� �C�<s+���<E�%�L �+����B��c����5�8Z��T0 k� �Û�Ǜ'$2(u e1�t A  ��    ��� �                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��_R ]�0�0� � �����3  Y Y     � �ˋ    ���� ��[    �6            %	 ��             �@�     ���  		'           ����   � �
	   � ��    ���. ���    ���   
        #  	��          
 �    ���  @
	"           1�   � $      �c     1\o �\     �             k��          �p�     ���  8
(         ��\�  � �	    ��    �� #��    �                 [	��           @�  !  ���   8
          ����   � �
	   .��    ������    �[<               #��           +@�  #  ���  X
	         �}S�  M M       B ��f    �|ș �k6    ��             	 �� �}         �     ���  0	
          ��W         V �C^    ��@� ��x    N�               	     !�        0     ��B   0

 
 
          H�       j ��     H�W ��]    ����              & 
	 S �               ��B@ (
 
          ���D        ~ Ș&    ���# ȉF    � �                �         P     ��@   8�         ���#        ���    ���#��                            �         	       ��@   (
           ����         � �Nh    ���� �:Z    .               �         
 ��      ��@   @



	A

         ��V��       � �5    ��V �5                              �� �                ��H    8		 1                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          %�   ��        ���  *� "���  *� �                x                j  �       �                          %    ��        �       "             "                                                �                          � �  � � � � � ���   	       
       
  �   � �� �L�E       B� �[� �$ f� �D f� �d g  Є g  Ф g@ A d� A$ d� Ф ]@���X ���� ����  ����. ����< ����J ����X � 
�� V� 
�\ W  � s` 
�\ W  
� W� 
�< W� 
�\ W� � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }`���� � �� �c@ �� d@ � d` �$  d� �d d� �� d� �� @`� �$ a@ �D  a` �� a� �� 0a� �  b  �D b` ބ �^@ Τ w@ �� `w` τ x  ��  }` �� }����� � )D  n  
�\ U� 
�� V  
�| V  
�\ V� 
�� V� 
�\ W  
�\ W� 
�� W� 
�| W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����   �����   ������  
�fD
��L���"����D" � j  "  B   J jF�"     "�j  " ��
��
��"    B�j l �  B �
� �  �  
�  1    ��     �        1    ��     �       ��   ��     � �          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �"(( 1      �� � �  ���        �tS  ���        �        ��        �        ��        �    ��     , P�C��        ��                          �w� $  ����                                     �                ���             1 ���%��  ��  2                22 Christan Ruuttu     1:34                                                                        2  2      �Tkj|lkrlKB �# KJ �c~ �( c� � �J� � �c� �	c� � �
cV � c^ � � k�" �k� c^ � � k�" �k� �B� � � B� � � B� � � B� � � B� � � B� � �Cd � C\ �c� � c� � �[ � �Z �K � �K � �K � �  K" � �!K# � �	"�$ �	#�; �$�" �%�M �&C. � � 'C6 � � (C7 � � )C8 � � *C9 � � +C: � �,"�a � -"�s �.�] �/
�l �0"�a � 1"�s �2"�] �3*�l4"� 5"�' �6� �7
� �8"( � � 9"O � �:"( � � ;"O � �<" � � =!� � � >"Q � � "6 �                                                                                                                                                                                                                         �� R         � $   @        �     [ P E `  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    ���   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, 6� * (�� L� t�@~@�@�� �                                                                                                                                                                                                                                                                                                                                �� �"�.�����                                                                                                                                                                                                                                 a    ,    � �  4�J �    -�                             �������������������������������������������������������                                                                                                                                   |  �� r            �          ��               	 
     ���������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ����           y                            ��  L�J      9  	                           ������������������������������������������������������                                                                                                                                        $   7�� (            �         �� �               	 	 � ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� ������������������            ?                                                                                                                                                                                                                                                 
                                        	                    �             


            �   }�                                                                '�  'w                     ������������  R�  'q����������������������������  R���������������������     'q������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" A C 6                                 � -'�� �\                                                                                                                                                                                                                                                                                       )n)n
  �        a            m                m            `                                                                                                                                                                                                                                                                                                                                                                                                        > �  >�  @�  (�  (�  EZm2 ���y��� � �N ���d�{�����X�����������������2                 y � :�r��	          �   &  AG� �   �                    �                                                                                                                                                                                                                                                                                                                                        N I   �                     !��                                                                                                                                                                                                                            Y��   �� � ���      �� 8      ���������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ����� ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ;      .   �                         8     �   �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$     `d  �@���6 ��  �@���6 �$ ^$ �y@  �@  �y@   � 
�" ��       j���� ��  j���� �$ ^$    j  ��             � ��� ��  e� � ��� �� � ��� Y! �  ��  �      �       "�����������J g���   �     f ^�         ��  ��      "      ��_��������J���J��u����      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                          �      �  a r!   f�"""""*��**"*�"�""�""v""*f   "  ""- ��"�"*"-""z"""""����            n   �  "  q  ��                          �  �                                 � gv"!g�vg�vggfvv|�b��r""gb"�vr�rgb��v���g���v���***�*q!q�"!a�!vwfqqr~� qw��q�~~q�����~~~�w~~w�w            �   ~   ��  ~~  �w      v    �                ggj�vvggvvgg!vg�g֪vvg�r�r��⢪rq**gjb�v�q*gjj*vv��gg�z�/�"!�"�*�""*z����qw�~q~ww��q~qwvq�w�`� ��� �w �~p w�p  ��                    �                        lggz�v��g        �       ggbvvrgggavvvqggav� �      ���w!z�w"""�!""*�"! ��        q� q�        `               �        �                      wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         7v` weV "fff"O�p"��p"��p"�p3�}p-��p=��p|� }�  }�  ��  ��  ��  ��  �  �  �  �  �  "              `  eV  fff O�  ��  ��  �  �} �� �� ��  |�  }�  ��    =   }   =   =              �������}�}�}�ww~r�� ∈�������������������}�� }�� ��� ��� ����   �   �   �   �   �   �   �   C""42""#2""#2""#2""#s3342"""3333    p   p   p   p   p   p   p    ��������� ��� }�� ��  ��  ����  ��  ��  ��  ��  ��  ��  ��                          � �� ��    "               wvf wfU 7Of`w��f"�� "�p-�}p���� ��� ����x��	�� �� �� "�        f  U` f` f` �p w���� `  eV  ff  O�  ��  �� ����}�                �  �  ��  �            �  �  �   �  ��  �                     �  �  �   � `  eV  ff  O�  ��  ��  ����}���������������p	���         `  eV  ff  O�  ��  ��  ���}�     �  �  �   �  ��  �   �            ��  ��  �   ��  �   ���������������p	���                    3333UUUU                        wwww                    333333333333333333333   w  G� ws@ ws� ws$7w@wwww"                               ����������� ��� �� ��  �    `  eV  ff  O�  ��  ��  � ��}�            """"                 �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                                                �����   �   �   �   ����                                     
�  

  
 � 
 
 
   
   
   
   
  ��                  ��   
   
   
   
   
   
 
 
 � 

  
�                 �   
    �   
    �   
    �   
   
   �  
   �  
   �  
   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    "!  "" "  """ "! ""! " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ "! ""! " ""  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  " ! " ""                "                                                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                       �� wڪ z�� ���
���	������
���̪��̹����ӈ��E �U ��U�UD�D 
��  ��  ˰ ",� """��"" ��  �    �   �   ��  ̨  ̋  �۰ �۰ ��� �=  30  DC  UD0 T4J 3DT�4U@ 3D� ;�  �   �   ��  ��  �   �   �   ""  �"  � ��� �                      ̰ ̻ ��                               �   �   ��  � " ��"  "                     �                             ���                         �  ��                    �����                         �     �                                       �   ���                            �   �                                                                                                         �  �  �  �� ݚ� }�Ȫ��˙������˼� ��  ��  ��  ��  ��  I� H� �E X�T X�S T�D �[ ˻  ˸  ��  
� �,"��"" "  �" �  ""� �� ˻ �˻ ��ݪ��کɨ��ˀ�̽ ��� ��  ̽  ̻  ̻  ˉ  ��  �D  DC  C3  #;  ;�� �� ��  �� "�  "  �"/ / ����� ��  �      �   �          �  �  "     "  "  "   "�  �  �   �   
                            �          �   �          �                    ��  ���� ��    �����                                                                                                                                                                                                                           �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �          
 "� ""� ""� "                       �                             ���                         �  ��                    �����                                                                                                                                                                                                                      ۻ� ۽� ��� H�DH�D�DP�E X�T H�P H�@ Ȥ� ̻� ˘ �� "*� �/�""/""/���                       ��  ۼ� ݻ� w�� b}ذgvz�w������ɨ�ͨ���ڋ��٭���ۻݻ� �   �          �   �   .   ."  ""  ""  ,   �   
            "  "  ""  "�   �           �   ��  �      �                                     �  �  �  ��  �  �  �  ��  �             �   �   �             � � "            � "�",�"+� ",                       "  .���"    �     �                                                                                                                                                                                          �  �  �  �� ݚ� }�Ȫ��˙������˼� ��  ��  ��  ��  ��  I� H� �E X�T X�S T�D �[ ˻  ˸  ��  
� �,"��"" "  �" �  ""� �� ˻ �˻ ��ݪ��کɨ��ˀ�̽ ��� ��  ̽  ̻  ̻  ˉ  ��  �D  DC  C3  #;  ;�� �� ��  �� "�  "  �"/ / ����� ��  �      �   �          �  �  "     "  "  "   "�  �  �   �   
                            �          �   �          �                    ��  ���� ��    �����                       ��                                 � ���� ��   � � �                                                                                                                                    ˰ ̻ ̻ �� {�  �� 
�� ��� ��� ������
���	��ܻ̍ݻ���"� 8"  8  �  D�  H�  X�  ��  �   �          "  "     �                        ��  ��� �̺�̻����ۻ�˽��̽��̝ ̙� �30 �EP �U@ �T0 EC0 T3  C:  K�  �"  �"/ ����˽� �"� "" �""� � �� ��      �   �� ��  �"  �            �   �"  ""  !� �� ��  �               �   ������  ��           �   �    �   �       �   �   �                .                                                                                                                                                                                                                                   �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                      �  �� ��  �    � ���                                                                                                                                                                                                           �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �      �   �                                �   �       �    �                     �   �  �  �                    ��  ��  ���       +  "  "     �  �                                                                                                                                                                                   �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                 �� �̽���ݪ۽w�}�֪�vv���p��� �  �� 	  
  �  ",  ""  �"   "                      ��  ��  �          ���� ��� ����         �EU �E  
�   �               �"�!/"�  �                       � ���� ��   � � �                                                                                                                                  �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �   �   "   "   "  !�    ��                                 �   �                      �������  ���    �                                                                                                                                                                                                                                               �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �        �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��  ��  ��� ���                                  � �������������               �  �     �   �  �  �                                                                                                                      �� �����ݼڜ��ک��ک��z�	��� 
�� 
�� 	�� ̘ ɪ  ��  �  �� �� ������������ ���  � � � �� �� ������ ��                      �   ��  ��  �̰ ��� ��˰�̻��̻���������ˉ�U��EP�ET �I� ٕ  �D� �L� ��� ��" ����/�"�"�""�����                         ��  ��� ��  �                                        �� ��           �   �                   �  ��  ��  ��  ��� ��� ��� ��˰ɜ˰��˻�̻���������3���DDD�                                                                                                                                                                                                             �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��           	 
          
        ((((((( 
	(((( ����������������             ! " # $ % & '   ( $ % ) ! " # * ('(&(%($(#("(! (((���������������� + , -   . / 0 1  	 2         3       4 (((((((2	10/(.(-(,(+���������������� 5 6   7   8 9 1 :   $ % ) ! " #   ; ) ! " # $ % ) (#("(!()(%($ :198(((7(6(5����������������    <     = 8 0 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>108(=((( (<���������������� L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L����������������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7����������������  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(�����������������333333333333333333333333333333333333333333333333333333333333����  
�fD
��L���"��������������������D" � j  "  B   J jF� ����
��� �����
���� ����
��� �����
��� 0 q����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqTkj|lkrlKB �$ KJ �c~ �( c� � �J� � J� � � 	J� �
J� � �c� �c� � �cV � c^ � � k�" �k� �B� � � B� � � B� � � B� � � B� � � B� � �Cd � C\ �c� � c� � �[ � �Z �K � �K � �K � �  K" � �!K# � �	"�$ �	#�; �$�" �%�M �&C. � � 'C6 � � (C7 � � )C8 � � *C9 � � +C: � �,"�a � -"�s �.�] �/
�l �0"�a � 1"�s �2"�] �3*�l4"� 5"�' �6� �7
� �8"( � � 9"O � �:"( � � ;"O � �<" � � =!� � � >"Q � � "6 �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3�����������������������������������������#��<�Z�K�\�K��6�G�X�S�K�X� � � � � � � � �-�2�3�������������������������������������������-�N�X�O�Y�Z�G�T��;�[�[�Z�Z�[� � � � � �-�2�3�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�2�3� �� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������,�-��.�/�0�1�2������������������������� �!�"�3�4�#�#�#�#�#�#�#�#�$������������������%�&�'�(�)�)�)�)�)�)�)�)�)�)�*�+������������������5�6���7�8�9�:�;�<�=�>�?�������������������� �!�"�#�#�#�#�#�#�#�@�4�#�$������������������%�A�B�C�D�E�F�G�H�I�J�K�L�M�N�O�����������������P�Q�R�S�T�U�V�W�X�Y�W�Z�[�\�]�^�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 