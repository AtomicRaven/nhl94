GST@�                                                            \     �                                               9 ��       �  d   6         ����e J���J�������������������        Fi     	#    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    
 �j
  ����
��
�"     "�j��   * ��
  �                                                                               ����������������������������������      ��    bb? QQ0 5 118 44               		 


     
               ��� 4    �                 nnY ))         88:�����������������������������������������������������������������������������������������������������������������������������=  0b  4  11                                         �  �  �  �                  F  
1          = �����������������������������������������������������������������������������                                ��  �       ��   @  #   �   �                                                                                '      )n)nY  
1F    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    �|E�7�C�8*1?����l;��s�|0Da��Ic��A��3��T0 k� �w��{���1"t'!(e1't   ��:    ��� $�|E�;�C�0*�?����l;��k�x1Da��Ic��A��3��T0 k� �o��s���1"t'!(e1't   ��:    ��� #�{E�?�C�()�;����l;��c�p1Da� @���1��3��T0 k� �k��o���1"t'!(e1't   ��:    ��� "�{E�?�C� (�7����l;��[�h1Da�@���1��3��T0 k� �g��k���1"t'!(e1't   ��:    ��� !�zErG�C�'�7����l;��G�X2I�x@���1��3��T0 k� �[��_���1"t'!(e1't   ��:    ���  �zErK�C�&�3� ��l;��?��P2I�p@���1{�3��T0 k� �W��[���1"t'!(e1't   ��:    ��� �yErK�C� %�+� ��l;��7��H2I�h@���Aw�3��T0 k� �S��W���1"t'!(e1't   ��:    ��� �yErO�C��$�'� ��l;��/��@3I�dA��As�3��T0 k� �K��O���1"t'!(e1't   ��:    ��� �yErS�C��$�� ��l;��'��83I�\A��Ao�3��T0 k� �G��K���1"t'!(e1't   ��:    ��� �xxErW�C��#�� ��l;����03I�TA��Ak�3��T0 k� �C��G���1"t'!(e1't   ��:    ��� �lxEr[�C��!�� ��l;���� 4I�H	A��Q_�3��T0 k� �;��?���1"t'!(e1't   ��:    ��� �dwEr_�C�� �� ��l;����4I�D	A��Q[�3��T0 k� �7��;���1"t'!(e1't   ��:    ��� �\wEr_�C����� ��l;�����4I�<
A��QW�3��T0 k� �/��3���1"t'!(e1't   ��:    ��� �TwErc�C����� ��l;�	���5EQ8A��QS�3��T0 k� �+��/���1"t'!(e1't   ��:    ��� �LvEbg�C����� ��l;�	��� 5EQ4A��QO�3��T0 k� �'��+���1"t'!(e1't   ��:    ��� �HvEbg�C�������l;�	����5EQ,A��aK�3��T0 k� �#��'���1"t'!(e1't   ��:    ��� �8vEbk�C������l;�	�׳��6EQ A��aC�3��T0 k� ������1"t'!(e1't   ��:    ��� �0uEbk�C�����{�l;�	�ϳ��6EQAS��a?�3��T0 k� ������1"t'!(e1't   �:    ��� 	(uEbo�C�����s�l;�	�ǳ��6EQAS��a;�3��T0 k� ���󭑕1"t'!(e1't  ��?    ����� uEbo�C��P��k�l;�	�ó��6EQAS��q7�3��T0 k� �׭�ۭ��1"t'!(e1't  ��?    �����tEbo�C��P��c�l;�	�����6EQAS��q3�3��T0 k� ��í��1"t'!(e1't  ��?    �����tEbo�C��P��[�l;�	�����7EP�AS��q/�3��T0 k� ������1"t'!(e1't  ��?    �����tEbs�C�xP��S�l;�᯳м7C��AS��q+�3��T0 k� ��������1"t'!(e1't  ��?    ������sEbs�C�pP��K�l;�᧳д7C��AS��q'�3��T0 k� �{�����1"t'!(e1't  ��?    ������sERs�C�lP��C�l;�ᣳЬ7C��AS���#�3��T0 k� �c��g���1"t'!(e1't  ��?    ������sERs�C�dP���;�l;�ᛳФ8C��AS����3��T0 k� �K��O���1"t'!(e1't  ��?    ������sERs�C�\P���3�l;�ᓳМ8C��AS����3��T0 k� �3��7���1"t'!(e1't  ��?    ������rERo�C�TP���/�l;�ᏳД8EP�AS����3��T0 k� ������1"t'!(e1't  ��?    ������rERo�C�LP���'�l;�ᇳЌ8EP�AS����3��T0 k� ������1"t'!(e1't  ��?    ������rERo�C�HP����l;�����8EP�AS����3��T0 k� ���󬑕1"t'!(e1't  ��?    ������rERk�C�@P����l;��w��|9EP�AS����3��T0 k� �׬�۬��1"t'!(e1't 	 ��?    ������qERk�C�8P����l;��o��t9EP�AS����3��T0 k� ����ì��1"t'!(e1't 	 ��?    ������qERg�C�0P����;��g��l9EP�AS����3��T0 k� ��������1"t'!(e1't 
 ��?    ������qC�g�C�(P{�����;��_��d9EP�AS����3��T0 k� ��������1"t'!(e1't 
 ��?    ������qC�c�C�$
Pw�����;��[��\9E@�AS����3��T0 k� �{�����1"t'!(e1't  ��?    ����~�qC�c�C�	Po�����;��S��T9E@�AS�����3��T0 k� �c��g���1"t'!(e1't  ��?    ����y�pC�_�C�Pk�����;��K��L8E@|AS�����3��T0 k� �K��O���1"t'!(e1't  ��?    ����t�pC�[�C�Pg�����;��C��D8E@tAS�����3��T0 k� �7��;���1"t'!(e1't  ��?    ����p|pC�W�C�Pc�����;��7��<8E@lAS�����3��T0 k� ���#���1"t'!(e1't  ��?    ����ltpC�S�C� P[�����;��/�048E@`AS����3��T0 k� ������1"t'!(e1't  ��?    ����h�hoC�O�C��PW�����7��'�0,8E@XAS����3��T0 k� ���󫑕1"t'!(e1't  ��?    ����e�`oC�K�E��PS�����7���0$8E@PAS����3��T0 k� �۫�߫��1"t'!(e1't  ��?    ����b�XoC�G�E��PO����|7���07E@DAS����3��T0 k� �ë�ǫ��1"t'!(e1't  ��?    ����_�PoC�C�E�� PK����|7���07E@<AS����3��T0 k� ��������1"t'!(e1't  ��?    ����\�HoC�?�E���PG����|7���07C�4AS�� �3��T0 k� ��������1"t'!(e1't  ��?    ����Y�<nC�;�E���PC����|7� ��06C�(AS�� �3��T0 k� �{�����1"t'!(e1't  ��?    ����V�4nC�7�E���P?����|7� �0 6C� AS�� �3��T0 k� �g��k���1"t'!(e1't  ��? 	   ����T�,nC�/�E���P;�����7� �?�6C�AS�� ߕ3��T0 k� �O��S���1"t'!(e1't  ��? 	   ����R�$nC�+�E߿�P7����7� �?�5C�AS�� ە3��T0 k� �7��;���1"t'!(e1't  ��? 	   ����P�nC�'�E߷�P3����7� ۳?�5E�AS�� ە3��T0 k� ���#���1"t'!(e1't  �? 	   ����P�nC��EO��P/���7�Pӳ��5E��AS�� ו3��T0 k� ������1"t'!(e1't  �? 	   ����P�mC��EO��P+�w��7�Pǳ��4E��AS�� Ӕ3��T0 k� �������1"t'!(e1't  ��? 	   ����P� mC��EO��P'�o��7�P����4E��AS�� Ӕ3��T0 k� �۪�ߪ��1"t'!(e1't  ��? 	   ����P��mC��EO��P#��g��7�P����4E��AS�� ϔ3��T0 k� �ê�Ǫ��1"t'!(e1't  ��? 	   ����P��mC��EO��P��_��7�P����3E��AS�� ϔ3��T0 k� ��������1"t'!(e1't  ��? 	   ����P��lC���EO��P��[��7�P����3E��AS�� ˓3��T0 k� ��������1"t'!(e1't  ��? 	   ����P��lD��EO��P��O��7�P����2E��AS�� ˓3��T0 k� �������1"t'!(e1't  ��? 	   ����P��lD��EO��P��G��7�P����2E߼AS�� Ǔ3��T0 k� �g��k���1"t'!(e1't  ��? 	   ����P��kD��EO{�P��?��7�P����2A_�AS�� Ǔ3��T0 k� �O��S���1"t'!(e1't  ��? 	   ����P��kD��EOw�P��7��7�P����1A_�AS�� Ó3��T0 k� �7��;���1"t'!(e1't  ��? 	   ����P0�jD��C�o�P��/��7�P����1A_�AS�� Ò3��T0 k� �#��'���1"t'!(e1't  ��? 	   ����P0�jD��C�g�P��'��7�P{���1A_�AS�� ��3��T0 k� ������1"t'!(e1't  ��?	   ����P0�jD��C�c�P����7�Ps���1A_�AS�� ��3��T0 k� �������1"t'!(e1't  ��? 	   ����P0�iD��C�[�_�����7�Pk���0A_�AS�� ��3��T0 k� �۩�ߩ��1"t'!(e1't 
 ��? 	   ����P0�iD��C�S�_��?��7�Pg���0A_�AS�� ��3��T0 k� �é�ǩ��1"t'!(e1't 
 ��? 	   ����P0�hD��C�O�_��?��7�P_��|0A_�AS�� ��3��T0 k� ��������1"t'!(e1't 
 ��? 	   ����P0�gD��C�O�_��?��7�PW��t/A_xAS�� ��3��T0 k� ��������1"t'!(e1't 	 ��? 	   ����P0�gD��C�G�_��>���7�PS��p/A_pAS�� ��3��T0 k� �������1"t'!(e1't 	 ��?    ����P0xfD��C�?�_��>���7�PK��l/A_hAS�� ��3��T0 k� �g��k���1"t'!(e1't  ��?    ����P0pfD��C�;�_��>���7�PC��d.A_dAS�� ��3��T0 k� �S��W���1"t'!(e1't  ��?    ����P0heD��C�3�_��>���7�P?��`.A_\AS�� ��3��T0 k� �;��?���1"t'!(e1't  ��?    ����P0`dD��C�+�_��>���7�P7��X.A_TAS�� ��3��T0 k� �#��'���1"t'!(e1't  ��?    ����P@XdD{�C�#�_��N���7�P3��T.A_PAS�� ��3��T0 k� ������1"t'!(e1't  ��?    ����P@LcDo�C��_��N���7�P+��P-A_HAS�� ��3��T0 k� �������1"t'!(e1't  ��?    ����P@DbDg�C��_��N���7�P'��H-A_DAS�� ��3��T0 k� �ߨ�㨑�1"t'!(e1't  ��?    ����P@<bD_�C��_��N���7�P��D-A_<AS�� ��3��T0 k� �Ǩ�˨��1"t'!(e1't  ��?    ����P@4aDW�C��_��N���7�P��@-A_4AS�� ��3��T0 k� ��������1"t'!(e1't  ��?   ����P@,`DO�C��_��N���7�P��<,A_0AS�� ��3��T0 k� ��������1"t'!(e1't  ��?    ����P@$_C�C�C���_��N���7�P��8,A_(AS�� ��3��T0 k� ��������1"t'!(e1't  ��?    ����P@_C�;�C���_��N���7�P��0,A_$AS�� ��3��T0 k� �k��o���1"t'!(e1't  (�?    ����P@^C�3�C���_��N���7�P��,,A_ AS�� ��3��T0 k� +k��o���1"t'!(e1't  ��?    ����P@]C�+�C���_��N���7�_���(+A_AS�� ��"s� T0 k� +o��s���1"t'!(e1't   ��?    ����P@\C�#�C���_��N���7�_���$+A_AS�� ��"s� T0 k� +s��w���1"t'!(e1't   ��?    ����P_�[C��C���_��^���7�_�� +A_AS�� ��"s� T0 k� +w��{���1"t'!(e1't   ��?    ����P_�[C��C���_��^{��7�_��+A_AS�� ��"s� T0 k� +{�����1"t'!(e1't   /�?    ����P_�ZC��C���_��^s��7�_��+A_AS�� ��"s� T0 k� +{�����1"t'!(e1't   ��?    ����P_�YC���C���_��^k��7�_��*A^�AS�� ��"s� T0 k� �������1"t'!(e1't   ��?    ����P_�XC���C���_��^g��7�_߳�*A^�AS�� ��"s� T0 k� ��������1"t'!(e1't   ��?    ����P_�WC���E޳�_��^_��7�_۳�*A^�AS�� ��"s� T0 k� ��������1"t'!(e1't   ��?    ����P_�VC���Eޯ�_��^W��7�_׳�*A^�AS�� ��"s� T0 k� ��������1"t'!(e1't   ��?    ����P_�UC���Eާ�_��^O��7�_ӳ� *A^�AS�� ��"s� T0 k� ��������1"t'!(e1't   ��?    ����P_�TC���Eޟ�_��^G��7�_ϳ��)A^�AS�� ��"s�T0 k� ��������1"t'!(e1't   ��?    ����P_�TC���Eޗ�_��^C��7�_˳��)A^�AS�� ��3�T0 k� ������1"t'!(e1't   ��?    ����P_�SC��Eޏ�_��^;��7�_ǳ��)A^�AS�� ��3�T0 k� �����đ�1"t'!(e1't   ��?    ����Po�RC��Eދ�_��n3��7�_����)A^�AS�� ��3�T0 k� �����Ƒ�1"t'!(e1't   ��?    ����Po�QC��Eރ�_��n+��7�_����)A^�AS�� ��3�T0 k� �����ȑ�1"t'!(e1't   ��?    ����Po�PC��C�{�_��n#��7�_����(A^�AS�� ��3�T0 k� �����ʑ�1"t'!(e1't   ��?    ����Po�OC��C�s�_��n��7�_����(A^�AS�� ��3�T0 k� �����̑�1"t'!(e1't   ��?   ����Po�NC��C�k�_��n��7�_����(A^�AS�� ��3�T0 k� �����Α�1"t'!(e1't   ��?    ����Po|MC���C�c�_��>��7�_����(A^�AS�� ��3�T0 k� �����Б�1"t'!(e1't   ��?    ����PotLC��C�_�_��>��7�_����(A^�AS�� ��3�T0 k� �����ґ�1"t'!(e1't   ��?    ����PolKD w�LW�_��>��7�_����(A^�AS�� ��3�T0 k� �����ԑ�1"t'!(e1't   ��?    ����PohJD o�LO�_��=���7�_����'A^�AS�� ��3�T0 k� �����֑�1"t'!(e1't   ��?    ����Po`ID c�LG�_��=���7�_����'A^�AS�� ��"��T0 k� �����ؑ�1"t'!(e1't   ��?    ����PoXHD [�LC�_��=���7�_����'A^�AS�� �"��T0 k� �����ڑ�1"t'!(e1't   ��?    ����P?PFD S�L;�_��=���7�_����'A^�AS�� �"��T0 k� �����ܑ�1"t'!(e1't   ��?    ����P?HED G�L3�_��=���7�_����'A^�AS�� �"��T0 k� �����ޑ�1"t'!(e1't   ��?    ����P?@DD ?�L/�_��=���7�_����'A^�AS�� �"��T0 k� ��������1"t'!(e1't   ��?    ����P?8CD 7�L'�_��=���7�_����'A^�AS�� �"��T0 k� �����⑕1"t'!(e1't   ��?    ����P?0BD /�L#�_��=���7�_����&A^�AS�� {�"��T0 k� �����䑕1"t'!(e1't   ��?    ����P?(AEP#�L�_��=���7�_����&A^�AS�� {�"��T0 k� �����摕1"t'!(e1't   ��?    ����P? @EP�L�_��M���7�_����&A^�AS�� {�"��T0 k� �����葕1"t'!(e1't   ��?    ����P??EP�L�_��M���7�_���&A^�AS�� {�"��T0 k� �����ꑕ1"t'!(e1't   ��?    ����P?>EP�L.�_��M���7�_{���&A^�AS�� w�"��T0 k� �����ꑕ1"t'!(e1't   *�?    ����P?=E_��L.�_��M���7�_w���&A^�AS�� w�3�T0 k� +����ꑕ1"t'!(e1't   /�?    ����P?;E_��L-��_��M���7�_s���&A^�AS�� w�3�T0 k� +����鑕1"t'!(e1't   ��?   ����P>�:E_��L-��_��M���7�_s���%A^�AS�� w�3�T0 k� +����鑕1"t'!(e1't   ��?    ����PN�9E_� L-�_��M���7�_o���%A^|AS�� w�3�T0 k� +����葕1"t'!(e1't   ��?    ����PN�8E_� L-�_��M���7�_k���%A^|AS�� s�3�T0 k� +����葕1"t'!(e1't   ��?    ����PN�7E_� L-�_��M���7�_g���%A^xAS�� s�3�T0 k� �����瑕1"t'!(e1't   ��?    ����PN�6EO�L-�_��M���7�_g���%A^tAS�� s�3�T0 k� �����瑕1"t'!(e1't   ��?    ����PN�4EO�L-߹_��M���7�_c���%A^pAS�� s�3�T0 k� �����摕1"t'!(e1't   ��?    ����PN�3EO�L-۸_�M���7�__���%A^pAS�� s�3�T0 k� �����摕1"t'!(e1't   ��?    ����PN�2EO�L-ӷ_{�M���7�__���%A^lAS�� o�3�T0 k� �����呕1"t'!(e1't   ��?    ����PN�2EO�L-Ϸ_w�M���7�_[���$A^hAS�� o�3�T0 k� �����呕1"t'!(e1't   ��?    ����PN�1EO�L-˶_s�M���7�_W���#A^dAS�� o�3�T0 k� �����䑕1"t'!(e1't   ��?    ����PN�1EO�L-Ƕ_o�M��7�_W���#A^dAS�� o�3�T0 k� �����䑕1"t'!(e1't   ��?    ����PN�0EO�L-õ_k�M{��7�_S���"A^`AS�� o�3�T0 k� �����㑕1"t'!(e1't   ��?    ����P^�0EO�L-��_g�Ms��7�_O���!A^\AS�� o�3�T0 k� �����㑕1"t'!(e1't   ��?    ����P^�/K��L-��_c�Mo��7�_O���!A^\AS�� k�3�T0 k� �����⑕1"t'!(e1't   ��?    ����P^�.K��L-��__�Mk��7�_K��� A^XAS�� k�3�T0 k� �����⑕1"t'!(e1't   ��?    ����P^�.K��L-��_[�Mg��7�_K��| A^TAS�� k�3�T0 k� ����ᑕ1"t'!(e1't   ��?    ����P^�.K��L-��_W�Mc��7�_G��xA^TAS�� k�3�T0 k� ����ᑕ1"t'!(e1't   ��?    ����P^�-K��L-��_S�M_��7�_C��tA^PAS�� k�3�T0 k� ���ᑕ1"t'!(e1't   ��?    ����P^�-K��L-��_O�M[��7�_C��pA^LAS�� k�3�T0 k� ������1"t'!(e1't   ��?    ����P^�,K��L-��_K�MW��7�_?��lA^LAS�� g�3�T0 k� ������1"t'!(e1't   ��?    ����P>�,K��L-��_G�MW��7�_?��lA^HAS�� g�3�T0 k� ���ߑ�1"t'!(e1't   ��?    ����P>�,K��L-��_C�MS��7�_;��lA^DAS�� g�3�T0 k� ���ߑ�1"t'!(e1't   ��?    ����P>�,K�|L-��C�MO��7�_;��hA^DAS�� g�3�T0 k� ���ޑ�1"t'!(e1't   ��?    ����P>�+K�xL-��?�MK��7�_7��dA^@AS�� g�3�T0 k� ���ޑ�1"t'!(e1't   ��?    ����P>�+K�tL-��;�MG��7�_7��`A^<AS�� g�3�T0 k� ���ݑ�1"t'!(e1't   ��?    ����P>�*K�pL-��7�MC��7�_3��`A^8AS�� g�3�T0 k� ���ݑ�1"t'!(e1't   ��?    ����P>|*K�lL-��3�M?��7�_3��\A^8AS�� c�3�T0 k� ���ܑ�1"t'!(e1't   ��?    ����P>x*LhL-�/�M;��7�_/��\A^4AS�� c�3�T0 k� ���#ܑ�1"t'!(e1't   ��?    ����P>t)LdL-{�/�M;��7�_/��XA^0AS�� c�3�T0 k� ���#ۑ�1"t'!(e1't   ��?    ����P>p)L`L-{�+�M7��7�_+��TA^0AS�� c�3�T0 k� �#��'ۑ�1"t'!(e1't   ��?    ����P>l(L`L-w�'�M3��7�_+��TA^,
AS�� c�3�T0 k� �'��+ۑ�1"t'!(e1't   ��?    ����P>l(L\L-s�#�M/��7�_'��PA^(
AS�� c�3�T0 k� �'��+ڑ�1"t'!(e1't   ��?    ����P>h(LXL-o�#�M+��7�_'��LA^$	AS�� c�3�T0 k� �+��/ڑ�1"t'!(e1't   ��?    ����P>d'LTL-k��M+��7�_#��LA^$	AS�� c�3�T0 k� �/��3ّ�1"t'!(e1't   ��?    ����PNd'LPL-g��M'��7�_#��HA^ 	AS�� _�3�T0 k� �/��3ّ�1"t'!(e1't   ��?    ����PN`'LLL-g��M#��7�_��DA^AS�� _�3�T0 k� �3��7ؑ�1"t'!(e1't   ��?    ����PN\&LHL-c�/�=��7�_��DA^AS�� _�3�T0 k� �7��;ؑ�1"t'!(e1't   ��?    ����PN\&LHL-_�/�=��7�_��@A^AS�� _�3�T0 k� �7��;ב�1"t'!(e1't   ��?    ����PNX&LDL[�/�=��7�_��<A^AS�� _�3�T0 k� �;��?ב�1"t'!(e1't   ��?    ����PNT&L@L[�/�=��7�_��<A^AS�� _�3�T0 k� �?��C֑�1"t'!(e1't   ��?    ����PNT%L<LW�/�=��7�_��8A^AS�� _�3�T0 k� �?��C֑�1"t'!(e1't   ��?    ����PNP%L8LS�/�=��7�_��8A^AS�� _�3�T0 k� �C��G֑�1"t'!(e1't   ��?   ����PNL%L8LO�/�=��7�_��4A^AS�� _�3�T0 k� �G��KՑ�1"t'!(e1't   ��?    ����PNH$L4LO�/�=��7�_��0A^AS�� [�3�T0 k� �G��KՑ�1"t'!(e1't   ��?    ����PND$L0C�K�.��=��7�_��0A^AS�� [�3�T0 k� �K��Oԑ�1"t'!(e1't   ��?    ����PND$L0C�G�.��=��7�_��,A^AS�� [�3�T0 k� �O��Sԑ�1"t'!(e1't   ��?    ����PN@$L,C�C�.��=��7�_��,A^AS�� [�3�T0 k� �O��Sӑ�1"t'!(e1't   ��?    ����PN<#L(C�?�.������7�_��(A^AS�� [�3�T0 k� �S��Wӑ�1"t'!(e1't   ��?    ����PN8#L$C�;�.������7�_��(A^ AS�� [�3�T0 k� �W��[ґ�1"t'!(e1't   ��?    ����PN8#L$C�7�.������7�_��$A]�AS�� [�3�T0 k� �W��[ґ�1"t'!(e1't   ��?    ����PN4#L C�3�.������7�_��$A]�AS�� [�3�T0 k� �[��_ґ�1"t'!(e1't   ��?    ����PN0"L C�/�.�����7�_�� A]�AS�� [�3�T0 k� �_��cё�1"t'!(e1't   ��?   ����PN,"LC�+�.�����7�_�� A]�AS�� [�3�T0 k� �_��cё�1"t'!(e1't   ��?   ����PN,"LC�'�.�����7�_��A]�AS�� W�3�T0 k� �c��gБ�1"t'!(e1't   ��?    ����PN("LC�#�.�����7�_��A]�AS�� W�3�T0 k� �c��gБ�1"t'!(e1't   ��?    ����PN$!LI��.�����7�_��A]�AS�� W�3�T0 k� �g��kϑ�1"t'!(e1't   ��?    ����PN$!LI��.�����7�_��A]�AS�� W�3�T0 k� �k��oϑ�1"t'!(e1't   ��?   ����PN !LI��.��ߴ�7�^���A]�AS�� W�3�T0 k� �k��oϑ�1"t'!(e1't   ��?    ����PN!LI��.��߳�7�^���A]�AS�� W�3�T0 k� �o��sΑ�1"t'!(e1't   ��?    ����PN L	I��.��۲�7�^���A]�AS�� W�3�T0 k� �s��wΑ�1"t'!(e1't   ��?    ����PN L	I��.��ױ�7�^���A]�AS�� W�3�T0 k� �s��w͑�1"t'!(e1't   ��?    ����PN L	I��.��װ�7�^���A]� AS�� W�3�T0 k� �w��{͑�1"t'!(e1't   ��?    ����PN L	I��.��ӯ�7�^���A]� AS�� W�3�T0 k� �{��̑�1"t'!(e1't   ��?    ����PN L 	I���.��ӯ�7�^���A]� AS�� W�3�T0 k� �{��̑�1"t'!(e1't   ��?    ����PNL 	I���.��ϯ�7�^���A]� AS�� W�3�T0 k� ����̑�1"t'!(e1't   ��?    ����PNL�	I���.��Ϯ�7�^���A]��AS�� W�3�T0 k� ����ˑ�1"t'!(e1't   ��?    ����PNL�	I���.���˭�7�^���A]��AS�� W�3�T0 k� �����ˑ�1"t'!(e1't   ��?    ����PNL�	I���.���ǭ�7�^���A]��AS�� S�3�T0 k� �����ʑ�1"t'!(e1't   ��?    ����PNK��	I���.���Ǭ�7�^��A]��AS�� S�3�T0 k� �����ʑ�1"t'!(e1't   ��?    ����PNK��	I���.���ǫ�7�^�� A]��AS�� S�3�T0 k� �����ɑ�1"t'!(e1't   ��?    ����PNK��	I���.���ë�7�^�� A]��AS�� S�3�T0 k� �����ɑ�1"t'!(e1't   ��?    ����PN K��
I���.���ê�7�^�� A]��AS�� S�3�T0 k� �����ɑ�1"t'!(e1't   ��?    ����PN K��
I���.���é�7�^���A]��AS�� S�3�T0 k� �����ȑ�1"t'!(e1't   ��?    ����PM�K��
I���.���é�7�^���A]��AS�� S�3�T0 k� �����ȑ�1"t'!(e1't   ��?    ����PM�C��
I���.���é#,7�^���A]��AS�� S�3�T0 k� �����Ǒ�1"t'!(e1't   ��?    ����P=�C��
I���.�����#,7�^���A]��AS�� S�3�T0 k� �����Ǒ�1"t'!(e1't   ��?    ����P=�C��
A���.�����#,7�^���A]��AS�� S�3�T0 k� �����Ǒ�1"t'!(e1't   ��?   ����P=�C��	A��������#,7�^���A]��AS�� S�3�T0 k� �����Ƒ�1"t'!(e1't   ��?    ����P=�C��	A��������#,7�^���A]��AS�� S�3�T0 k� �����Ƒ�1"t'!(e1't   ��?    ����P=�C��	A��������#,7�^���A]��AS�� S�3�T0 k� �����ő�1"t'!(e1't   ��?    ����P=�C��	A��������#,7�^���A]��AS�� S�3�T0 k� �����ő�1"t'!(e1't   ��?    ����P=�C��A��������#,7�^���A]��AS�� S�3�T0 k� �����đ�1"t'!(e1't   ��?    ����P=�C��A���^�����#,7�^���A]��AS�� S�3�T0 k� �����đ�1"t'!(e1't   ��?    ����P=�C��A���^�����#,7�^���A]��AS�� O�3�T0 k� �����Ñ�1"t'!(e1't   ��?   ����P=�C��A���^������7�^���A]��AS�� O�3�T0 k� �����Ñ�1"t'!(e1't   ��?    ����P=�C��BL��^������7�^���
A]��AS�� O�3�T0 k� �����Ñ�1"t'!(e1't   ��?    ����P=�C��BM�^������7�^���
A]��AS�� O�3�T0 k� ������1"t'!(e1't   ��?    ����P=�C��BM�^������7�^���
A]��AS�� O�3�T0 k� ������1"t'!(e1't   ��?    ����P=�C��BM�^���å�7�^���
A]��AS�� O�3�T0 k� ��������1"t'!(e1't   ��?    ����P=�C��BM�^���ä�7�^���
A]��AS�� O�3�T0 k� ��������1"t'!(e1't   ��?    ����P=�C��F�^���Ǥ�7�^߳��
A]��AS�� O�3�T0 k� ��������1"t'!(e1't   ��?   ����P=�C��F�^���Ǥ�7�^߳��	A]��AS�� O�3�T0 k� ��������1"t'!(e1't   ��?    ����P=�C��F�^���Ǥ�7�^߳��	A]��AS�� O�3�T0 k� ��������1"t'!(e1't   ��?    ����P=�C��F�^���Ǥ�7�^߳��	A]��AS�� O�3�T0 k� �ǿ�˿��1"t'!(e1't   ��?    ����PM�C��F�^���ˤ�7�^߳��	A]��AS�� O�3�T0 k� �˿�Ͽ��1"t'!(e1't   ��?    ����PM�C��F�^���ˤ#7�^߳��	A]��AS�� O�3�T0 k� �˿�Ͽ��1"t'!(e1't   ��?    ����PM�C��F�^���ϣ#7�^۳��	A]��AS�� O�3�T0 k� �Ͼ�Ӿ��1"t'!(e1't   ��?    ����PM�C��F�^���ϣ#7�^۳��A]��AS�� O�3�T0 k� �Ӿ�׾��1"t'!(e1't   ��?    ����PM�C��F�^���ϣ#7�^۳��A]��AS�� O�3�T0 k� �ӽ�׽��1"t'!(e1't   ��?   ����PM�C��F�^���ӣ#7�^۳��A]��AS�� O�3�T0 k� �׽�۽��1"t'!(e1't   ��?    ����PM�C��F�^���ӣ#7�^۳��A]��AS�� O�3�T0 k� �׽�۽��1"t'!(e1't   ��?    ����PM�C��F�^���ע#7�^۳��A]��AS�� O�3�T0 k� �ۼ�߼��1"t'!(e1't   ��?    ����PM�C�� L}�^���ۢ#7�^۳��A]��AS�� O�3�T0 k� �߼�㼑�1"t'!(e1't   ��?    ����PM�C�� L}�^���ߢ#7�^׳��A]��AS�� O�3�T0 k� �߼�㼑�1"t'!(e1't   ��?    ����PM�C��L}�^���ߢ#7�^׳��A]��AS�� O�3�T0 k� ���绑�1"t'!(e1't   ��?    ����PM�C�w�L}�^���ߢ#7�^׳��A]��AS�� O�3�T0 k� ���绑�1"t'!(e1't   ��?    ����PM�C�s�L}#�^�����7�^׳��A]��AS�� O�3�T0 k� ���뺑�1"t'!(e1't   ��?    ����PM�C�k�L}#�^�����7�^׳��A]��AS�� K�3�T0 k� ���ﺑ�1"t'!(e1't   ��?    ����PM�C�g�L}'�^�����7�^׳��A]��AS�� K�3�T0 k� ���ﺑ�1"t'!(e1't   ��?    ����PM�C�_�L}+�^�����7�^׳��A]��AS�� K�3�T0 k� ���󹑕1"t'!(e1't   ��?    ����PM�C�[�L}+�^�����7�^ӳ��A]��AS�� K�3�T0 k� ���󹑕1"t'!(e1't   ��?    ����PM�C�S�L}/�^�����7�^ӳ��A]��AS�� K�3�T0 k� �������1"t'!(e1't   ��?    ����PM�C�O�L}/�^�����7�^ӳ��A]��AS�� K�3�T0 k� ��������1"t'!(e1't   ��?    ����PM�C�G�L}3�^�����7�^ӳ��A]��AS�� K�3�T0 k� ��������1"t'!(e1't   ��?    ����PM�C�C�L}7�^������7�^ӳ��A]��AS�� K�3�T0 k� ��������1"t'!(e1't   ��?    ����PM�C�;�L}7�^������7�^ӳ��A]��AS�� K�3�T0 k� ��������1"t'!(e1't   ��?   ����PM�C�3�L�;�^������7�^ӳ��A]��AS�� K�3�T0 k� �������1"t'!(e1't   ��?    ����PM�C�/�L�;�^������7�^ӳ��A]��AS�� K�3�T0 k� �������1"t'!(e1't   ��?    ����PM�C�'�L�?�^������7�^ӳ��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�C��L�?�^�����7�^ϳ��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�C��L�C�^�����7�^ϳ��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�C��L�G�^�����7�^ϳ��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�C��L�G�^�����7�^ϳ��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�C��L�K�^�����7�^ϳ��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�C���L�K�^�����7�^ϳ��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�C���L�O�^�����7�^ϳ��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�EM��L�O�^�����7�^ϳ��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�EM��L�S�^�����7�^ϳ��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�EM��L�S�^�����7�^˳��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�EM��L�W�^�����7�^˳��A]��AS�� K�3�T0 k� ������1"t'!(e1't   ��?    ����PM�EM��L�W�^�����7�^˳��A]��AS�� K�3�T0 k� ���#���1"t'!(e1't   ��?    ����PM�EM��L�[�^����7�^˳��A]��AS�� K�3�T0 k� ���#���1"t'!(e1't   ��?    ����PM�EM��L�[�^� ��7�^˳��A]��AS�� K�3�T0 k� �#��'���1"t'!(e1't   ��?    ����PM�EM��L�_�^� ��7�^˳��A]��AS�� K�3�T0 k� �#��'���1"t'!(e1't   ��?    ����PM�EM��L�_�^� ��7�^˳��A]��AS�� K�3�T0 k� �'��+���1"t'!(e1't   ��?    ����P=�EM��L�_�^� ��7�^˳��A]��AS�� K�3�T0 k� �+��/���1"t'!(e1't   ��?    ����P=�E=��L�c�^� ��7�^˳��A]��AS�� K�3�T0 k� �+��/���1"t'!(e1't   ��?    ����P=�E=��L�c�^{� ��7�^˳��A]��AS�� K�3�T0 k� �/��3���1"t'!(e1't   ��?    ����P=�E=��L�g�^{����7�^˳��A]��AS�� K�3�T0 k� �/��3���1"t'!(e1't   ��?    ����P=�E=��L�g�^{����7�^˳��A]��AS�� K�3�T0 k� �3��7���1"t'!(e1't   ��D    ����P=�E=��L�k�^{����7�^ǳ��A]��AS�� K�3�T0 k� �3��7���1"t'!(e1't   ��D    ����P=�E=��L�k��{����7�^ǳ��A]��AS�� K�3�T0 k� �3��7���1"t'!(e1't   ��D    ����P=�E={�L�k��w����7�^ǳ��A]��AS�� K�3�T0 k� �3��7���1"t'!(e1't   ��D    ����P=�E=s�L�o��w� ��7�^ǳ��A]��AS�� K�3�T0 k� �;��?���1"t'!(e1't   ��D    ����P=�E=o�L�o��s� ��7�^ǳ��A]��AS�� K�3�T0 k� �C��G���1"t'!(e1't   ��D    ����P=�E=g�L�o��s� ��7�^ǳ��A]��AS�� K�3�T0 k� �G��K���1"t'!(e1't   ��D   ����P=�CMc�L�s��o� ��7�^ǳ��A]��AS�� K�3�T0 k� �O��S���1"t'!(e1't   ��D    ����P=�CM[�L�s��o� ��7�^ǳ��A]��AS�� K�3�T0 k� �S��W���1"t'!(e1't   ��D    ����P=�CMW�L�w��k� ��7�^ǳ��A]��AS�� K�3�T0 k� �S��W���1"t'!(e1't   ��D    ����P=�CMO�L�w��k� ��7�^ǳ��A]��AS�� K�3�T0 k� �S��W���1"t'!(e1't   ��D    ����P=�CMK�L�w��g� ��7�^ǳ��A]��AS�� K�3�T0 k� �S��W���1"t'!(e1't   ��D    ����P�E=C�L�{�>g� ��7�^ǳ��A]��AS�� K�3�T0 k� �W��[���1"t'!(e1't   ��D    ����P�E=?�L�{�>c� ��7�^ǳ��A]��AS�� K�3�T0 k� �W��[���1"t'!(e1't   ��D    ����P�E=7�L�{�>_� ��7�^ǳ��A]��AS�� K�3�T0 k� �W��[���1"t'!(e1't   ��D    ����P�E=3�L��>_� ��7�^ǳ��A]��AS�� K�3�T0 k� �W��[���1"t'!(e1't   ��D    ����P�E=/�L��>[����7�^ó��A]��AS�� K�3�T0 k� �C��G���1"t'!(e1't   ��D    ����P=�E='�L��>[����7�^ó��A]��AS�� K�3�T0 k� �7��;���1"t'!(e1't   ��D    ����P=�E=#�L}��>W����7�^ó��A]��AS�� K�3�T0 k� �+��/���1"t'!(e1't   ��D    ����P=�E=�L}��>W����7�^ó��A]��AS�� K�3�T0 k� �#��'���1"t'!(e1't   ��D    ����P=�E-�L}��>S����7�^ó��A]��AS�� G�3�T0 k� ���#���1"t'!(e1't   ��D    ����P=�E-�L}��>S����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D   ����P=�E-�L}��>O����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����P=|E-�L}��>O����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����P=xE-�BM��>K����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����P=xK��BM��NK����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����P=tK��BM��NG����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����P=tK��BM��NG����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����P=pK��BM��NC����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����P=p
K���E}��NC����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMl
K���E}��N?����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMh	K���E}��N?����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMh	K���E}��N?����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMdK��E}��N;����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMdK��Em��N;����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PM`K��Em��N7����7�^ó��A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PM`K��Em��N7����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PM\K��Em��N7����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PM\K��Em��N3����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMXK��Em��N3����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMXK�ߣE]��N/����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMXK�ߢE]��N/����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMTK�ۢE]��N/����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMTK�סE]��N+����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMPK�סE]��N+����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMPK�ӠE]��N+����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMLK�ӟEM��N'����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMLK�ϟEM��N'����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMLK�˞EM��N'����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMHK�˞EM��N#����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMHK�ǝEM��N#����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMDK�ǝEM��N#����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMDK�ÜEM��N����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PMDK�ÜEM��N����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����PM@ K̿�EM��N����7�^����A]��AS�� G�3�T0 k� ������1"t'!(e1't   ��D    ����P a�jS���Ea����9���l;��ǽ��NE���B�D"7�3��T0 k� ������1"t'!(e1't   ��/    ��� � a�jS���Ea��� :���l;��Ͼ��NE���B�L"7�3��T0 k� ������1"t'!(e1't   ��/   ��� � �jS���Ea���:���l;��׿мNE���B�T"7�3��T0 k� ������1"t'!(e1't   ��/    ��� � �jS���Ea���;���l;������ME��B�h"7�3��T0 k� ��	��	��1"t'!(e1't   ��/    ��� � �jS���Ea��� ;���l;������ME��B�p"7�3��T0 k� ��	��	��1"t'!(e1't   ��/    ��� � �jS���Ea���(<���l;������LE�#�B�x�7�3��T0 k� ��	��	��1"t'!(e1't   ��/    ��� ���jS���EQ���0<��l;������LE�+�B���7�3� T0 k� ��
� 
��1"t'!(e1't   ��/    ��� ���jS���EQ���8=��l;�����LE�3�B���7�3� T0 k� �
�
��1"t'!(e1't   ��/    ��� ���jS���EQ���L=��l;����KE�G�B���7�3� T0 k� ����1"t'!(e1't   ��/    ��� ���jS���EQ���T>�#�l;�#��KE�O�B���7�3�T0 k� �� ��1"t'!(e1't   ��/    ��� ��jS���EQ���\>�+�l;�+��JEs[�B���;�3�T0 k� �$�(��1"t'!(e1't   ��/    ��� ��jS���EQ���h>�/�l;�3��JEsc�B���;�3�T0 k� �,�0��1"t'!(e1't   ��/    ��� ��iS���EQ���p?�7�l;�;��IEsk�B���;�3�T0 k� �4�8��1"t'!(e1't   ��/    ��� ��iS���EQ���x?�?�l;�C�� IEss�B���;�3�T0 k� �<�@��1"t'!(e1't   ��/    ��� ���iS���EQ����@�O�l;��S��0HPӇ�B���?�3�T0 k� �L�P��1"t'!(e1't   ��/    ��� ���iS���EQ��Δ@�W�l;��[��8GPӏ�B��C�3�T0 k� �T�X��1"t'!(e1't   ��/    ��� ���hS���EQ��ΠA�[�l;��g��@GPӗ�B��C�3�T0 k� �X�\��1"t'!(e1't   ��/    ��� ���hS���EQ��ΨA�c�l;��o��HFPӟ�B��G�3�T0 k� �`�d��1"t'!(e1't   ��/    ��� ���hS���EQ��ΰA�k�l;��w��PFPӧ�B��G�3�T0 k� �h�l��1"t'!(e1't   ��/    ��� �q�gS���EQ��μB�s�l;����XEPӯ�B�K�3�T0 k� �p�t��1"t'!(e1't   ��/    ��� �q�gS���EQ����B�{�l;�����\EP��B�K�3�T0 k� �x�|��1"t'!(e1't   ��/    ��� �q�fS���EQ����Bދ�l;�����lCP���B�O�3�
T0 k� �����1"t'!(e1't   ��/    ��� �q�eS���EQ����Cޓ�l;�ѣ��tCP���B�(�S�3�
T0 k� �����1"t'!(e1't   ��/    ��� �q�dS���EQ����C���l;�ѫ��|BP���B�0�W�3�T0 k� �����1"t'!(e1't   ��/    ��� �q�cS���EQ����C���l;�ѳ��AP���B�8�W�3�T0 k� �����1"t'!(e1't   ��/    ��� �a�cS���EQ����D���l;�ѻ��AP��B�@�[�3�T0 k� �����1"t'!(e1't   ��+    ��� �a�bS���EQ���D���l;�����@P��B�H�[�s�T0 k� �����1"t'!(e1't   ��+    ��� �a�`S�� EQ���E���l;�����?P���B�\�_�s�T0 k� �����1"t'!(e1't   ��+    ��� �a�_S�� EQ��� E���l;����	�>P��B�d�c�s�T0 k� �����1"t'!(e1't   ��+    ��� 1�^S��A����,E���l;����	�>P��B�l�c�s�T0 k� �����1"t'!(e1't   ��+    ��� 1�]S��A����4E���l;����	�=P��B�t�g�s�T0 k� �����1"t'!(e1't   ��+    ��� 1�[S��A����HF���l;���	��<P��B҈Bk�s�T0 k� �����1"t'!(e1't   ��+    ��� 1�ZS��A����PF���l;���	��<P�#�BҐBo���T0 k� �����1"t'!(e1't   ��+    ��� 2 YS� A���XF���l;���
�;Et+�BҘBo���T0 k� �����1"t'!(e1't   ��+    ��� 2 XS� A���dG���l;���
�;Et/�BҠBs���T0 k� �����1"t'!(e1't   ��+    ��� 2 US�A���tG��l;�r/�
�:Et?�BҰ"w���T0 k� �����1"t'!(e1't   ��+    ��� �B TS�A����G��l;�r7�
�:EtC�BҸ"{�øT0 k� �����1"t'!(e1't   ��+    ��� �B SS�BA����H��l;�r7�	��:EtK�I�"�øT0 k� �����1"t'!(e1't   ��+    ��� �B RS�BA����H��l;�r;�	��:EtO�I�"��ôT0 k� �����1"t'!(e1't   ��+    ��� �B OS�BA����H�/�l;�rG�	��9Et[�I�"��ðT0 k� �����1"t'!(e1't   ��+    ��� �b NS�BA����I�7�l;�rK�	��9Ed_�I���ìT0 k� �|����1"t'!(e1't   �+    ��� �b LS�D�����I�?�l;�rO�
�9Edg�I�����T0 k� �p	�t	��1"t'!(e1't   ��/    ��� �a�KS�D�����I�G�l;�BS�
 9Edk�I"�����T0 k� �h�l��1"t'!(e1't   ��/    ��� �a�KS�D�����J�W�l;�B_�
8Eds�I"�����T0 k� �T�X��1"t'!(e1't   ��/    ��� ���KS�D�����J�_�l;�Bc�
7Edw�I# 	2����T0 k� �O��S���1"t'!(e1't   ��/    ��� ���JS�D�����J�c�l;�Bg�	�7Ed{�I#	2����T0 k� �C��G���1"t'!(e1't   ��/    ��� ���IS�D�����J�k�l;�o�	�6Ed�I	2����T0 k� �;��?���1"t'!(e1't   ��/    ��� ���IS�	D�����J�s�l;�s�	�6Ed��I	2����T0 k� �/��3���1"t'!(e1't   ��/    ��� ���GS� 	D����J���l;��	�5Ed��I 	B����T0 k� ����1"t'!(e1't   ��/    ��� ���FS� 
D����K���l;���� 4Ed��I(	B����T0 k� ����1"t'!(e1't   ��/    ��� ���EU2 
D����K���l;�����$4ET��E�,	B����T0 k� ���1"t'!(e1't   ��/    ��� ���DU2$
D����(K���l;�����(3ET��E�4	B����T0 k� �����둕1"t'!(e1't   ��*    ��� ��BU2(D����8J���l;�����02ET��E�@	2����T0 k� �����쑕1"t'!(e1't   ��*    ��� ��AU2(D����DJ���l;�����41ET��E�H	2����T0 k� �����푕1"t'!(e1't   ��*    ��� ��?U2(D����LJ���l;����r80ET��E�H	2����T0 k� �����푕1"t'!(e1't   ��*    ��� ��>U2,D����TJ���l;����r<0ET��E�L	2����T0 k� �����1"t'!(e1't   ��*    ��� ��=U2,F���`J���l;����r@/ET��E�L	2����T0 k� �����1"t'!(e1't   ��*    ��� ��<U2,F���hJ���l;����rD.ET��E�P	B����T0 k� �����1"t'!(e1't   ��*    ��� ��9U20F���|I���l;��˸rL,C��E�X	B����T0 k� �����1"t'!(e1't   ��*    ��� ��8E"0F��ЄI���l;��ӸrP+C��E�\	B����T0 k� �����1"t'!(e1't   ��*    ��� ���7E"4F��ЌI���l;�	۷rP*C��E\	B����T0 k� ����1"t'!(e1't   ��*    ��� �� 5E"4F�ИH���l;�	�rT)C��E`	2����T0 k� ����1"t'!(e1't   ��*    ��� �� 4E"8F�РH���l;�	�rX(C��Ed	2����T0 k� ����1"t'!(e1't   ��*    ��� ��2E�<D��дG �l;�	�r`%C��Ed	2����T0 k� ����1"t'!(e1't   ��*    ��� ��0E�@D���G �l;�	��bd$C��E�h	2����T0 k� ����1"t'!(e1't   ��*    ��� ��/E�DD����F �l;�	"��bd#C��E�l	B����T0 k� ����1"t'!(e1't   ��*    ��� ��.E�HD� ��F �l;�	#�bh!C��E�p	B����T0 k� ����1"t'!(e1't   ��*    ��� ��,E�PD���E /�l;�	#�blC��E�x	B����T0 k� ����1"t'!(e1't   ��*    ��� ��+E�TD���D 3�l;�	#�blC��I�|	B��3�T0 k� ����1"t'!(e1't   ��    ��� ��)E�XD� ��D ;�l;�	�bpC�{�I�	2��3�T0 k� ����1"t'!(e1't   ��    ��� �� (E�\D�$��CC�l;�	�btC�w�I�	2��3�T0 k� ����1"t'!(e1't   ��    ��� ��(&E�`D�$�BS�l;�	#�bxC�o�I�	2��3�T0 k� ����1"t'!(e1't   ��    ��� ��,%E�`D�$�AW�l;�	'�b|C�k�J�	2��3�T0 k� ����1"t'!(e1't   ��    ��� ��0$E�`D�(� A_�l;�	#+�R�C�g�J���3�T0 k� ������1"t'!(e1't   ��    ��� ��4$E�dD�(�(@g�l;�	#/�R�C�c�J���3�T0 k� ������1"t'!(e1't   ��    ��� ��@"E�hD�(�<?w�l;�	#7�R�C�[�J���3�T0 k� ������1"t'!(e1't   ��    ��� ��D!E�lD�(qD>�l;�	#;�R�C�W�I���3�T0 k� ������1"t'!(e1't   ��    ��� ��H!E�p
D�,qL=��l;�	;�R�DS�I�R��3�T0 k� �����푕1"t'!(e1't   ��    ��� ��H!E�p	D�,qT<��l;�	?�R�DO�I�R��3�T0 k� �����ꑕ1"t'!(e1't   ��    ��� ��L!E�tD�0qh;��l;�	C�R�DC�I�R��3�T0 k� ����葕1"t'!(e1't   ��    ��� ��P C�tD�0qp:	��l;�	G�B�D?�J�R��3�T0 k� ����瑕1"t'!(e1't   ��    ��� ��T C�xD�0qx8	��"�;�	#K�B�D7�J�
R��3�T0 k� ����摕1"t'!(e1't   ��    ��� ��X C�xD�4q�7	��"�;�	#K�B�D3�J�
���3�T0 k� ����㑕1"t'!(e1't   ��    ��� ��\ C�xD�4q�6	��"�;�	#K�B�D+�J�
���3�T0 k� ��������1"t'!(e1't   ��    ��� ��d C�xD�8q�4	��"�;�	#O�B�D�@�
���3�T0 k� �����ޑ�1"t'!(e1't   ��    ��� ��h C�|D�8q�2	 ��"�;�	S�B�D�@�	���3�T0 k� �����ݑ�1"t'!(e1't   ��    ��� ��l C�| E�8q�1	 ��"�;�	S�B�D�@�	���3�T0 k� �����ۑ�1"t'!(e1't   ��    ��� ��l C��E�<a�0	 ��"�;�	S�B�D�@����3�T0 k� ����ؑ�1"t'!(e1't   ��    ��� ��p C�{�E�<	a�-	 ��"�;�	W�B�D��E�����3�T0 k� ����ב�1"t'!(e1't   ��    ��� ��t!C�{�E�@	a�+	��"�;�	#W���D��E�����3�T0 k� ����֑�1"t'!(e1't   ��    ��� ��x!C�{�Er@	a�*	��l;�	#W���D��E�����3�T0 k� ����ԑ�1"t'!(e1't   ��    ��� ���"C�w�ErDa�'	��l;�	#W���D��E�����3�T0 k� ����ӑ�1"t'!(e1't   ��    ��� �B�#C�w�ErHa�%	��l;�	#W���D��E�����3�T0 k� ����ґ�1"t'!(e1't   ��    ��� �B�#C�w�ErHa�$	 ��l;�	W���D��E�����3�T0 k� ����ё�1"t'!(e1't   ��    ��� �B�%C�s�ErLa� 	 ��l;�	W���D��E�� ���3�T0 k� ����Б�1"t'!(e1't   ��    ��� �B�&C�o�ErPa�	!�l;�	W���C��E������3�	T0 k� ����ϑ�1"t'!(e1't   ��    ��� �B�'C�o�ErPa�	!�l;�	W���C��E������3�T0 k� ����Α�1"t'!(e1't   ��    ��� �B�(C�k�EbPQ�	�l;� �W���C��E������3�T0 k� ����Α�1"t'!(e1't   ��    ��� �B�)E2g�EbTQ�	�l;� �W���C��E������3�T0 k� ����̑�1"t'!(e1't   ��    ��� �R�+E2c�EbTR 	�"�;� �W���C��Eã����3�T0 k� ����ˑ�1"t'!(e1't   ��    ��� �R�,E2c�EbXR	�"�;� �W���C�{�Eã����3�T0 k� ����ˑ�1"t'!(e1't   ��    ��� �R�.E2_�EbX�	!�"�;�W���I�g�Eã����3�T0 k� ����ȑ�1"t'!(e1't   ��    ��� R�/E2[�EbX�	!�"�;�W���I�_�Eã�ҿ�3�T0 k� ����Ƒ�1"t'!(e1't   ��    ��� }R�1E2[�EbX�	!�"�;�W���I�W�C���һ�3� T0 k� ����ő�1"t'!(e1't   ��    ��� {R�2E2W�EbT�	!�"�;�W���I�O�C���һ�c� T0 k� ����đ�1"t'!(e1't   ��    ��� yR�5E2S�ERT�
	�"�;�W�ҔI�?�C���ҳ�c��T0 k� �w��{�1"t'!(e1't   ��    ��� wR�6E2O�ERP�		#�"�;�W�ҔI�7�C���ү�c��T0 k� �s��w���1"t'!(e1't   ��    ��� uR�8E2O�ERP�	#�"�;�SW�ҐI�/�E3��ҫ�c��T0 k� �o��s���1"t'!(e1't   ��    ��� sb�9E2K�ERL�	#�l;�SW�ҐI�+�E3��ҧ�c��T0 k� �k��o���1"t'!(e1't   ��    ��� qb�=E2G�ERH!�	!'�l;�SW�ҌI��E3��ҟ�c��T0 k� �c��g���1"t'!(e1't   ��    ��� ob�>E2G�ERD"�	!'�l;�SW�҈E��E3����c��T0 k� �_��c���1"t'!(e1't   ��    ��� mb�@E"G�ER@#� 	!'�l;��W�҄E��E3����c��T0 k� �[��_���1"t'!(e1't   ��    ��� k��BE"C�ER<$��	!'�l;��S�҄E��E3����c��T0 k� �W��[���1"t'!(e1't   ��    ��� i��EE"C�ER4&��	'�l;��O��|E���E3����c��T0 k� �K��O���1"t'!(e1't   ��    ��� g��GE"?�ER0'��	'�l;��O��x E���IS����c��T0 k� �G��K���1"t'!(e1't   ��    ��� e��IE"?�ER,(��	'�l;��K��t E���IS����c��T0 k� �C��G���1"t'!(e1't   ��    ��� c��KE"?�EB()��	'�l;��K��p!E���IS��Rw�c��T0 k� �G��K���1"t'!(e1't   ��    ��� a��ME"?�EB$*�	'�l;��G��l!E���IS��Rw�c��T0 k� �G��K���1"t'!(e1't   ��    ��� _��QP2;�EB,� a'�l;��C��d"E���IS��Ro�c��T0 k� �C��G���1"t'!(e1't   ��    ��� ]��SP2;�EB-�� a'�l;��?��`#D2��Ic��Rg�c��T0 k� �C��G���1"t'!(e1't   ��    ��� [��VP27�C�-�� a'�l;��;��X#D2��Ic��Rc�c��T0 k� �?��C���1"t'!(e1't   ��    ��� Y��XP27�C�.�� a'�l;��7��T$D2��Ic��R_�c��T0 k� �;��?�1"t'!(e1't   ��:    ��� W��\P23�C� /Q�� �'�l;��/��L%D2��Ic��RS�c��T0 k� �/��3���1"t'!(e1't   ��:    ��� U��^PB3�C��0Q�� �'�l;��+��D%D2��IS��RO�c��T0 k� �+��/���1"t'!(e1't   ��:    ��� S��`PB3�C��0Q�� �'�l;��'��@&D2��IS��RG�c��T0 k� �#��'���1"t'!(e1't   ��:    ��� Q��bPB3�C��0Q�� �'�l;��#��8&D2��IS��RC�c��T0 k� ���#���1"t'!(e1't   ��:    ��� O��ePB/�C��1Q�� �'�l;����4'D2�IS��R;�c��T0 k� ������1"t'!(e1't   ��:    ��� M��gPB/�C��1Q��'�l;���,'D2w�IS��R7�c��T0 k� ������1"t'!(e1't   ��:    ��� K��kPB/�C��2Q��'�l;��� (D2c�Ic��R'�c��T0 k� ������1"t'!(e1't   ��:    ��� I��mPB+�C��2Q��'�l;���(DB[�Ic��B#�c��T0 k� �������1"t'!(e1't   ��:    ��� G��oPB+�C��2Q��'�l;���)DBS�Ic��B�c��T0 k� ��������1"t'!(e1't   ��:    ��� E��rP2+�C��2Q��'�l;����)DBK�Ic��B�c��T0 k� ��������1"t'!(e1't   ��:    ��� C��tP2+�C��2A��Q'�l;����)DBC�Ic��B�c��T0 k� ��������1"t'!(e1't   ��:    ��� A��vP2'�C��2A��Q'�l;��� *DB;�IS��B�c��T0 k� ��������1"t'!(e1't   ��:    ��� ?��zP2'�C��2A��Q'�l;���+DB'�IS��a��c��T0 k� �ӿ�׿��1"t'!(e1't   ��:    ��� =��|E"'�C��1A��Q'�l;���+DB�IS��a�c��T0 k� �Ͼ�Ӿ��1"t'!(e1't   ��:    ��� ;��}E"'�C��1A���'�l;�۳�+DB�IS��a�c��T0 k� �Ǿ�˾��1"t'!(e1't   ��:    ��� 9��E"'�C��1A���#�l;�׳�,DB�Ic��a�c��T0 k� �ý�ǽ��1"t'!(e1't   ��:    ��� 7�܁E"'�C��1A���#�l;�ϳ�,DB�Ic��a߮c��T0 k� ������1"t'!(e1't   ��:    ��� 5�ԀE'�C��0A����l;����-DQ��Ic��aӭc��T0 k� ������1"t'!(e1't   ��:    ��� 3�ԀE'�C�|0A{���l;����-DQ��Ic��Qϭc��T0 k� ������1"t'!(e1't   ��:    ��� 1��E'�C�t/As���l;����.DQ��IS��QǬc��T0 k� ������1"t'!(e1't   ��:    ��� /��E+�C�l/Ao���l;����.DQ��IS��Që3��T0 k� ������1"t'!(e1't   ��:    ��� -��E+�C�d.1g���l;����.DQ��IS��Q��3��T0 k� ������1"t'!(e1't   ��:    ��� +��~E+�C�\.1_���l;����/DQ��IS��Q��3��T0 k� ������1"t'!(e1't   ��:    ��� )Ҽ}E�/�C�P,1S���l;����/DQ��Ic��A��3��T0 k� ������1"t'!(e1't   ��:    ��� '�}E�3�C�H,1K���l;�⃳�0DQ��Ic��A��3��T0 k� �������1"t'!(e1't   ��:    ��� &�|E�7�C�@+1G���l;��{��0DQ��Ic��A��3��T0 k� �{�����1"t'!(e1't   ��:    ��� %                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��vJ ]�4�4� X �*  ��   � �	   ��P·     ?��Q!%    �-�r           m���P�         ���    ���  8

�          ����  � �
	   ��/�^    ����0)
    �]�   
       s ���P�         ��    ���  0

           ����  T T    �bo0    ���i�cT    ��p          ���P�        
0�  �  ���   (
"          ���e   � �	    ��S�    �������    ����   	         %���P          ��  
  ���  H
w          ����   � �
      .�C��    ��/��C�E    �y��           e
 ���P            �    ���   (
         ��m  ��
      B�|�    ��m�|�           	                  ���_              \  ���    0

 2            ���:          V��b~    ���:��i�      ��            q =         -0     ��@   8
(          Y�    	     j�l�      `�l��    ���N           	   :         �      ��@   @


         ��ɖ        ~�cY    �����cM    ���L          
�� �         ��     ��@    

'           ����  �	   � ��W    ���� ��W                     	�� �         	 �     ��@   8

          ��y   x	     � Ɇ    ��y ��      ��           
     �         
 �      ��J   X
          [+ ��
	     � �=i     [+ �=i                          ���y        �@   +  ��@    0 0                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         ���[  ��        ��CM�    ���P�CSb    �y�� "                 x                j  �       �                         ��    ��       ��D      ��  �D           "                                                 �                         �P�/�b���C����l�c �  ����C�D    
    	         
    I~ ?��G       ;� ``� <� a� <� a� <�  a� �d _� �� _� ɤ  ]  �� ]` �� d� Ǆ  d@ �� d� �� d� �  d� �� p� �d  x� פ x� $� �o� %� p� 
�< V� 
�< V� 
�| W  
�� W� 
�\ W� � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }` 
�| W� 
� W� 
�\ W����� � 
�\ W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����P������ �  ������  
�fD
��L���"����D" � j  "  B   J jF�"     
�j 
 ���
��
��"     "�j��   * �
� �  �  
� ����  ��     ��C      ����  ��     ��C      ����  ��     �           � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �D      ��0 �  ���        � � �  ��        �        ��        �        ��        � 
 
 f�
    �����        ��                         �$ ( � ��                                    �                 ����           ���C
���%��  ���P��                5 Nicklas Lidstrom    1:57                                                                        5  5     � �
� �2�!2�8CBCD$ CL �J� � � J� � 	J� � �
J� � � J� � � J� � � � � �C. � �C4 � �C8 � � � � �B�4 � B�: �B�- �B�5 � B�= �k~$ � k�$ �K � � K � � K � �K � �cj6 � cr. �C �  C" �!C#  �"C% � #C' |$cV � � %c^ �&"� � '"� � �(� � �)
� �*"� � +"� � �,"� � �-*� � �."  y �/!� y � 0"@ y � 1"O � � 2"J � � 3"K � � 4"B �5"  y  6" �(7!� yP 8"I �`  "P � }:!� u;", u *L { *L ~>"- ~ *$M                                                                                                                                                                                                                         �� R @      �    @ 
         �     b P E e  ��        
            �������������������������������������� ���������	�
��������                                                                                          ��    ��K�� ��������������������������������������������������������   �4, 8  H �� ����@�@���A+�?�J�s������������                                                                                                                                                                                                                                                                                                  �@�                                                                                                                                                                                                                                             4    6    � �  .�J     W�                             ������������������������������������������������������                                                                                                                                    �  ��                �        �   �            	     ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� �������           g      	          T        � �  4�J      =m  	                           ������������������������������������������������������                                                                                                                                 
       ]  �   )  �                  ��               	 
     ��  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���                                                                                                                                                                                                                                                  	                                                               
        �             


            �   }�                 }�  y�                                          y�                         ��������    ����  + ����   ����������������  V��������������������  N���������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" R > / 	                                � �W� �\        �U�!&R�1U1'                                                                                                                                                                                                                                                             )n)nY  
1F        c            k                  m            `                                                                                                                                                                                                                                                                                                                                                                                                         > �  >�  <�  @8  H#�  EZmt ������0�= �N @��� i�����"����������������        .  �� � : ��          �   & AG� �   `   
           A\�                                                                                                                                                                                                                                                                                                                                     _ X    m    
   	             !��                                                                                                                                                                                                                            Y��   �� � Ѱ��      �� X      ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� ���������  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���      �     $��˼��̼���˻̼�̻�̻�˼�����̼�l�˼����k���������̺��˼���f��ff��˻������˻���f��ff�fffffffffff��̼��l��fflffffffflffffffffffff���˻��̼���˻̼f̼�f˻��l��fl̼�k����̻���̻�˼���˼̼������˼�����˻̼���˻�������������˻����ʦff��ff��ff�fff�ffȼffw�ff��ff�ffffff�ff�z�lx�w��w�xuwX�uwwwwuWfffffffl����wWWUww��xWwWuwuwxWwUff��fl�ˆf�lXf�fw�ffwVflwYffWyff̼�̻̼���k˻������˼�˼���̼��˪����������������˻��������������ff��ff��ff��ffw�ffw��fW���W���W�u�w�wWuwUwWwuUU��k��xƺx�hɋ�ȧ�wuww�wWuxwuUWUUwW���y��ux�i�U�gxxflwY�lwxfkWwfl�ufk��f˩�Ǽ�w�������̼̻�k̻������̼�̻̼�����˺�����������������������ʪ���������w��������fgw��jU����x��fw�ffw����wWxxwwwwuwxXww��wwz�����wwww�u��wwxw�ww��xXWwW���x�W����wxXW�w��WYy�w�WfwXY�w�|�xu��wwf�wVk�����̼̻���̻������̻���˻�˻���˺�������������������������������ffw�ffw��fw��fw���w���U�������Ww�wuwwwzwx��w����xxy���xX���ux�uUWUw��ww���w���x��w���wxuUw�UUX�xVj�wV̻u�k�w�����˻����u���U�˻��̼���������������̻������˻�������˺��˺���������U̧UU�UW�U{�����u���w���w�X�wX�XwU[�w˵�U��Yuww��wuw�wwU�WWWuwWwwWWWXuuuwUWUUw��u��uW��wuUWWWwwwu�wXWwuuUuUWUu���U�˻u���u���u�{\W��Uu���Wuū�˻�������̼����l���z�̼�|�˻����m�    ?      2   � ��                       X        ���������J    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$     `d  �@���6 ��  �@���6 �$ ���  ��       � �N ^$   ��  ����  ��  ����  �$ ^$��    �     
^V        *   3� � ��� �� � ��� �$  � �  �� �  �      �   d   6���� e����J   g��� 	        f ^�         �� b��      6      ��v��������J���J������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                                             �                       �e iV�U�i                    ��������eeY�                 fU��Ul���ř�Yf�    V  UY e�V ��P �Uf Ŗf f�U                �  �  �\  �� 
]�    �U�eVl�Vl�f�f��f�iUl�f��VfU��f�V�����Ɯfli��e�fl\�Vf\ilVlUV����eU������elfl��fl�Y��eUV��f�e��fU�UVf�feYfU�l�fUVf�f�feUfY�l�ffP \UU �eP fe� �V  i`  V   `    \l �l� ��� ��l ��V �lV \e 
V��ll��V�fVllUVYlefll��VlfleVeV�eU��e����f�l���flf��V��f�ff��\l\UleU��f�fVlU�l�f�fY�feleU`iU` U`  �leZfeV eU` ej  V                                �                �l   e                       Uf��leUUV�eUeY�� Y�            eeV�Ul�Plƕ �e` �`              P                                                                                             wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            """ "!   " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                              """ "!   " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       """ "!   " ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                          �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                   �     �                         � �������������  �                                                                                                                                       "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��             �  �˰ ��� �wp ���                            ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                     �� ���
�������˽������̽�]��+I۲"T�""T32.T33>@4C CDT �E@ ��  ʐ  �       "   "�� � ��� �wp ��� �vz �w� �����˻���˰�̰� ��  ��  ��� � �+ �+ �  .   "�   �   �   �    � ��  �                     �  �˰ ���                 ��  ��  ���           U   U  U  U  	T  ,� ,� "  " "  ��  �                �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����            �����                         �     �                                       �   ���                            �   �                                                                                                     �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                            �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                  ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .   ��  �   ��  �                                  ���                � ���� ��   � � �                           �   �                                                                                                              �  ��� ��� ��� �ݪ�                       �   �    �z� 
�� ������������ ˍ� ��� ���������ˉ����� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��                    ˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                                         �  ��  �� ��  ��        �   �     �   �                                                   �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  ��  ��  �                       ���  +"  "" ���������                   �                        ���� ��� ����                              "  .���"    �     �                                          ����     �   �  �  �  ��  �   �                                                                                                        �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                ��� ���� ��    �     �                                                                                                                                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                  �� ��� ��                      "   "   "  �� ��                   ����������             ��  �   ��  �                    ��   �  ��  �  �  �         � �������������  �                                                                                                                                                 �   �  
� 
�� ���	���    �   ��  ��  �ڠ rj� gj��w���������������˽,̲" �""  "  
�  
�   �   �   J   
           ����̻ۻ�˽��˽�̻��뻽���K���RDD>�UD4NUDD�T4�K 3˸ Ȣ   "" �   �   �   �   �   �   "   "   "   "   ".  C � ;� �ˊ  ��  
�"         0    "    0      " �/����      �             "�"�����   �� �          ����   �       �                                   �    ���  ��                    ��  ��  ���                   ���                � �������������  �                                                                                                                                         �� ̚�
���	��������� �ܷ �� +� "� "+  ��UH"+��""��"+���   ��  ̸� ��� �͌��ݩ�g���gz��w���ت��ݚ���ɜЉ��К˽ ȭ� ��9 �UB �UB �T@ ED/ ��� ��� ������   ""  ""� �  �� ��   ��                                         � ��                +��"�"/� ""� "" �   �             ��  ���  �                      � ����  �                                 �                 ���� ��� ����                               � ��                  �  �˰ ��� �wp ���                       ����     �   �  �  �  ��  �   �                                                                                                               �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��                  �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""����������D��M��M""""����������""""�����ADMA����""""����DD�M�""""��������AD�DM�""""�����������A�A�""""������AD�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��M��M�������D����3333DDDD�DD�M�D�������3333DDDDD�������M�DM�D����3333DDDD��A�M�M���M�����3333DDDDMM������D��D����3333DDDDA�A�A�D��M�D�����3333DDDD�������������D������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=LL����������D����3333DDDD    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����������A������ x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx""""�������I�I������ w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww""""�������I��D���I�������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(�D�M�D���M������3333DDDD �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""�����AMAD������ M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M""""������������������ � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�fFfFDfFFfFffdFffff3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DDFFDfFFfdFffff3333DDDD 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5""""wwwwwwwGGD x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x""""wwwwwwqwAqwAwA w w x y�������H���������������������������������H������yxww""""wwwwqwqAwAqAqAq  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(A�A�A�A��LD�����3333DDDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,�A�LDL�L�D�L�����3333DDDD +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+""""wwwwwwDGAD 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5""""wwwwqqDAAq =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
� �2�!2�8CBCD$ CL �J� � � J� � 	J� � �
J� � � J� � � J� � � � � �C. � �C4 � �C8 � � � � �B�4 � B�: �B�- �B�5 � B�= �k~$ � k�$ �K � � K � � K � �K � �cj6 � cr. �C �  C" �!C#  �"C% � #C' |$cV � � %c^ �&"� � '"� � �(� � �)
� �*"� � +"� � �,"� � �-*� � �."  y �/!� y � 0"@ y � 1"O � � 2"J � � 3"K � � 4"B �5"  y  6" �(7!� yP 8"I �`  "P � }:!� u;", u *L { *L ~>"- ~ *$M3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������.�O�T�U��-�O�I�I�G�X�K�R�R�O� � � � � �.�/�=�����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3����������������������������������������� ��8�O�I�Q�R�G�Y��6�O�J�Y�Z�X�U�S� � � � �.�/�=�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������-�2�3� �� �������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������.�/�=� ��"������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            