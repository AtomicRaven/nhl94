GST@�                                                           �[�                                                      #��     �              ����e J���J�����������p�������        �g      #    ����                                d8<n    �  ?     Ra����  �
fD�
�L���"����D"� j   " B   J  jF�"    
 �j� � 
 ���
��
�"   "D�j��
� " ��
  �                                                                               ����������������������������������      ��    bbo QQ g 11 44               		� 

                      ��                      nn� ))         888�����������������������������������������������������������������������������������������������������������������������������=o  0  4o  1    +     '           �                    �	  �7  �V  �	                  n  	          : �����������������������������������������������������������������������������                                �z  �   s  E�   @  #   �   �                                                                                '     )n)n�  	n    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE 7 �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    E^�gMXo��? l�,a� 	 �P[�,3��1A�g�BB�T0 k� �s��w�e2D# 3I)@5   ��O    � <�hE^�gMTo��? m�(a� 	 �P[�,3��1A�k�BB�T0 k� �s��w�e2D# 3I)@5   ��O    � <�hE^|hMTo��?�n�(a� 	 �O[�,3��1A�k�BB�T0 k� �w��{�e2D# 3I)@5   ��O    � <�hENthMTo��>�p�(a� 	 �O[�,3��1A�k�BB�T0 k� �{���e2D# 3I)@5   ��O    � <�hENhhMTo��>�q�(a� 	 �O[�,3��1A�k�BB�T0 k� �{���e2D# 3I)@5   ��O    � <�hEN`iMPo��>�r�(a� 	 �N[�-3��1A�k�BB�T0 k� �����e2D# 3I)@5   ��O    � <�hENXiMPo��>�s�$a� 	 �N[�-3��1A�k�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hENPiMPo��>�u�$a� 	 �N[�-"���1A�k�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hC�DjMPo��=�v�$a� 	 �M[�-"���1A�k�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hC�<jMLo��=�w�$`� 	 �M[�-"���1A�k�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hC�4jMLo��=�x�$`� 	 �M[�-"���1A�k�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hC�,kMLo��=�y�$`� 	 �L[�-"���1A�k�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hC� kMLo��=�z�$`� 	 �L[�-"���1A�k�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK�kMHo��<�| � `� 	 �L[�-"���1A�k�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK�kMHo��<�} � `� 	 �L[�."���1A�k�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK�lMHo��<�~ � `� 	 �K[�."���1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK��lMHo��<� � `� 	 �K[�."���1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK��lMHo��<� � `� 	 �K[�."���1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK��mMDo��<� � `� 	 �J[�.3��1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK��mMDo��<� � `� 	 �J[�.3��1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK��mMDo��<� �`� 	 �J[�.3��1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK��mMDo��<� �`� 	 �J[�.3��1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK��nMDo��<� �`� 	 �I[�.3��1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK��nM@o��<�~ �`� 	 �I[�/3��1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK��nM@o��<�~ �`� 	 �I[�/3��1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hK��oM@o� <�~ �`� 	 �I[�/3��1A�o�BB�T0 k� ������e2D# 3I)@5   ��O   � <�hL�oM@o�=�~ �_� 	 �H[�/3��1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL�oM@o�=�} �_� 	 �H[�/3��1A�o�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hE=pk,S�>_�\�<��|8 �\k�3���<Dm��C���T0 k� �  � e2D# 3I)@5   ��    ����JE-hi,O�>W�\�<��|<�Pl�3���4Dm��C�{�T0 k� � !�!e2D# 3I)@5   ��    ����JE-`h,K�>O�\�<ü|<>Hl�3���,Dm�D s�T0 k� � #�#e2D# 3I)@5   ��    ����JE-\g,G�>K�\�<ý|<>@l�3���$Dm{�D k�T0 k� � %�%e2D# 3I)@5   ��    ����JE-Tf,C�>C�\�<ǿ!�<>8l�"s���Dms�D c�T0 k� � &�&e2D# 3I)@5   ��    ����JE-Pe,?�>;�\�<��!�@>0l�"s���Dmk�D [�T0 k� � (�(e2D# 3I)@5   ��    ����KE-Db,7�N+�\�<��!�@> l�"s��� Dm_�D K�T0 k� �+�+e2D# 3I)@5   ��    ����KE-@a,3�N#�\�L��!�@>l�"s�� �DmW�D C�T0 k� �,�,e2D# 3I)@5   ��    ����KE-8_,/�N�L�L��!�D>l�"s�� �D=S�D ;�T0 k� �.�.e2D# 3I)@5   ��    ����KE-4^,+�N�L�L��!�D>l�"s�� �D=K�D 3�T0 k� �/�/e2D# 3I)@5   ��    ����KE-0],+�N�L�L��!�D> l�"s�� �D=G�D +�T0 k� �1�1e2D# 3I)@5   ��    ����KE-(Z,'�N�L�L��!�D=�l�!"s�� �D=7�D �T0 k� �4�4e2D# 3I)@5   ��    ����KE-$X,#�M��L�L��!�DM�l""s�� �D=3�D�T0 k� �5�5e2D# 3I)@5   ��    ����KE-$W,�M�L�L��|DM�k$3�� �E�+�D�T0 k� �7�7e2D# 3I)@5   ��    ����KE- U,�M�L�L��|DM�k%3�� �E�'�D�T0 k� �8�8e2D# 3I)@5   ��    ����KE-T�M�L�L��|DM�k&3�� �E��D��T0 k� �9�9e2D# 3I)@5   ��    ����KEQ�M��L�L��|HM�k)3�� �E��D��T0 k� ��5��5e2D# 3I)@5   �    ����IEO�]��L� \��|HM�j*3���E��D��T0 k� ��3��3e2D# 3I)@5  ��    ����GEM�]��L��\��|HM�j,3���E��D��T0 k� ��1��1e2D# 3I)@5  ��    ����FEL�]��<��\��|HM�j-3���E���D��T0 k� ��/��/e2D# 3I)@5  ��    ����EEK�]��<��\��|LM�i.3��xE���D��T0 k� ��-��-e2D# 3I)@5  ��    ����DEH�=��<��<��|L	M�i13��hE��D��T0 k� �l)�p)e2D# 3I)@5  ��    ����CEF =��<��<��|L	]�h.23��`E��E_��T0 k� �X'�\'e2D# 3I)@5  ��    ����BB�E�=��L��<��|L	]|h.33��XE��E_��T0 k� �D%�H%e2D# 3I)@5  ��    ����AB�D�=��L{�<��|L	]tg.43��LE�۷E_��T0 k� �0#�4#e2D# 3I)@5  ��    ����@B�B�=��Lw�<��|L
]lg.53��DE�׸E_��T0 k� �!� !e2D# 3I)@5  ��    ����?B�@�=��Lo�<��|P	]\f.83��4E�˻EO��T0 k� ����e2D# 3I)@5  ��    ����>B�>�-��Lo�,��|P
]Tf.93���,E�üEO��T0 k� ����e2D# 3I)@5  ��    ����=B�=�-��Lk�,��|P
]Le.:3���$E���EO�T0 k� ����e2D# 3I)@5  ��    ����<B�<�-��<g�,��|T
]De.;3���E���EOw�T0 k� ����e2D# 3I)@5  ��    ����;B�:�-��<c�,���P
]<d.<3���E���EOo�T0 k� ����e2D# 3I)@5  ��    ����:B�8�-�<[�,���P
](d.>3��� D���C�_�T0 k� ����e2D# 3I)@5  �    ����9B�7�	-{�<W�,���P
] c.?3����D���C�W�T0 k� ,|��e2D# 3I)@5  ��    ����8E�6�	-w�<S�,���P
�c.@3����D���C�O�T0 k� ,x�|e2D# 3I)@5  ��    ����8E�4�	-s�<O�,� �P
�c.A3����D���C�K�T0 k� ,x�|e2D# 3I)@5  ��    ����8E� 3	-o�<K�- �P
�b.B3����D���C�C�T0 k� ,t�xe2D# 3I)@5  ��    ����8E�$2	�o�,G�-�P
� b.C3����E���C�;�T0 k� ,p�te2D# 3I)@5  ��    ����8E�(/�g�,?�-�T
��a.E3����E���C�+�T0 k� ,l�pe2D# 3I)@5  ��    ����8E�,.�g�,;�	=
�T
��a.F3����E��C�#�T0 k� �h�le2D# 3I)@5  ��    ����8E�0,�c�,;�	=�T
��a.G3����E�{�C��T0 k� �d�he2D# 3I)@5  ��    ����8E�4+-c��7�	=�T
��`>H3����Fw�C��T0 k� �d�he2D# 3I)@5  ��    ����8E�8)-c��3�	=�T
��`>I3����Fs�C��T0 k� �`�de2D# 3I)@5  ��    ����8B�@&-_��/�	=�T
��_>K3����Fk�EN��T0 k� �X�\e2D# 3I)@5  ��    ����8B�@%�-_��/�	M�T
�_>L3����Fg�EN��T0 k� <X�\e2D# 3I)@5  ��    ����8B�D$�-[��+�	M�T
�_>M3����Fc�EN��T0 k� <T�Xe2D# 3I)@5  ��    ����8B�H"�-X�+�	M�X
�^>O3���xF_�EN��T0 k� <P�Te2D# 3I)@5  ��    ����8I=P � -X�'�	M�X
�]. Q3���dFW�EN��T0 k� <L�Pe2D# 3I)@5  ��    ����8I=P�$-X�$ 	=�X
�]. S3��\FW�EN��T0 k� �H �L e2D# 3I)@5  ��    ����8I=T�$X
$ 	=�X
�\. T3��TFS�EN��T0 k� �D!�H!e2D# 3I)@5  ��    ����8I=X�(X
  	=�X
�\. U3��LFO�EN��T0 k� �D"�H"e2D# 3I)@5  ��    ����8IM\�0\ 	=�\
�p[.$X3��<FK�EN��T0 k� �<#�@#e2D# 3I)@5  ��    ����8IM`�4\ 	M�\
�hZ.(Z3��_0FK�EN��T0 k� ,8$�<$e2D# 3I)@5  ��    ����8IMd�8\ 	M�\
�`Z.([3��_(FG�E>��T0 k� ,8%�<%e2D# 3I)@5  ��    ����8IMd �<\ 	M�\
�XY.(]3��_ E�G�E>��T0 k� ,4&�8&e2D# 3I)@5  ��    ����8I=h!�D` 	M �`
�HX.0`3��_E�C�E>��T0 k� ,0'�4'e2D# 3I)@5  ��    ����8I=l!�L�d� 	=!�`
�@W.0b3��_E�C�E>��T0 k� �,(�0(e2D# 3I)@5  ��    �  �8I=l"�P�d� 	=!�`
�8W4c3��_ E�C�E>�T0 k� �()�,)e2D# 3I)@5  ��    � �8I=p"�X�l� 	="�`
�(U8g3��^�E�C�E>s�T0 k� �$+�(+e2D# 3I)@5  ��    � �8IMp#�`�l� 		=#|`
� T<h3��^�E�C�E>k�T0 k� �(� (e2D# 3I)@5  ��3    � �8IMp#�d�p< 		M#|`�S@j3��^�E�C�E>c�T0 k� L&� &e2D# 3I)@5  ��3    � �8IMt$p!�t< 		M$|`�QHm3��N�E�C�E>W�T0 k� L%� %e2D# 3I)@5  ��3    � �8IMt$t!�x< 		M$|`�PLn3��N�E�C�E>S�T0 k� L#� #e2D# 3I)@5  ��3    � �8Ex$|"�|< 
	M$�`��OPp3��N�E�G�E>K�T0 k� L#� #e2D# 3I)@5  ��3    � �8Ex$�"��,	=%�`��NTq3��N�E�G�E.G�T0 k� � !�$!e2D# 3I)@5  ��3    � �8E�%�$��,	=%�`��K`t3��N�E�G�E.;�T0 k� �$"�("e2D# 3I)@5  ��3    � �8E�%�$��,	=%�`�Jdv3��N�E�G�E.3�T0 k� �$!�(!e2D# 3I)@5  ��3    � �8E�%�%��,	=%�\�Ilw3��N�E�G�E./�T0 k� �$"�("e2D# 3I)@5   ��3    � �8E��&�&���	M&�\�Ftz3��N�E�H E.'�T0 k� ,&� &e2D# 3I)@5   -�3    � �8E��&�'���	M&�\�E|{3��NxE�HE.#�T0 k� ,(�(e2D# 3I)@5   ��3    � �8E��'�'ݠ�	M&�\�C�|3��NpE�HE.�T0 k� ,*�*e2D# 3I)@5   ��3    � �8E��(��(ݨ�	M&�X�@�3��N\E�LE.�T0 k� ,.�.e2D# 3I)@5  ��3    � �8Dݜ(��)ݬ� �&�X�?��3��>TE�LE.�T0 k� �0�0e2D# 3I)@5  ��3    � �8Dݠ)��)ݰ� �%�X�=���3��>LE�PE.�T0 k� �2�2e2D# 3I)@5  ��3    � �8Dݬ*��*ݼ�" �%�P�:��3��><E�PE.�T0 k� �6�6e2D# 3I)@5  ��3    � �8Dݰ+��*���$ � %�L�9��3��>4E�TE�T0 k� �8�8e2D# 3I)@5  ��3    � �8Dݴ,��+���&�$%�Hۤ7��3��>,CLTE��T0 k� <8�8e2D# 3I)@5  ��3    � �8Dݸ-��+���(�$&�D۠6��~3��>$ CLTE��T0 k� <9�9e2D# 3I)@5  ��3    � �8D��.��+���,�,&�@ۜ2��~3��>"CLXE��T0 k� < <�<e2D# 3I)@5  ��3    � �8D��/��,���.�0&�8ۘ1��~3��>"CLXB���T0 k� < =�=e2D# 3I)@5  ��3    � �8D��0��,���0�4&�4�/��}3��>#CL\B���T0 k� � >�>e2D# 3I)@5  ��3    � �8D��2��,���4�8'�,�,��}3��>#CL\B��T0 k� ��B� Be2D# 3I)@5  ��3    � �8D��4��,���6�<'�(�,��|3��>$CL\B��T0 k� ��D��De2D# 3I)@5  ��3    � �8D��5��,���8�<(�$�,� |3��. $CL`B��T0 k� ��F��Fe2D# 3I)@5  ��3    � �8D��7��,� �9�@(�$��-�|3��-�%CL`B��T0 k� +�G��Ge2D# 3I)@5   ��3    � �8D��;��,�L=�D)���-�{3��-�&CLdB��T0 k� +�L��Le2D# 3I)@5   ��3    � 	�8D��=� ,�
L?�H)���.� {3��-�&C\dB��T0 k� +�N��Ne2D# 3I)@5   ��3    � 
�8D��?� ,�	LA�L*���.�({3��-�'C\d B��T0 k� +�P��Pe2D# 3I)@5   /�3    � �8D��A�,� LC�L*���.�0{3��-�(C\d B��T0 k� ��R��Re2D# 3I)@5   ��3    � �8D�D�,�,K�G�P+���/�@z3��-�)C\k�B��T0 k� ��V��Ve2D# 3I)@5   ��3    � �8D�F�,�4K�I�T+���0�Hz3��-�*C\k�B��T0 k� ��X��Xe2D# 3I)@5   ��3    � �8D�H�,�<K�K�T+���0�Tz3���*C\k�B��T0 k� ��Z��Ze2D# 3I)@5   ��3    � �8E�J�,�D;�M�X+���1�\y3���+C\o�B��T0 k� ��\��\e2D# 3I)@5   ��3    � �8E�M�+�P;�Q�\,���2�ly3���-C\o�B���T0 k� ��a��ae2D# 3I)@5   ��3    � �8E�$O�+�X ;�S�\,���3�ty3���-C\o�B���T0 k� ��d��de2D# 3I)@5   ��3    � �8E�(Q�*�c�;�U�\,� ��3�|y3����.Cls�B���T0 k� ��f��fe2D# 3I)@5   ��3    � �8E�0R�*�k�;�W�`,� ��4τx3����/Cls�B���T0 k� ��h��he2D# 3I)@5   ��3    � �8E�4T� *�s�;�Y�`,� ��5όx3����/Cls�B���T0 k� ��j��je2D# 3I)@5   ��3    � �8E�@W� *��;�\�d,����6Ϡx3����1Clw�B��T0 k� ��n��ne2D# 3I)@5   ��3    � �8E�HY�$*���;�^=d,����7Ϩw3����1Clw�B��T0 k� ��p��pe2D# 3I)@5   ��3    � �8E�P[�$)~��;�`=d,����8߰w3����2Clw�B��T0 k� ��r��re2D# 3I)@5   ��3    � �8E�T\�$)~��;�b=h+����9߸w3����3Clw�B��T0 k� ��t��te2D# 3I)@5   ��3    � �8E�\^�$(~��+�d=h+����:��w3����3E�w�B��T0 k� ��u��ue2D# 3I)@5   ��3    � �8E�d_�('~��+�f=h+����;��w3����4E�{�B��T0 k� ��v��ve2D# 3I)@5   ��3    � �8E�pb�('~��+�j=l+����=��v3����5E�{�B��T0 k� ��y��ye2D# 3I)@5  �3    �  �<E�xd(&~��+�l=l*���>��v3����6E�{�B��T0 k� �z�ze2D# 3I)@5  ��?    � !�@E�|e,%~����n=l*���?	�v3����6E��B�#�T0 k� �{�{e2D# 3I)@5  ��?    � "�DE��g,$~����p=l)���@	�v3����7E��B�'�T0 k� � }�$}e2D# 3I)@5  ��?    � #�HE��h,$�����q=p)���A	�v3����8E��B�+�T0 k� �,~�0~e2D# 3I)@5  ��?    � $�LE��i,#�����s=p)���B	 v3����8E��B�/�T0 k� �8�<e2D# 3I)@5  ��?    � %�PE��k0"�����uMp(���C	v3����9E��B�3�T0 k� �D��H�e2D# 3I)@5  ��?    � &�TE��l0!�����uMp(���E	v3����9E��B�7�T0 k� �T��X�e2D# 3I)@5  ��?    � '�XE��n4 �����uMp'���F	 v3����:Ẽ�B�;�T0 k� �`��d�e2D# 3I)@5  *�? 	   � (�\E��o8~����uMp'���H	 v3����:Ẽ�B�C�T0 k� �l��p�e2D# 3I)@5  ��? 	   � )�`E��q8~����uMp&����J	  v3����;Ẽ�B�G�T0 k� �x��|�e2D# 3I)@5  ��? 	   � *�dE��t<~����u]p&����O	 (v3����<E<��B�O�T0 k� ̔����e2D# 3I)@5  ��? 	   � +�hE��u�@~����v]p&����Q	0v3����<E<��B�W�T0 k� ̠����e2D# 3I)@5  ��? 	   � ,�lE��v�D���v]p&����S	4v3����=E<��B�[�T0 k� ̬����e2D# 3I)@5  ��? 	   � -�pE��x�H���v]p&����V	8v3��� =E<��B�_�T0 k� ܼ����e2D# 3I)@5  ��? 	   � .�tE��y�H���v]p&����X	<v3���>E<��B�g�T0 k� �Ȃ�̂e2D# 3I)@5  ��? 	   � /�xE��{�Lo���vMl%� ��Z	Dv3���>E<��B�k�T0 k� �Ԃ�؂e2D# 3I)@5  ��? 	   � 0�|E��|�Po���vMl%� ��\	 Hv3���?E<��B�s�T0 k� �����e2D# 3I)@5  ��? 	   � 1��E��~�To���vMl%� �^	 Lv3���?CL��B�w�T0 k� �����e2D# 3I)@5  ��? 	   � 2��E���Xo#���vMh%� �`	 Pv3���@CL��B��T0 k� ���� �e2D# 3I)@5   ��? 	   � 3��E����\o'�� vMh%��b	 Pv3���@CL��B���T0 k� ����e2D# 3I)@5   ,�?    � 4��E� ��`o+��v=h%��d	 Tv3��� ACL��B���T0 k� ����e2D# 3I)@5   ��?    � 5��E���do/��v=d&��f	Xv3���(ACL��B���T0 k� � ��$�e2D# 3I)@5   ��?    � 6��E��ho3��v=d&��f	\v3���,BE<��B���T0 k� �0��4�e2D# 3I)@5   ��?    � 7��E��lo3��w=d&��$g	`v3���0BE<��B���T0 k� �<��@�e2D# 3I)@5  ��?    � 8��E��po7��w=`&��(h	`v3���8BE<��B���T0 k� �H��L�e2D# 3I)@5  ��?    � 9��E� ~�x
_;��xM`'��0i	dv3���<CE<��B���T0 k� �T��X�e2D# 3I)@5  ��?    � :��E�(~�|	_;��xM`'��8j	 dv3���DCE<��B���T0 k� �`��d�e2D# 3I)@5  ��?    � ;��E�,~��_?��yM`(��@l	 hv3���HDE<��B���T0 k� �p��t�e2D# 3I)@5  ��?    � <��E�4}��_?��yM\(��Dm	 hv3���PDE,��B���T0 k� |����e2D# 3I)@5  ��?    � <��E�8}��_C��yM\)��Ln	 lv3���TDE,��B�ǁT0 k� �����e2D# 3I)@5  ��?    � <��E�H|��_C��xMX*��Xp	 lv3���`EE,��E׀T0 k� �����e2D# 3I)@5  ��?    � <��E�L|��_G� lxMX+��`q	pv3���hEE,��EۀT0 k� �����e2D# 3I)@5  ��?    � <��E�T|��_G� lxMX,��dr	pv3���pFE,��E�T0 k� ݼ��e2D# 3I)@5  ��?    � <��E�X{��_G� lwMX-��ls	pv3���tFE,��E�T0 k� ����e2D# 3I)@5  ��?    � <��E�`{�� _G� lwMT.��pt	pv3���|GE,��E�T0 k� ����e2D# 3I)@5  ��?    � <��E�d{���_G� l w�T/��xu	tv3����GE,��E��T0 k� ����e2D# 3I)@5  ��?    � <��E�lz���OG�, w�T0��|w	 tv3����GE,��E�T0 k� ����e2D# 3I)@5  ��?    � <��E�tz���OG�,$w�P0���x	 tv3����HE,��E�T0 k� �� e2D# 3I)@5  ��?    � <��E�xz���OG�,(w�P1���y	 tv3����HE,��E�T0 k� �e2D# 3I)@5  ��?    � <��E��y���OC�,(v�L2���y	 tv3����HE,��E�T0 k� ~�~e2D# 3I)@5   ��?    � <��E��y���OC�,,v�L4���z	 tv3����IE,��E�#�T0 k� $~�(~e2D# 3I)@5   ��?    � <��E��x���OC�0v�H5���{ `tv3����IE��E�+�T0 k� 0~�4~e2D# 3I)@5   ��?    � <��E��x���OC�0v�H6���| `tv3����IE��E�3�T0 k� �<~�@~e2D# 3I)@5   ��?    � <��E��x���O?�4v�D7���} `tv3����JE��E�;�T0 k� �H~�L~e2D# 3I)@5   /�?    � <��E��w���O?�4u�D8���~ `tv3����JE��E�C�T0 k� �T~�X~e2D# 3I)@5   ��?    � <��E��w��O;�8u�@9��� `tv3����JE��E�K�T0 k� �`~�d~e2D# 3I)@5   ��?    � <��E��w��?;� <u�<:���� �tv3����JE��E�S�T0 k� �p~�t~e2D# 3I)@5   ��?    � <��E��v��?;� <u�8;���� �tv3����KE��E�W�T0 k� �|}��}e2D# 3I)@5   ��?    � <��E��v��?7� @u�8<��� �tv3����KE��E�_�T0 k� Έ}��}e2D# 3I)@5   ��?    � <��E��v�#�?7� @u�4=��� �tv3����KE��E�g�T0 k� Δ}��}e2D# 3I)@5   ��?    � <��E��u�+�?3� Dt�0>��� �tv3����LE��D�o�T0 k� Π}��}e2D# 3I)@5   ��?    � <��E��u�/�?3� Dt�,?��� tv3���LB���D�w�T0 k� ά}��}e2D# 3I)@5   ��?    � <��E��u�7�?3� Ht�(@���~ tv3���LB���D��T0 k� ��}��}e2D# 3I)@5   ��?    � <��E��u�?�?/� Ht�$A���~ tv3���LB���D߇�T0 k� ��}��}e2D# 3I)@5   ��?    � <��E��t�G�?/� Lt� B�%<�~ tv3���MB���Dߏ�T0 k� ��}��}e2D# 3I)@5   ��?    � <��E��t�O�?/� Lt�C�%<�~ tv3���$MB�ÄDߗ�T0 k� ��|��|e2D# 3I)@5   ��?    � < E��t�W�?+� Pt�C�%<�}Ptv3���,MB�ǃDߟ�T0 k� ��|��|e2D# 3I)@5   ��?    � < E��s�_�/+� Ps�D�%<�}Ptv3���4MB�ˁDߧ�T0 k� ��|��|e2D# 3I)@5   ��?    � < E��s�g�/+� Ts�E� %<�}Ptv3���@NB�πD߫�T0 k� �|�|e2D# 3I)@5   ��?    � < E��s�o�/'� Ts�F� %<�}Ppv3���HNB�׀D߳�T0 k� �|�|e2D# 3I)@5   ��?    � < E� r�w�/'� Xs� F� %<�|Phv3���PNB�ہD߻�T0 k� �|� |e2D# 3I)@5   ��?    � < E�r��/'� Xs��G� %<�|�dv3���XNB�߁D�ÍT0 k� �(|�,|e2D# 3I)@5   ��?    � < E�r���/'� \s��G� %=|�\v3���`OB��D�ˎT0 k� �4|�8|e2D# 3I)@5   ��?    � < E�q����'� \s��G�$%=|�Tv3���hOB��D�ӎT0 k� �D{�H{e2D# 3I)@5   ��?    � < E�q����'� `s��H�$%={�Tv3���pOB��D�ۏT0 k� �P{�T{e2D# 3I)@5   �?    � < Qp����'� `r��H�$%={�Pv3���|OB��D��T0 k� �\{�`{e2D# 3I)@5   ��?    � <  Qo����'� `r��H�$%={PPv"s��߄OB���D��T0 k� �h{�l{e2D# 3I)@5   ��?    � < #Qn����'� dr��I�$%={PLw"s��ߌPB���D��T0 k� �t{�x{e2D# 3I)@5   ��?    � < &Qm����+� dr��I�$%=zPLw"s��ߔPB��D���T0 k� ��{��{e2D# 3I)@5   ��?    � < )Ql����+� hr��I�$%= zPHw"s��ߜPB��D���T0 k� ��{��{e2D# 3I)@5   ��?    � < ,Qk����+� hr��I�$%=$zPHw"s��ߤPB��D��T0 k� ��{��{e2D# 3I)@5   ��?    � < /Qj����+� hr��I�(%=(zPHw"s��߬QB��D��T0 k� ��z��ze2D# 3I)@5   ��?    � < 2Qi����/� lr��H�(%=,yPDw"s����QB��D��T0 k� ��z��ze2D# 3I)@5   ��?    � < 5Q h����/�lr��H�(%=0yPDx"s����QB�'�D��T0 k� ��z��ze2D# 3I)@5   ��    � < 8Q g����/�pq��H�(%=4yPDx"s����QB�+�D�#�T0 k� ��z��ze2D# 3I)@5   ��    � < ;Q f���3�pq��H�(%=8yP@x"s����QB�3�D�+�T0 k� ��z��ze2D# 3I)@5   ��   � < >Q e���3�tq��G|(%=<xP@x"s����QB�;�D�3�T0 k� ��z��ze2D# 3I)@5   ��   � < AQ d���7�xq��G|(%=@xP@x3����RB�?�D�7�T0 k� ��z��ze2D# 3I)@5   ��   � < DQ c��7��xq��F|(%=DxP<x3����RB�G�D�?�T0 k� ��z��ze2D# 3I)@5   ��    � < GQ a��;��|q��F|(%=HwP<y3����RB�O�D�G�T0 k� �y�ye2D# 3I)@5   ��    � < JQ0a��;���p��E|(%=LwP8y3����QB�W�D�O�T0 k� �y�ye2D# 3I)@5   ��    � < MQ0a��?���p��E|(%=PwP8y3��� QB�_�D�S�T0 k� �y� ye2D# 3I)@5   ��    � < PQ0b�#�C���p��D|(%=PwP8y3���PB�g�D�[�T0 k� �(y�,ye2D# 3I)@5   $�    � < NQ0b�+�C���o��C|(%=TwP8y3� �PB�k�D�c�T0 k� �$y�(ye2D# 3I)@5   ��    � < LQ0b�3�G�|�o��B|(%=XvP4y3� �OB�s�E k�T0 k� �$y�(ye2D# 3I)@5   ��    � < KQ0b�;�K�|�o��B|(%=\vP4y3� � OB�{�E o�T0 k� �$y�(ye2D# 3I)@5   ��    � < JQ0b�?�O�|�n��A|(�`vP4z3��(NB݃�E w�T0 k� �$y�(ye2D# 3I)@5   ��    � < IQ0b�G�S�|�n��@|(�dvP0z3��0NB݋�E �T0 k� � y�$ye2D# 3I)@5   ��    � < HQ0 b�K�S�|�m��?|(�dvP0z"���8NBݓ�E ��T0 k� � y�$ye2D# 3I)@5   ��    � < GQ0$b�W�[�|�l�|=|(
�lvP,z"���HMBݟ�E ��T0 k� � y�$ye2D# 3I)@5   ��    � < FQ0(b�[�_�|�k�x<|(
�pv�,z"���PLBݧ�E ��T0 k� � y�$ye2D# 3I)@5   ��    � < EQ0(b?_�c�|�j�t;|(	�tu�,z"���XLBݯ�E ��T0 k� �x�xe2D# 3I)@5   ��    � < CQ0,b?g�g���i�p9|(	�xu�(z"���dLBݷ�E ��T0 k� �x�xe2D# 3I)@5   ��    � < AQ0,b?k�k���h�p8|(�xu�${"���lLBݿ�E ��T0 k� �x�xe2D# 3I)@5   ��    � < ?Q00b?o�o���g�l7|(�|u�${"���tKB�ǊDз�T0 k� �y�ye2D# 3I)@5   ��    � < =Q00b?s�s���f�h5|(-�t@ {"���|KB�ˊDл�T0 k� �~�~e2D# 3I)@5   ��    � < ;Q04b?w�/w���e�d4|(-�t@{"����KB�ӊD�ìT0 k� � ���e2D# 3I)@5   ��    � < 9Q08b?��/�|�c�`1|(-�t@z"����KB��D�ϮT0 k� ���� �e2D# 3I)@5   ��    � < 6Q0<b?��/��|�b�\0|(-�t@z3���KB��D�ׯT0 k� ������e2D# 3I)@5   ��    � < 3Q0<b?��/��|�a�X.|(-�t@z3� �KB��D�߰T0 k� �����e2D# 3I)@5   ��    � < 0Q0@b?�����|�`�T-|(�s@y3� �KB���D��T0 k� �����e2D# 3I)@5   ��    � < -Q0@b?�����|�^�T+|(�sy3� �KB���D��T0 k� ����e2D# 3I)@5   ��    � < *Q0Db?�����|�]�P)|(�sy3� �KB��D��T0 k� �܇���e2D# 3I)@5   ��    � < 'Q0Db/�����|�\�L(|(�sy3� �JB��D���T0 k� �ԇ�؇e2D# 3I)@5   ��    � < $Q0Hb/�����|�ZH&�(�s x3�0�JB��D���T0 k� �̆�Іe2D# 3I)@5   ��    � < !Q0Lb/� ���l�WD"�(��s�x3�0�IB�'�D��T0 k� ����Će2D# 3I)@5   ��    � < Q0Pb/�O��l�VD!�(��s�x3�0�IB�/�D��T0 k� ������e2D# 3I)@5   ��    � < Q0Pb��O��l�U@�(��s�w3�0�HB�3�D��T0 k� ������e2D# 3I)@5   ��    � < Q0Tb��O��l�S@�(��s�w3�0�HB�;�D�#�T0 k� ������e2D# 3I)@5   ��    � < Q0Tb��O��l�Q<�(��s�w3�0�GB�C�D�'�T0 k� ������e2D# 3I)@5   ��    � < Q0Xb��O��l�P<�(��s�w3�0�GB�K�D�/�T0 k� ������e2D# 3I)@5   ��    � < Q0\b��
���l�M<�(��s�v3�1FB�[�D�;�T0 k� ������e2D# 3I)@5   ��    � < Q0`b�����l�K<�$��r/�v3�1EEc�D�C�T0 k� ������e2D# 3I)@5   ��    � < Q0`b�����l�J<�$��r/�v3�1EEg�D�G�T0 k� ������e2D# 3I)@5   ��    � <  Q0db�����l�H�<�$��r/�u3�1DEo�D�O�T0 k� ������e2D# 3I)@5   ��    � <��Q0db�����\�F�<� ��r/�u3�1$DEw�D�S�T0 k� ������e2D# 3I)@5   ��    � <��Q0hb�����\�C�@� �rߴu3�10CE��D�c�T0 k� ����e2D# 3I)@5   ��    � <��Q0lb�����\�B�@!� �r߬t3�14BE��D�g�T0 k� ��{��{e2D# 3I)@5   ��    � <��Q0lb�����\�@�@!� �rߨt3�1<BE��D�o�T0 k� ��x��xe2D# 3I)@5   ��    � <��Q0pb�������>�@!� �rߠt3�1@BE��D�s�T0 k� �xv�|ve2D# 3I)@5   ��    � <��Q0pb�������=�@!� �$rߘt3�1HAE��D�w�T0 k� �pt�tte2D# 3I)@5   ��    � <��Q0tb�������;�D!��,rߐs3�1LAE��D��T0 k� �ls�pse2D# 3I)@5   ��    � <��Q0xb�� �����9�D!� �4rߌs3�1T@E���D��T0 k� �dr�hre2D# 3I)@5   ��    � <��Q0|b��$�����6�L!� �Dr�|s3�1\?E�ÏD��T0 k� �Tq�Xqe2D# 3I)@5   ��    � <��Q0|b��&�����4�L!��Lr�ts3�1d?E�ǏE��T0 k� �Lp�Ppe2D# 3I)@5   ��    � <��Q0�b��(�����2�P!��Tr�lr3�1h?E�ϏE��T0 k� �Dp�Hpe2D# 3I)@5   ��    � <��Q0�b��*�����0�T!� 	\r�dr3�1l>I�׏E��T0 k� �<p�@pe2D# 3I)@5   ��    � <��Q0�b��,�����.�T� 	dr�\r3�1t>I�ۏE��T0 k� �8k�<ke2D# 3I)@5   ��    � <��Q0�b�.����,�X� 	hr�Tr3�1x>I��E��T0 k� �0f�4fe2D# 3I)@5   ��    � <��Q0�b�0����*�\� 	pr�Lq3�1|=I��E��T0 k� �(c�,ce2D# 3I)@5   ��    � <��Q0�b�2����(�\� 	tr�Dq3�1�=I��E��T0 k� � a�$ae2D# 3I)@5   ��    � <��Q0�b�3����&�`� 	.|r�<p3�1�<J�E��T0 k� �^�^e2D# 3I)@5   ��    � <��Q0�bp 5����$�`� 	.�r�4p3�1�<J��E��T0 k� �]�]e2D# 3I)@5   ��    � <��Q0�bp 7����#�`� 	.�r�,p3�1�<J��E��T0 k� �[�[e2D# 3I)@5   ��    � <��Q0�b� 9�� �!�d� 	.�r�$o3�1�;J��E��T0 k� ��\� \e2D# 3I)@5   ��    � <��Q0�b�;����d� 	.�r�n3�1�;J�E��T0 k� ��\��\e2D# 3I)@5   ��    � <��Q0�b�<����d� ��r�n3�1�;E��E��T0 k� ��]��]e2D# 3I)@5   ��    � <��Q0�b�>����d� ��r�m3�1�:E��E��T0 k� ��]��]e2D# 3I)@5   ��    � <��Q0�b�@��	��h!� 	��r�m3�1�:E��E��T0 k� ��]��]e2D# 3I)@5   ��    � <��Q0�b�A�����h!� 	��r��l3�1�:E��E��T0 k� ��\��\e2D# 3I)@5   ��    � <��Q0�b�C�����h!� 	��s��l3�1�:E��E��T0 k� ��\��\e2D# 3I)@5   ��    � <��Q0�b�E�����h!� 	��s��k3�1�9E�#�E��T0 k� ��\��\e2D# 3I)@5   ��    � <��Q0�b�F�����h!� 	��s��j3�1�9E�+�E��T0 k� ��[��[e2D# 3I)@5   ��    � <��Q0�bpH�����h!� 	��t��i3�1�9E/�E��T0 k� ��Z��Ze2D# 3I)@5   ��    � <�~Q0�bpI����Lh!� 	��u��g3�1�8E3�E��T0 k� ��X��Xe2D# 3I)@5   ��    � <�|Q0�bpK����Lh!� 	��v��f3�1�8E7�E��T0 k� ��W��We2D# 3I)@5   ��    � <�zQ0�bpL����
Lh!� 	��u��d3�1�8E?�E��T0 k� ��V��Ve2D# 3I)@5   ��    � <�xQ0�bpN����Lh!� 	��u��c3�1�7EC�E��T0 k� ��T��Te2D# 3I)@5   ��    � <�vQ0�b�O����Lh!� 	��u��b3�1�7EG�E��T0 k� ��S��Se2D# 3I)@5   ��    � <�tQ0�c�R��!�� h� 	.�t��_3�1�7ES�E�T0 k� ��P��Pe2D# 3I)@5   ��    � <�rQ0�c�S�"�� h� 	.�tμ]3�1�6EW�E�T0 k� ��N��Ne2D# 3I)@5   ��    � <�pQ0�c�U�$��  h� 	.�tθ\3�1�6E[�E�T0 k� ��M��Me2D# 3I)@5   ��    � <�nQ0�c�V�&�� h� 	.�tΰZ3�1�6E_�E�T0 k� ��K��Ke2D# 3I)@5   ��    � <�lQ0�c�X�(�� h� 	.�tάY3���6Ec�E��T0 k� �xJ�|Je2D# 3I)@5   ��    � <�jQ0�c�Y�)�� h� 	�tΨW3���6Eg�E��T0 k� �tH�xHe2D# 3I)@5   ��    � <�hQ0�c�Z�+�� h� 	�tΠU3���5Eok�E��T0 k� �pF�tFe2D# 3I)@5   �    � <�hQ0�c�[�-�� lh� 	�tޜT3���5Eoo�E��T0 k� �dD�hDe2D# 3I)@5   �    � <�hQ0�cP]�.�� lh� 	�tޔR3���5Eos�E�#�T0 k� �\A�`Ae2D# 3I)@5   ��    � <�hQ0�cP^�0�� lh� 	�tސQ3���5Eow�E�'�T0 k� �T@�X@e2D# 3I)@5   ��    � <�hQ0�cP_��1�#� lh� 	 �sތO3���5Eo{�E�+�T0 k� �P>�T>e2D# 3I)@5   ��    � <�hQ0�cP`��3�'� lh� 	 �sބN3���5Eo�E�/�T0 k� �L<�P<e2D# 3I)@5   ��    � <�hQ0�cPb��5�+��l� 	 �sހL3���5Eo��E�/�T0 k� �D;�H;e2D# 3I)@5   ��   � <�hQ0�c@c��6�/��l� 	 �s�xJ3�� 5Eo��E�3�T0 k� �@9�D9e2D# 3I)@5   ��    � <�hQ0�c@d�x8�3��l� 	 �s�tI3� 5Eo��BB7�T0 k� �88�<8e2D# 3I)@5   ��    � <�hQ0�c@e�t9�7��l� 	 �s�pG3�5Eo��BB;�T0 k� �46�86e2D# 3I)@5   ��    � <�hQ0�c@g�l:�;��p� 	 �s�hF3�5A���BB?�T0 k� �,5�05e2D# 3I)@5   ��    � <�hQ0�c@h�d<M?��p� 	 �s�dD3�5A���BB?�T0 k� �(3�,3e2D# 3I)@5   ��    � <�hQ0�c@i�`=MC��t� 	 �s�\C3�4A���BBC�T0 k� �$1�(1e2D# 3I)@5   ��    � <�hQ0�c@k�X?MG��t� 	 �s�XA3�4A���BBG�T0 k� �0� 0e2D# 3I)@5   ��    � <�hQ0�c@l�P@MK�x� 	 �s�T?3�4A���BBK�T0 k� �.�.e2D# 3I)@5   ��    � <�hQ0�c@ nLAMO�x� 	 �s�L>3�4A���BBK�T0 k� �-�-e2D# 3I)@5   ��    � <�hQ0�c@ oDC�S�|� 	 �s�H<3�4A���BBO�T0 k� �+�+e2D# 3I)@5   ��    � <�hQ0�cO�p<D�W�|� 	 �s^@;3�4A���BBS�T0 k� �/�/e2D# 3I)@5   ��G    � <�hQ0�c��r4E�[��� 	 �s^<93�4A���BBW�T0 k� �3�3e2D# 3I)@5   ��G    � <�hQ@�c��s,F�_���� 	 �s^483�4A���BBW�T0 k� �5�5e2D# 3I)@5   ��G    � <�hQ@�c��u(H�c���� 	 �s^063� 4A���BB[�T0 k� �6�6e2D# 3I)@5   ��G    � <�hQ@�c��v I�g���� 	 �r^(53� 4A���BB_�T0 k� �7�7e2D# 3I)@5   ��G    � <�hQ@�c��xJ�k���� 	 �r^$43�$4A���BB_�T0 k� � 7�7e2D# 3I)@5   ��G    � <�hQ@�c��yK�k���� 	 �r^23�(4A���BBc�T0 k� ��7� 7e2D# 3I)@5   ��G    � <�hQ@�c��zL�o���� 	 �r^13�(4A���BBg�T0 k� ��6��6e2D# 3I)@5   ��G    � <�hQ@�c��| M�s���� 	  r^03�,4A�íBBg�T0 k� ��6��6e2D# 3I)@5   ��G    � <�hQ@�c��}�N�w���� 	  rN.3�,3A�ǮBBk�T0 k� ��7��7e2D# 3I)@5   ��G    � <�hQ@�c���P�{���� 	 rN -3�03A�ǯBBk�T0 k� ��7��7e2D# 3I)@5   ��G    � <�hU�c�܀�Q�{���� 	 rM�,3�03A�˯BBo�T0 k� ��8��8e2D# 3I)@5   ��G    � <�hU�c�؀�R����� 	 rM�+3�43A�ϰBBs�T0 k� ��8��8e2D# 3I)@5   ��G    � <�hU�c���S����� 	 rM�*3�43A�ϰBBs�T0 k� ��8��8e2D# 3I)@5   ��G    � <�hU�c���T����� 	 rM�)3�83A�ӱBBw�T0 k� ��8��8e2D# 3I)@5   ��G    � <�hU c���U����� 	 rM�(3�83A�ײBBw�T0 k� ��7��7e2D# 3I)@5   ��G    � <�hU c��~�V��ܬ!� 	 rM�'3�<3A�ײBB{�T0 k� ��6��6e2D# 3I)@5   ��G    � <�hUc��~�W��ܰ"� 	 rM�&3�<3A�۳BB{�T0 k� ��6��6e2D# 3I)@5   ��G    � <�hUc�~�X��ܰ#� 	 rM�&3�@3A�߳BB�T0 k� ��5��5e2D# 3I)@5   ��G    � <�hUc�}�Y��ܴ$� 	 r�%3�@3A�ߴBB�T0 k� ��4��4e2D# 3I)@5   ��G    � <�hUc�}�Z��ܸ%� 	 r�$3�@3A��BB��T0 k� ��4��4e2D# 3I)@5   ��G    � <�hUc�}�[��ܸ'� 	 r�$3�D3A��BB��T0 k� ��3��3e2D# 3I)@5   ��G    � <�hUc�}�[��ܼ(� 	 r�#3�D3A��BB��T0 k� �t3�x3e2D# 3I)@5   ��G    � <�hUc��|�\��ܼ)� 	 r�#3�H3A��BB��T0 k� �l2�p2e2D# 3I)@5   ��G    � <�hUc��|�]����*� 	 r�#3�H3A��BB��T0 k� �d2�h2e2D# 3I)@5   ��G    � <�hUc��|�x^����+� 	 r�"3�L3A��BB��T0 k� �\1�`1e2D# 3I)@5   ��G    � <�hUc��|�p_����,� 	 r�"3�L3A��BB��T0 k� �T1�X1e2D# 3I)@5   ��G    � <�hUc��{�h`����-� 	 q�"3�L3A��BB��T0 k� �L1�P1e2D# 3I)@5   ��G    � <�hUc��{�`a����.� 	 q�|!3�P2A��BB��T0 k� �H,�L,e2D# 3I)@5   ��G    � <�hUc�|{�Xa����/� 	 q�t!3�P2A���BB��T0 k� �D(�H(e2D# 3I)@5   ��G    � <�hUc�t{�Pb����0� 	  q�l!3�T2A���BB��T0 k� �@%�D%e2D# 3I)@5   ��G    � <�hUc�lz�Hc����1� 	  q�d!3�T2A���BB��T0 k� �<#�@#e2D# 3I)@5   ��G    � <�hUc�dz�@d����2� 	  q�\!3�T2A���BB��T0 k� �4"�8"e2D# 3I)@5   ��G    � <�h@ac�`z�8e����3� 	 $q�T 3�X2A���BB��T0 k� �,!�0!e2D# 3I)@5   ��G    � <�h@ac`z�0e����4� 	  q�H 3�X2A���BB��T0 k� �$�(e2D# 3I)@5   ��G    � <�h@ac\z�(f����5� 	  p�@ 3�X2A��BB��T0 k� ��e2D# 3I)@5   ��G    � <�h@acXz�g����6� 	 p�8 3�\2A��BB��T0 k� ��e2D# 3I)@5   ��G    � <�h@acTz�g����7� 	 o�0 3�\2A��BB��T0 k� ��e2D# 3I)@5   ��G    � <�h@�cL{�h�����8� 	 o�(3�\2A��BB��T0 k� ��� e2D# 3I)@5   ��G    � <�h@�cH{�i�����9� 	 n� 3�`2A��BB��T0 k� ����e2D# 3I)@5   ��G    � <�h@�cD{��j�����9� 	 n�3�`2A��BB��T0 k� �� �� e2D# 3I)@5   ��G    � <�h@�c@|��j�����:� 	 m�3�`2A��BB��T0 k� ��!��!e2D# 3I)@5   ��G    � <�h@�c8|��k�����;� 	 m�3�d2A��BB��T0 k� ��"��"e2D# 3I)@5   ��G    � <�hAc4|��k�����<� 	 l� 3�d2A��BB��T0 k� �� �� e2D# 3I)@5   �G    � <�hAc0|��l�����=� 	 l��3�d2A��BB��T0 k� ����e2D# 3I)@5  ��O    � <�hAc(}��l�����>� 	 k��3�h2A��BB��T0 k� ����e2D# 3I)@5  ��O    � <�hAc$}��m�����>� 	 k��3�h2A��BB��T0 k� ����e2D# 3I)@5  ��O    � <�hAc}��m�����?� 	 j��3�h2A��BB��T0 k� ����e2D# 3I)@5  ��O    � <�hC�c}�n�����@� 	 j��3�l2A��BB��T0 k� ����e2D# 3I)@5  ��O    � <�hC�c~�n�����A� 	 j��3�l2A��BB��T0 k� ����e2D# 3I)@5  ��O    � <�hC�c�~�n�����A� 	 i��3�l2A��BB��T0 k� ����e2D# 3I)@5  ��O    � <�hC�c�~�n�����B� 	 i��3�l2A��BB��T0 k� ����e2D# 3I)@5  ��O    � <�hC�c��~�n�����C� 	 h��3�p2A��BB��T0 k� �|��e2D# 3I)@5  ��O    � <�hC�c����n�����C� 	 h�3�p2A��BB� T0 k� �p�te2D# 3I)@5  ��O    � <�hC�c����n�����D� 	  g�3�p2A��BB� T0 k� �h�le2D# 3I)@5  ��O    � <�hC�c���|n�����E� 	  g�3�p2A�#�BB� T0 k� �`	�d	e2D# 3I)@5  ��O    � <�hC�c���tn�����F� 	  g�3�t2A�#�BB� T0 k� �T�Xe2D# 3I)@5  ��O    � <�hC� c���lnM��� F� 	 �f�3�t1A�#�BB� T0 k� �L�Pe2D# 3I)@5  $�O    � <�hC��c�Ԁ�dnM��� G� 	 �f�3�t1A�'�BB�T0 k� �P�Te2D# 3I)@5  ��O    � <�hC��c���\nM��� G� 	 �f�3�t1A�'�BB�T0 k� �P�Te2D# 3I)@5  ��O    � <�hC��c���TmM���H� 	 �e�3�x1A�'�BB�T0 k� �T�Xe2D# 3I)@5  ��O    � <�hC��c��LmM���I� 	 �e�3�x1A�+�BB�T0 k� �X�\e2D# 3I)@5  ��O    � <�hC��c�~�DmM���I� 	 �e�3�x1A�+�BB�T0 k� �\�`e2D# 3I)@5  ��O    � <�hC��c�~�<lM���J� 	 �d�|3�x1A�+�BB�T0 k� �`�de2D# 3I)@5  ��O    � <�hC��c>�~4lM���K� 	 �d�x3�|1A�/�BB�T0 k� �`�de2D# 3I)@5  ��O    � <�hC��c>�}0kM���K� 	 �d\t3�|1A�/�BB�T0 k� �d�he2D# 3I)@5  ��O    � <�hC��c>�}(jM���L� 	 �c\l3�|1A�/�BB�T0 k� �h�le2D# 3I)@5  ��O    � <�hC��c>�} jM���L� 	 �c\h3�|1A�3�BB�T0 k� �l�pe2D# 3I)@5  ��O    � <�hC��c>�|iM���M� 	 �c\d3�|1A�3�BB�T0 k� �l�pe2D# 3I)@5  ��O    � <�hC��c>�|i]���M� 	 �b\\3��1A�3�BB�T0 k� �p�te2D# 3I)@5  ��O    � <�hD �c>||h]���N� 	 �b\X3��1A�3�BB�T0 k� �t�xe2D# 3I)@5  ��O    � <�hD �c>x{g]���N� 	 �b\T3��1A�7�BB�T0 k� �x�|e2D# 3I)@5  ��O    � <�hD �c>p{f]���O� 	 �a\P3��1A�7�BB�T0 k� �|��e2D# 3I)@5  ��O    � <�hD �c>h{ e]���O� 	 �a\L3��1A�7�BB�T0 k� �|��e2D# 3I)@5  ��O    � <�hD �c>dz�e]���P� 	 �a\D3��1A�7�BB�T0 k� ����e2D# 3I)@5  ��O    � <�hL�c>\z��d]���P� 	 �`\@3��1A�;�BB�T0 k� �� �� e2D# 3I)@5   ��O   � <�hL�c>Xz��c]���Q� 	 �`\<3��1A�;�BB�T0 k� �� �� e2D# 3I)@5   ��O    � <�hL�cNPz��b]�� �Q� 	 �`\83��1A�;�BB�T0 k� �� �� e2D# 3I)@5   .�O    � <�hL�cNLy��a]�� �R� 	 �`\43��1A�;�BB�T0 k� �� �� e2D# 3I)@5   ��O    � <�hL�cNDy��a]�� �R� 	 �_\03��1A�?�BB�T0 k� �����e2D# 3I)@5   ��O    � <�hL�cN@y��`m�� �S� 	 �_\,3��1A�?�BB�T0 k� �����e2D# 3I)@5   ��O    � <�hL|cN<y��_n� �S� 	 �_\(3��1A�?�BB�T0 k� �����e2D# 3I)@5   ��O    � <�hLtcN4x��^n� �T� 	 �_\$3��1A�?�BB�T0 k� �����e2D# 3I)@5   ��O    � <�hLlcN0x��^n� �T� 	 �^\ 3��1A�C�BB�T0 k� �����e2D# 3I)@5  ��O    � <�hLhcN,x��]n� � U� 	 �^\3��1A�C�BB�T0 k� ܣ����e2D# 3I)@5  ��O    � <�hL`cN$w��\n� � U� 	 �^\3��1A�C�BB�T0 k� ܧ����e2D# 3I)@5  ��O    � <�hLXcN w��\n� � U� 	 �^\3��1A�C�BB�T0 k� ܧ����e2D# 3I)@5  ��O    � <�hL TcNw��[n� � V� 	 �]\3��1A�C�BB�T0 k� ܫ����e2D# 3I)@5  ��O    � <�hL LcNw��Zn� �$V� 	 �]\3��1A�G�BB�T0 k� ܯ����e2D# 3I)@5  ��O    � <�hL DcNw��Zn� �$W� 	 �]\3��1A�G�BB�T0 k� �����e2D# 3I)@5  ��O    � <�hL @cNv��Yn� �$W� 	 �]\3��1A�G�BB�T0 k� �����e2D# 3I)@5  ��O    � <�hL 8cNv��X~� �$W� 	 �]\3��1A�G�BB�T0 k� �����e2D# 3I)@5   ��O    � <�hL 4cNv��X~� �$X� 	 �\\ 3��1A�G�BB�T0 k� �����e2D# 3I)@5   ��O    � <�hL ,cM�v��W~� �(X� 	 �\\ 3��1A�K�BB�T0 k� �����e2D# 3I)@5   ��O    � <�hL $cM�u��W~� �(Y� 	 �\[�3��1A�K�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL  cM�u��V~� �(Y� 	 �\[�3��1A�K�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL cM�u��U~ �(Y� 	 �[[�3��1A�K�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL cM�u��U~ �(Z� 	 �[[�3��1A�K�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL cM�u��T~ �,Z� 	 �[[�3��1A�O�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL cM�t��T~ �,Z� 	 �[[� 3��1A�O�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL  cM�t��S~ �,[� 	 �[[� 3��1A�O�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�t��S~	 �,[� 	 �[[� 3��1A�O�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�t��RN �,[� 	 �Z[�!3��1A�O�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�t��RN �0\� 	 �Z[�!3��1A�O�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�s��QN �0\� 	 �Z[�!3��1A�S�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�s��QN �0\� 	 �Z[�!3��1A�S�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�s��PN �0]� 	 �Z[�"3��1A�S�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�s��P��0]� 	 �Y[�"3��1A�S�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�s��O��0]� 	 �Y[�"3��1A�S�BB�T0 k� ������e2D# 3I)@5   ��O   � <�hL/�cM�s��O��4^� 	 �Y[�#3��1A�S�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�r��N��4^� 	 �Y[�#3��1A�W�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�r��N��4^� 	 �Y[�#3��1A�W�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�r��M��4^� 	 �Y[�#3��1A�W�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�r��M�!�4_� 	 �Y[�$3��1A�W�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�r��L�#�4_� 	 �X[�$3��1A�W�BB�T0 k� ������e2D# 3I)@5   ��O    � <�hL/�cM�r��L�%�4_� 	 �X[�$3��1A�W�BB�T0 k� �����e2D# 3I)@5   ��O    � <�hL/�cM�q��K�'�8`� 	 �X[�$3��1A�W�BB�T0 k� ����e2D# 3I)@5   ��O    � <�hL/�cM�q��K�)�8`� 	 �X[�%3��1A�[�BB�	T0 k� ����e2D# 3I)@5   ��O    � <�hL/�c=�q��K�+�8`� 	 �X[�%3��1A�[�BB�	T0 k� ����e2D# 3I)@5   ��O    � <�hL/�c=�q��J�-�8`� 	 �X[�%3��1A�[�BB�	T0 k� ����e2D# 3I)@5   ��O    � <�hL/�c=�q��J�/�8a� 	 �X[�%3��1A�[�BB�	T0 k� ����e2D# 3I)@5   ��O    � <�hL/|c=�q��I�1�8a� 	 �W[�&3��1A�[�BB�	T0 k� ����e2D# 3I)@5   ��O    � <�hL/xc=�q��I�3�8a� 	 �W[�&3��1A�[�BB�	T0 k� ����e2D# 3I)@5   ��O    � <�hL/pc=�p��I�5�<a� 	 �W[�&3��1A�[�BB�	T0 k� ����e2D# 3I)@5   ��O    � <�hL/hc=�p��H�7�<a� 	 �W[�&3��1A�[�BB�	T0 k� ����e2D# 3I)@5   ��O    � <�hL/dc=�p��H�9�<b� 	 �W[�'3��1A�_�BB�	T0 k� ����e2D# 3I)@5   ��O    � <�hL/\c=�p��H�;�<b� 	 �W[�'3��1A�_�BB�	T0 k� ���#�e2D# 3I)@5   ��O    � <�hL/Xc=�p��G�=�<b� 	 �W[�'3��1A�_�BB�	T0 k� �#��'�e2D# 3I)@5   ��O    � <�hLPc=�o��G�?�<b� 	 �W[�'3��1A�_�BB�	T0 k� �'��+�e2D# 3I)@5   ��O    � <�hLDc=xo��F�C�<c� 	 �V[�(3��1A�_�BB�
T0 k� �+��/�e2D# 3I)@5   ��O    � <�hL@c=xn��F�E�@c� 	 �V[�(3��1A�_�BB�
T0 k� �/��3�e2D# 3I)@5   ��O    � <�hL8c=tn��E�G�@c� 	 �V[�(3��1A�_�BB�
T0 k� �3��7�e2D# 3I)@5   ��O    � <�hL4c=tn��E�I�<c� 	 �V[�(3��1A�_�BB�
T0 k� �3��7�e2D# 3I)@5   ��O    � <�hC�,c=po��E�J�<c� 	 �V[�(3��1A�c�BB�
T0 k� �7��;�e2D# 3I)@5   ��O    � <�hC�(c=po��E�L�<c� 	 �V[�)3��1A�c�BB�
T0 k� �;��?�e2D# 3I)@5   ��O    � <�hC� c=po��D�N�<c� 	 �V[�)3��1A�c�BB�
T0 k� �;��?�e2D# 3I)@5   ��O    � <�hC�c=lo��D�P�8c� 	 �V[�)3��1A�c�BB�
T0 k� �?��C�e2D# 3I)@5   ��O    � <�hC�c=lo��D�R�8c� 	 �U[�)3��1A�c�BB�
T0 k� �C��G�e2D# 3I)@5   ��O    � <�hC�c=lo��C�S�8c� 	 �U[�)3��1A�c�BB�
T0 k� �G��K�e2D# 3I)@5   ��O    � <�hC�c=ho��C�U�8b� 	 �U[�)3��1A�c�BB�
T0 k� �G��K�e2D# 3I)@5   ��O    � <�hC��c=ho��C�W�4b� 	 �U[�*3��1A�c�BB�
T0 k� �K��O�e2D# 3I)@5   ��O    � <�hC��c=ho��B�X�4b� 	 �U[�*3��1A�c�BB�
T0 k� �O��S�e2D# 3I)@5   ��O    � <�hC��c=do��B�Z�4b� 	 �U[�*3��1A�c�BB�
T0 k� �O��S�e2D# 3I)@5   ��O   � <�hC��c=do��B�\�4b� 	 �U[�*3��1A�g�BB�
T0 k� �S��W�e2D# 3I)@5   ��O    � <�hC��cMdo��B]�4b� 	 �T[�*3��1A�g�BB�T0 k� �W��[�e2D# 3I)@5   ��O    � <�hC��cM`o��A_�0b� 	 �T[�*3��1A�g�BB�T0 k� �W��[�e2D# 3I)@5   ��O    � <�hC��dM`o��A`�0b� 	 �S[�+3��1A�g�BB�T0 k� �[��_�e2D# 3I)@5   ��O   � <�hC��dM`o��Ab�0b� 	 �S[�+3��1A�g�BB�T0 k� �_��c�e2D# 3I)@5   ��O    � <�hC��eM\o��Ac�0b� 	 �R[�+3��1A�g�BB�T0 k� �_��c�e2D# 3I)@5   ��O    � <�hC��eM\o��@e�0a� 	 �R[�+3��1A�g�BB�T0 k� �c��g�e2D# 3I)@5   ��O    � <�hC��eM\o��@ f�,a� 	 �R[�+3��1A�g�BB�T0 k� �g��k�e2D# 3I)@5   ��O    � <�hC��fM\o��@ h�,a� 	 �Q[�+3��1A�g�BB�T0 k� �k��o�e2D# 3I)@5   ��O    � <�hE^�fMXo��@ i�,a� 	 �Q[�,3��1A�g�BB�T0 k� �k��o�e2D# 3I)@5   ��O    � <�hE^�gMXo��? j�,a� 	 �P[�,3��1A�g�BB�T0 k� �o��s�e2D# 3I)@5   ��O    � <�h                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��
V ]�(6(5 � �� o�  � �     ��g!     of��iS�    S޺             ,
 Z�h           <��  &  ��� 
	           o��   � �	    ��P?@     o�)�PlW     8�Y            Z�h         ��    ���   0
&          =H0   / /      �B�U     =f�Ar/    �i          #  Z�h         0�     ���   8	          }�   � �    �|L�     ~-��|j(    ���D            8 Z�h          %��    ���  84          _�       .�G�     _���G!-    �H�4               0 Z�h          ��     ���   8
	
 
          	6�  ��     B�z�     	6��z�           
                   �o             !  ���     

 0             H�Y           V��5�     H�`��W�    �i��                  �          ��      ��@   0           /u    
	  j����     /\����3    n                 ��          ��     ��H    		�           Y� ��      ~ ��c     Y� ��c                           ����        ,`      ��@    0)           1   S	     � ��     1 ���       �               	 A �         	 `     ��@   H


         ��u�        � �    ��i1 �     � �                  d 5        
 �  �  ��@   8           �^ $ O     � ��V     � ���     � �                
 	   �         v�     ��@   P

 		                ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��1  ��        ��n,�  C�����m�I  C���	�                  x                j  �   �   �                         ��    ��        ��o      ��  �n           "                                                �                         �g�P�B�|�G����� � �  ����n�o    	   
          
  �   � �k ��n       �� �[� ¤ 0\� � ]  �$ ]@ �� 0\� �D  ]@ �� ]� � d� �$ d� E�  d@��� ����  ����. ����< ����J ����X � 
�| W� 
�\ W� �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ � }`���� � 
�| V ���� ����� � �� �^@ �� _@ �$ `y� ��  z� ބ �c@ �$ }@ ��  }` ��  }����� � � }` gD `j� h k� h$ 0k� 3� �c@ 4� d@ *d �^@ +d _@ +� _` 
�\ W� 
�| W� 
�| W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����h�� <�� �  ������  
�fD
��L���"����D" � j  "  B   J jF�"     
�j � � 
��
��
��"   "D�j�
�� " �
� �  �  
�      ��     ��@  �    _    ��     ��G       /    ��     ���          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �O� �      ��3 �  ���        � �T ��        �        ��        �        ��        �    ��     ������        ��                         ��  0 $� ���                                     �                ����            	����%��   <�h��       !         19 John Cullen  y  k   1:26                                                                        3  3      �C
� �Tcj �t cr �J� �J� �2 CB �:CC �R CI �:	CJ �
C � � C �C.  C60 �B�-
 B�3 �B�& �B�. � B�6 �J�- �J�5 � J�/ � J�% � � � � � � �C8 �C"8 � C%> � C&H �cV"� "�) "�!*�"t""� �t #"� �d$� �d%
� � p &*Gt0 '*IdH (*OdH *(lH **OdH *(l ,*,t0 -*DdH .*RdP  *l`0*
l` *6tH2*2t`3*
l` *6t` *6tH6*2t` *6t@8*<dH9*2t` *6t � ;*~ �  *Kv � =*~ �  *Kv �  *Hv                                                                                                                                                                                                                         �� P         �    @         1     X P E _  ���� 
               �������������������������������������� ���������	�
��������                                                                                          ��    ��� 
  ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, 1� 0 a����@�@p���@����@�@������                                                                                                                                                                                                                                                                                                                         )A��x"���                                                                                                                                                                                                                                     �  
  .     ��  :�J      �                             ������������������������������������������������������                                                                                                                             
         c   �                  �  �                  
     ��������� ������� ������� ���������� ��������   ������ � ��������� ��������� ���������������������� ������� �������� �������������� �����������  ������������������� �������� ������ ���������������� ������ ������ �� �           �                �  	  #    ��  E�J      4�  	                           ������������������������������������������������������                                                                                                                                            g    ��              �         � �    �        
 	    �� ������������ �������� ��� �� ������������ ����� �������������������������� ��������������������������������������������������������� �� � ����� ����� ������� ���  ���������������� ���� ���� ��� ������������             �                                                                                                                                                                                                                             	                                                                               �             


             �  }�    �               '�                                     Rx     'v                        ����������������    ����������������������������   ������������������������������������  + ������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" R > / 	                                � ���� �[�                                                                                                                                                                                                                                                                                      )n)n�  	n              l                                    m                                                                                                                                                                                                                                                                                                                                                                                j             j          > �  >�  
(~    j  (~  EZm6  �N ~�����;����(��������� ���d���������8��          0   }�F :�� H        ��   & AG� f ��              lt�                                                                                                                                                                                                                                                                                                                                     K H   �                     !��                                                                                                                                                                                                                            Y   �� �~ ���      �� 7  �� 
��������� ������� ������� ���������� ��������   ������ � ��������� ��������� ���������������������� ������� �������� �������������� �����������  ������������������� �������� ������ ���������������� ������ ������ �� ��� ������������ �������� ��� �� ������������ ����� �������������������������� ��������������������������������������������������������� �� � ����� ����� ������� ���  ���������������� ���� ���� ��� ������������    ��      $��˪����ɻ���������˪������������ʻ������ɻ����������������ƪ��f��˫�������f��fƦfffffffffffffff˪������f����fflffffffffffffffffʚʫ������������i���l���fʪ�fj���˺j����˪��������˻�����������������������������������ʹ����������f���f��ff��ff��ff��ff�fff�fffffffffffffffffffffffff�flffffff�fffffffffffffffffffff�ff���f����fj��ff��ffʪffj�ffj�fff�fff�fff��ʻ̼̪����˻���ʻ�����ʻ��������������������������������ʛ����ʺffl�ffl�ffɫff��ff��ff��fk��fi�fl���ʼ��ʧw�UWU�UUU�f�U���UuW���������xy���UUWwUuxxX�f̩̊���Uy�ffʜffi�ffk�ffj�ffk��fjȶfj��f�������������������ʪ�������������ʺ������������������������������fi���i���Ɉ�������������h����z��gʘ�����X��Ux��wW�uUX��uz���xZw���ʫ�����w��xwx��wx��wX˹x��xw���f���i���y�����������������������ʻ������ʺ�������ˬʺ�����ʻ����ʙ����������������������������������j���l����������������������x����y����w����������w���w���wx��x�����|�������������������w�����̺��j��fk��ff���i��f���ɺ˙���ʛ�����˫ʺ����������������ʻ�������������������wuUZUUUVUUUVUUUV�������������fi�feU�kUY�eU�weU�X���u�������̇��̉������U���w�xyy��������ʻ���ʘ������������wx�uw�ɺ�����������|f��U����Ux�eUx��U����������ʺ����j���feW�fUUUkUUU8      F   &   4   #����                       7     �   �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f          p����        5� � ��    �@���6      � �N ^$ �@  �@  �@   �  �     �    ����� ��   ����� �$ ^$��   �  �� | 
p � �&      $   # [� �� �� [� �� �$   ��#       �  ��   ���� e����J   g���        f ^�         �� <            ��
��������J���J��e���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                               	                 �  ��� �UU���U              �	���UUU�UUUUUU      	� ��U�UUUUUUUUUUUUUUUUUUU    ��� U^��UUU�UUU^UUUUUUUUUUUU            �   �   ^�  U�  UY�    � 	UU 	��  	�  	�  �^ 	��    �	UY�������UUUUUUU��UU��UU�U�UUUUUUUUUUUUUUUUUUUUUUUUUUUU^UUUYUU^�U^� U� ^�  �  ��  �   �   ��UU ��U �U  �U  ��            U^� UU� UU� UU� ���                    	   �       	   	   	    �UUU�UU���U  	�� �����U�UUU�UUUUUUYUUUYUUUYUUU^UUU^UUUUUUUUUUUU�   �   �   �   �   � �^���U^��            	����UUU�UUU�UUUUUU^            ��  U�  Y�  �  �      �   �   �   	                ���Y���U��Y�^�U��U ��^ 	� 	� UUUU�UUUUUUUU^�U^����� �        UUUUUUUUUUUUUUUUUUUU�������    UUU�UU^�UU�U� Y�  ��          �                               wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "! " ""  "!  " ! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ "!    " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "! " ""  "!  " ! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        "  " �" ��" ��- �ۼ w۽��ݹ����� ��� ��  ˼  ��  ˼  ��  H�  �D  J�  J�  �  �  �  �  
�  �  �  �  ,�  " "" �" �"�   ˰  ��  wp ��ډ�v���r�̸��˰��� ��  ��  ��  ��  ̸  ��  ��  DC  C4@ T4@ T40 T30 T30 S;� H�  ��  ��  ��  ""  "  �""� "�/��        �   �   �      �  �   �   �   �   �              �   �   �   �             ���� �                        " "" """ �"  �   �   �                              � ��                  �  �˰ ��� �wp ���                                                                                                                                                                   �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �               ���                            ���������������������  ��  ��  ��  �   �    �          �         �                                                                                                     �   �  �  �  	�  �  EH  ET DU CE DD4 DD3 DC0 �3 ɰ �  ,�  +�  "/  ������ � ̹�p�˚��̹���ː�̼�̻���ۜ��۩�ݍ���=��J�ܰT�� EJ�0 EJ� I�  ��  �"  ""  "/  "�� ���                    ̰ ̻ ̻	���̚�w          �.���       �  �      �  ��  �  ��  �            �  �   �   ��  �             ��  ��  �                            �   �    �   �       �   �   �                .                  �   �               �  ��� ݼ� w{� �װ vw�                    �   ���                            �   �                                                                                                   "  " �" ��" ��- �ۼ w۽��ݹ����� ��� ��  ˼  ��  ˼  ��  H�  �D  J�  J�  �  �  �  �  
�  �  �  �  ,�  " "" �" �"�   ˰  ��  wp ��ډ�v���r�̸��˰��� ��  ��  ��  ��  ̸  ��  ��  DC  C4@ T4@ T40 T30 T30 S;� H�  ��  ��  ��  ""  "  �""� "�/��        �   �   �      �  �   �   �   �   �              �   �   �   �             ���� �                        " "" """ �"  �   �   �                              � ��                  �  �˰ ��� �wp ���                                                                                                                                                                               �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                /���"/�  ��                    �                                                                            �               �  �  ��  �   �   �           �     �                                                                                                                                                                                                    �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �          �  � � �� ��     �   �������  �                     �  �   �  �  ��  �  ��  �                                                                                                                                                                                                     �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �   �   �   ˰  ˙  ɪ  ��� ټ� �̰ �̰ ��� ��  ��                              ��                     �   �                      �������  ���    �                    �   ���       ���� �                                                                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                    ""  ."  �"    �   ��  �   �                  �  �  �  �                                       �  �   ��                     �    � �  ��                  ���                     �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                           �� �����ݼڜ��ک��ک��z�	��� 
�� 
�� 	�� ̘ ɪ  ��  �  �� �� ������������ ���  � � � �� �� ������ ��                      �   ��  ��  �̰ ��� ��˰�̻��̻���������ˉ�U��EP�ET �I� ٕ  �D� �L� ��� ��" ����/�"�"�""�����                         U   T           �  �       �           �   /�  /   �  �                   �   �        �           �   �  �  �   �               �   �                     �                                                                                                                                                                                          	�  �� �� ���ܙܽɪ�͚�����͙ͼ̨��̄DC"�D32�C33�333�33P330X̽ 
�� ˪  "   ""/"""�����vv ��p ��  ��  ̽  ˸  ɚ  ��  ؛  -�� .ܰ .��  �"  �   .   "�                   � �  ��            Z   Z   Z   Z  Z  �� �� �� "� "" "" ""/ ����   �   � ���� �� ����                    �� ��������p��}`                            ��          �  ��� ̻� ��� rbp wgz�               �������  ���    �        � ��                    ���� �                                                   ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                    �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    �  �   �  �     �                                       ��                     �   �                      �������  ���    �                    ��  ��  ���                    � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        �� wڪ z�� ���
���	������
���̪��̹����ӈ��E �U ��U�UD�D 
��  ��  ˰ ",� """��"" ��  �    �   �   ��  ̨  ̋  �۰ �۰ ��� �=  30  DC  UD0 T4J 3DT�4U@ 3D� ;�  �   �   ��  ��  �   �   �   ""  �"  � ��� �                      ̰ ̻ ��                               �   �   ��  � " ��"  "                                    ��  "   "   "  �� ��                   ����������                                ��  ��  ���  �  �  �   �   ��  �                            �   ���                            �   �                                                                                                               �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""��������������������""""������DDM�D��""""�������MM�M�M""""��������DD�A��""""�������MAA�MA""""��������AA�A""""����������M�MA""""������������M���M���M���"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUQUUQUUUUUUQUUUUUUUU3333DDDDUUUUDEEDDTEUUUU3333DDDDAEAEQQUDTDUUUU3333DDDDQUQUQDUDDUUUU3333DDDDAADAUAUEDUTUUUU3333DDDDADAEAQAUEDUTUUUU3333DDDDUDUQEUQUUQUEUDUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""������������������""""������������������������""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""���������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��������������D�����3333DDDDI����D��DI����3333DDDDADAIA����D������3333DDDD��������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=LL����������D����3333DDDD    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����������A������ x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx""""�������I�I������ w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww""""�������I��D���I�������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(�D�M�D���M������3333DDDD �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""�����AMAD������ M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M""""������������������ � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�fFfFDfFFfFffdFffff3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DDFFDfFFfdFffff3333DDDD 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5""""wwwwwwwGGD x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x""""wwwwwwqwAqwAwA w w x y�������H���������������������������������H������yxww""""wwwwqwqAwAqAqAq  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(A�A�A�A��LD�����3333DDDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,�A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
� �Tcj �t cr �J� �J� �2 CB �:CC �R CI �:	CJ �
C � � C �C.  C60 �B�-
 B�3 �B�& �B�. � B�6 �J�- �J�5 � J�/ � J�% � � � � � � �C8 �C"8 � C%> � C&H �cV"� "�) "�!*�"t""� �t #"� �d$� �d%
� � p &*Gt0 '*IdH (*OdH *(lH **OdH *(l ,*,t0 -*DdH .*RdP  *l`0*
l` *6tH2*2t`3*
l` *6t` *6tH6*2t` *6t@8*<dH9*2t` *6t � ;*~ �  *Kv � =*~ �  *Kv �  *Hv3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������=�N�K�U�X�K�T��0�R�K�[�X�_� � � � � � �-�1�B�������������������������������������������1�G�X�_��;�U�H�K�X�Z�Y� � � � � � � � �-�1�B�����������������������������������������$��4�U�N�T��-�[�R�R�K�T� � � � � � � � � �=��;�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������=��;� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�1�B� �� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            