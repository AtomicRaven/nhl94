GST@�                                                            \     �                                                ��      �  ��  �         ����e ����J�����������x�������        f      #    ����                                d8<n    �  ?     p�����  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    B�jl �   B ��
  l�                                                                              ����������������������������������      ��    bbo QQ g 11 44               		� 

                      ��                      nn� ))         888�����������������������������������������������������������������������������������������������������������������������������o=  0  o4   1  +      '           �                    	�  7�  V�  	�                  E            : �����������������������������������������������������������������������������                                ��  �       M�   @  #   �   �                          �                                                     '     )n)n�  E    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    �*  E�0?b�40r|,�өA P`$ ��/��Zc`T0 k� �%�%��d  e1�t B  ��H    �  ��+  E�0@b�40r|,�өA  P\$ ��/��Zc`T0 k� �%�%��d  e1�t B  ��H    �  ��,  E�,Ar� �0r|,�ϩA  P\% ��/��Zc`T0 k� �%�%��d  e1�t B  ��H    �  ��-  E�,Ar� �0r|,�ϩA  PX% ��/��Zc`T0 k� �&�&��d  e1�t B  ��H    �  ��.  LQ,Br� �0r|,�ϩA�PX% ��/��Zc`T0 k� �&�&��d  e1�t B  ��H    �  ��0  LQ(Cr� �4r|,�ϩA�PX% ��/��Zc\T0 k� �&�&��d  e1�t B  ��H    �  ��1  LQ(Cr� �4r|,�ϩA�PT& ��/��Zc\T0 k� �&�&��d  e1�t B  ��H    �  ��2  LQ$Dr� �4r|,�ϩA�PT& ��/��Zc\T0 k� �'�'��d  e1�t B  ��H    �  ��3  LQ$Er� �4r|,�ϩA�PT& ��/��Zc\T0 k� �'�'��d  e1�t B  ��H    �  ��4  LQ Er�! �4s|,�ϩA�PP' ��/��Zc\T0 k� �'�'��d  e1�t B  ��H    �  ��5  LQ Fr�# �4s|,�˩A�PP' ��/��Zc\T0 k� �(�(��d  e1�t B  ��H    �  ��6  LQ Gr�% �8s|,�˩A�PP' ��/��Zc\T0 k� �(�(��d  e1�t B  ��H    �  ��7  LQGr�& �8s|,�˩A�PL' ��/��Zc\T0 k� �(�(��d  e1�t B  ��H    �  ��8  LQHB�( �8s|,�˩A�PL( ��/��Zc\T0 k� �)�)��d  e1�t B  ��H    �  ��9  LQHB�* �8s|,�˩A�PL( ��/��Zc\T0 k� �)�)��d  e1�t B  ��H   �  ��:  LQIB�, �8s|,�˩A�PH( ��/��Zc\T0 k� �)�)��d  e1�t B  ��H    �  ��;  LaIB�. �8s|,�˪A�PH) ��/��Zc\T0 k� � )�)��d  e1�t B  ��H    �  ��<  LaJB�0 �<s|,�˪A�PH) ��/��Zc\T0 k� � *�*��d  e1�t B  ��H    �  ��=  LaK2 �<s|,�˪A�PH) ��/��Zc\T0 k� � *�*��d  e1�t B  ��H    �  ��=  LaK4 �<t|,�˪A�PD) ��/��Zc\T0 k� � *�*��d  e1�t B  ��H    �  ��>  LaL5 �<t|,�ǪA�PD* ��/��Zc\T0 k� ��*� *��d  e1�t B  ��H    �  ��?  LaL7 �<t|,�ǪA�PD* ��/��Zc\T0 k� ��+� +��d  e1�t B  ��H    �  ��@  LaM9 �<t|,�ǪA�P@* ��/��Zc\T0 k� ��+� +��d  e1�t B  ��H    �  ��A  LaM; �<t|,�ǪA�P@* ��/��Zc\T0 k� ��+��+��d  e1�t B  ��H    �  ��B  LaN= �@t|,�ǪA�P@+ ��/��ZcXT0 k� ��+��+��d  e1�t B  ��H    �  ��B  LaN�? �@t|,�ǪA�P@+ ��/��ZcXT0 k� ��,��,��d  e1�t B  ��H    �  ��C  LaO�@ �@t|,�ǪA�P<+ ���/��ZcXT0 k� ��,��,��d  e1�t B  ��H    �  ��D  LaO�B �@t|,�ǪA�P<+ ���/��ZcXT0 k� ��,��,��d  e1�t B  ��H    �  ��E  LaP�D �@t|,�ǪA�P<+ ���/��ZcXT0 k� ��,��,��d  e1�t B  ��H    �  ��F  LaP�|E �@t|,�ǪA�P<, ���/��ZcXT0 k� ��,��,��d  e1�t B  ��H    �  ��F  LaQ�|G �@t|,�ǪA�P8, ���/��ZcXT0 k� ��-��-��d  e1�t B  ��H    �  ��G  LaQ�xI �@u|,�ǪA�P8, ���/��ZcXT0 k� ��-��-��d  e1�t B  ��H    �  �|H  LaQ�xJ �@u|,�êA�P8, ���/��ZcXT0 k� ��-��-��d  e1�t B  ��H    �  �|I  LaR�tL �Du|,�êA�P8, ���/��ZcXT0 k� ��-��-��d  e1�t B  ��H    �  �|I  La R�tN �Du|,�êA�P4- ���/��ZcXT0 k� ��-��-��d  e1�t B  ��H    �  �|J  La S�pO �Du|,�êA�P4- ���/��ZcXT0 k� ��.��.��d  e1�t B  ��H    �  ��|K  La S�pQ �Du|,�êA�P4- ���/��ZcXT0 k� ��.��.��d  e1�t B  ��H    �  ��xK  L`�T�pR �Du|,�ëA�P4- ���/��ZcXT0 k� ��.��.��d  e1�t B  ��H    �  ��xL  L`�T�lT �Du|,�ëA�P4- ���/��ZcXT0 k� ��.��.��d  e1�t B  ��H    �  ��xM  L`�TlU �Du|,�ëA�P0. ���/��ZcXT0 k� ��.��.��d  e1�t B  ��H    �  ��xM  L`�UhV �Du|,�ëA�P0. ���/��ZcXT0 k� ��/��/��d  e1�t B  ��H    �  ��xN  L`�UhX �Du|,�ëA�P0. ���/��ZcXT0 k� ��/��/��d  e1�t B  ��H    �  ��tO  L`�VhY �Hu|,�ëA�P0. ���/��ZcXT0 k� ��/��/��d  e1�t B  ��H    �  ��tO  L`�Vd[ �Hu|,�ëA�P0. ���/��ZcXT0 k� ��/��/��d  e1�t B  ��H    �  ��tP  L`�Vd\ �Hu|,�ëA�P,. ���/��ZcXT0 k� ��/��/��d  e1�t B  ��H    �  ��pQ  L`�W`^ �Hv|,�ëA�P,/ ���/��ZcXT0 k� ��0��0��d  e1�t B  ��H    �  ��pR  L`�W`` �Hu|,���A�P,/ ���/��ZcXT0 k� ��0��0��d  e1�t B  ��H    �  ��lR  L`�X`a �Hu|,���A�P,/ ���/��ZcXT0 k� ��0��0��d  e1�t B  ��H    �  ��lS  L`�X\b �Hu|,���A�P(/ ���/��ZcXT0 k� ��0��0��d  e1�t B  ��H    �  ��hS  L`�X\d �Hu|,���A�P(/ ���/��ZcXT0 k� ��0��0��d  e1�t B  ��H    �  ��hT  L`�Y\e �Hu|,���A�P(0 ���/��ZcXT0 k� ��0��0��d  e1�t B  ��H    �  ��dT  L`�YXe �Hv|,���A�P(0 ���/��ZcXT0 k� ��1��1��d  e1�t B  ��H    �  ��`U  L`�YXf �Hv|,���A�P(0 ���/��ZcXT0 k� ��1��1��d  e1�t B  ��H    �  ��`U  L`�ZXf �Hv|,���A�P(0 ���/��ZcXT0 k� ��1��1��d  e1�t B  ��H    �  ��\V  L`�ZXf �Hv|,���A�P$0 ���/��ZcTT0 k� ��1��1��d  e1�t B  ��H    �  ��XV  L`�ZXf �Hv|,���A�P$0 ���/��ZcTT0 k� ��1��1��d  e1�t B  ��H    �  ��TW  LP�[Xg �Dw|,���A�P$0 ���/��ZcTT0 k� ��1��1��d  e1�t B  ��H    �  ��PW  LP�[Xg �Dw|,���A�P$1 ���B�ZcTT0 k� ��2��2��d  e1�t B  ��H    �  ��PX  LP�[Xg �Dw|,���A�P$1 ���B�ZcTT0 k� ��2��2��d  e1�t B  ��H    �  ��LX  LP�\Xg �Dw|,���A�P$1 ���B�ZcTT0 k� ��2��2��d  e1�t B  ��H    �  ��HY  LP�\\g �Dw|,���A�P$1 ���B�ZcTT0 k� ��2��2��d  e1�t B  ��H    �  ��DY  LP�\\g �@w|,���A�P 1 ���B�ZcTT0 k� ��2��2��d  e1�t B  ��H    �  ��@Z  E��]\g �@w|,���A�P 1 ���B�ZcTT0 k� ��2��2��d  e1�t B  ��H    �  ��<Z  E��]\g �@v|,���A�P 1 ���B�ZcTT0 k� ��2��2��d  e1�t B  ��H    �  ��8[  E��]\g �@v|,���A�P 2 ���B�ZcTT0 k� ��2��2��d  e1�t B  ��H    �  ��4[  E��^\f �@v|,���A�P 2 ���B�ZcTT0 k� ��3��3��d  e1�t B  ��H    �  ��,\  E��^\f �<v|,���A�P 2 ���R�ZcTT0 k� ��3��3��d  e1�t B  ��H    �  ��(\  F �_\f �<u|,���A�P 2 ���R�ZcTT0 k� ��3��3��d  e1�t B  ��H    �  ��$\  F �_\f �<u|,���A�P2 ���R�ZcTT0 k� ��3��3��d  e1�t B  ��H    �  �� ]  F �`\f �<u|,���A�P2 ���R�ZcTT0 k� ��3��3��d  e1�t B  ��H   �  ��]  F �`\f �<u|,���A�P2 ���R�ZcTT0 k� ��3��3��d  e1�t B  ��H    �  ��^  F �a\f �8t|,���A�P2 ���R�ZcTT0 k� ��3��3��d  e1�t B  ��H    �  ��^  F �b\f �8t|,���A�P3 ���R�ZcTT0 k� ��3��3��d  e1�t B  ��H    �  ��^  F �b\f �8t|,���A�P3 ���R�ZcTT0 k� ��4��4��d  e1�t B  ��H    �  �_  E��c\f �8t|,���A�P3 ���R�ZcTT0 k� ��4��4��d  e1�t B  ��H    �  � _  E��d\f �8t|,���A�P3 ���R�ZcTT0 k� ��4��4��d  e1�t B  ��H    �  ��`  E��d\f �4t|,���A�P3 ���R�ZcTT0 k� ��4��4��d  e1�t B  ��H    �  ��`  E��e\f �4t|,���A�P3 ���R�ZcTT0 k� ��4��4��d  e1�t B  ��H    �  ��`  E��e\f �4t|,���A�P3 ���R�ZcTT0 k� ��4��4��d  e1�t B  ��H    �  ��a  E��f�\f �4t|,���A�P3 ���R�ZcTT0 k� ��4��4��d  e1�t B  ��H    �  ���a  E��g�`f �4s|,���A�P3 ���R�ZcTT0 k� ��4��4��d  e1�t B  ��H    �  ���a  E��g�`f �4s|,���A�P3 ���R�ZcTT0 k� ��4��4��d  e1�t B  ��H    �  ���b  B��h�`f �0s|,���A�P4 ���R�ZcTT0 k� ��4��4��d  e1�t B  ��H    �  ���b  B� h�`f �0s|,���A�P4 ���R�ZcTT0 k� ��5��5��d  e1�t B  ��H    �  ���b  B� i�`f �0s|,���A�P4 ���R�b�TT0 k� ��5��5��d  e1�t B  ��H    �  ���c  B�i�`f �0s|,���A�P4 ���R�b�TT0 k� ��5��5��d  e1�t B  ��H    �  ���c  B�j�`f�0r|,���A�P4 ���R�b�TT0 k� ��5��5��d  e1�t B  ��H    �  �Ҹc  B�j�`f�0r|,���A�P4 ���R�b�TT0 k� ��5��5��d  e1�t B  ��H    �  �Ұd  B�k�`f�0r|,���A�P4 ���R�b�TT0 k� ��5��5��d  e1�t B  ��H    �  ��d  B�k�`f�,r|,���A�P4 ���R�b�TT0 k� ��5��5��d  e1�t B  ��H    �  ��d  B�l`f�,r|,���A�P4 ���R�b�TT0 k� ��5��5��d  e1�t B  ��H    �  ��d  B�l\f�,r|,���A�P4 ���R�b�TT0 k� ��5��5��d  e1�t B  ��H    �  ��d  B� mXf�,r|,���A�P4 ���R�b�TT0 k� ��5��5��d  e1�t B  ��H    �  ��d  B�$mXf�,r|,���A�P5 ���R�b�TT0 k� ��5��5��d  e1�t B  ��H    �  �	��d  B�(nTf�(r|,���A�P5 ���R�b�TT0 k� ��6��6��d  e1�t B  ��H    �  �	��d  B�,nTf�(r|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �	��d  B�0oTf�(r|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �	��d  B�4oPf�$r|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �	��d  B�<pPf�$r|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �2�d  B�@pPf�$r|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �2�d  B�DqPf�$r|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �2�d  B�LqPf�$r|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �2�d  B�PrLf�$q|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �2�d  B�TrLf�$q|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �2�d  B�\rLf�$q|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �2�d  E�`sLf� q|,���A�P5 ��R�ZcTT0 k� ��6��6��d  e1�t B  ��H    �  �2�d  E�hsLf� q|,���A�P6 ��R�b�TT0 k� ��6��6��d  e1�t B  ��H    �  �2�d  E�ltLf� q|,���A�P6 ��R�b�TT0 k� ��7��7��d  e1�t B  ��H    �  �2�d  E�ttLf� q|,���A�P6 ��R�b�TT0 k� ��7��7��d  e1�t B  ��H    �  �2�d  E�|tLf� q|,���A�P6 ��R�b�TT0 k� ��7��7��d  e1�t B  ��H    �  �2�d  E��uLf�q|,���A�P6 ��R�b�TT0 k� ��7��7��d  e1�t B  ��H    �  �2�d  E��uRLf�q|,���A�P6 ��R�b�TT0 k� ��7��7��d  e1�t B  ��H    �  �2�d  E��uRLf�q|,���A�P6 ��R�b�TT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  E��vRLf�q|,���A�P6 ��R�b�TT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  E��vRLf�q|,���A�P6 ��R�b�TT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  E��vRHf�q|,���A�P6 ��R�b�TT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  E��wHf�q|,���A�P6 ��R�b�TT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  E��wHf�q|,���A�P6 ��R�ZcTT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  E��wHf�q|,���A�P6 ��R�ZcTT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  B��wHf�q|,���A�P6 ��R�ZcTT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  B��wHf�q|,���A�P6 ��R�ZcTT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  B��wHf�q|,���A�P6 ��R�ZcTT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  B��wHf�q|,���A�P7 ��R�ZcTT0 k� ��7��7��d  e1�t B  ��H    �  �B�d  B��wHf�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��wHf�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��xHf�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��x"Hf�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��x"Hf�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��y"He�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��y"He�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��y"He�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��y"He�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��y"He�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��y"He�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��y"He�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��z"He�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��z"He�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��z"He�q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��z"He� q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��z"He� q|,���A�P7 ��R�ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��z"He� q|,���A�P7 ��R �ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��z"He� q|,���A�P7 ��R �ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��z"He�$q|,���A�P7 ��R �ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�d  K��z"He�$q|,���A�P8 ��R �ZcTT0 k� ��8��8��d  e1�t B  ��H    �  �B�c  K��z"He�$q|,���A�P8 ��R �ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �B�c  K��z"He�$q|,���A�P8 ��R �ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �B�c  K��z"He�$q|,���A�P8 ��R �ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �B�c  K��z"He �$q|,���A�P8 ��R �ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �B�c  K��z"He �$q|,���A�P8 ��R$�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �B�c  K��z"He �$q|,���A�P8 ��R$�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �B�c  K��z"He �$q|,���A�P8 ��R$�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �B�c  K��z"He �$q|,���A�P8 ��R$�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �B�c  K��z"He �$q|,���A�P8 ��R(�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �B�c  K��z"He �$q|,���A�P8 ��R(�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��z"He �(q|,���A�P8 ��R(�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��z"He �(q|,���A�P8 ��R(�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��z"He �(q|,���A�P8 ��R,�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��z"He �(q|,���A�P8 ��R,�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��z"He �(q|,���A�P8 ��R,�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��z"He �(q!�,���A�P8 ��R,�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��z"He �(p!�,���A�P8 ��R0�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��z"He �(p!�,���A�P8 ��R0�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  ���c  K��z"He �(p!�,���A�P8 ��R0�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  ���c  K��z"He �(p!�,���A�P8 ��R4�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  ���c  K��z"He �(p!�,���A�P8 ��R4�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  ���c  K��z"He �(p!�,���A�P8 ��R4�ZcTT0 k� ��9��9��d  e1�t B  ��H    �  ���c  K��z"Hd �(o!�,���A�P8 ��R4ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��zHd �,o!�,���A�P8 ��R8ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��zHd �,o!�,���A�P8 ��R8ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��zHd �,o!�,���A�P8 ��R8ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�c  K��zHd �,o|,���A�P9 ��R8ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�b  K��zHd �,o|,���A�P9 ��R<ZcTT0 k� ��9��9��d  e1�t B  ��H    �  �2�b  K��zHd �,n|,���A�P9 ��R<ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �2�b  K��zHd �,n|,���A�P9 ��R<ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �2�b  K��zHd �,n|,���A�P9 ��R<ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �2�a  K��zHd �,n|,���A�P9 ��R@~ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �2�a  K��zHd �,n|,���A�P9 ��R@~ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �B�a  K��zHd �,n|,���A�P9 ��R@~ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �B�`  K��zHd �,n|,���A�P9 ��R@~ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �B�`  K��zRHd �,n|,���A�P9 ��RD}ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �B�`  K��zRHd �,n|,���A�P9 ��RD}ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �B�`  K��zRHd �,n!�,���A�P9 ��RD}ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �B�`  K��zRHd �,n!�,���A�P9 ��RD}ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �B�`  K��zRHd �,n!�,���A�P9 ��RH}ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �B�`  K��zRHd �,n!�,���A�P9 ��RH}ZcTT0 k� ��:��:��d  e1�t B  ��H    �  �B�`  B��zRHd �,n!�,���A�P9 ��RH}ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ���`  B��zRHd �,n!�,���A�P9 ��RH}ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ���`  B��zRHd �,n!�,���A�P9 ��RL}ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ���`  B��yRHd �,n!�,���A�P9 ��RL}ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ���`  B��yRHd �,n!�,���A�P9 ��RL|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ���`  B��yRHd �,n!�,���A�P9 ��RL|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��`  B��yRHd �,n!�,���A�P9 ��RP|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��`  B��yRHd �,n|,���A�P9 ��RP|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��`  B��yRHd �,n|,���A�P9 ��RP|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��`  B��yRHd �,n|,���A�P9 ��RP|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��_  B��yRHd �,n|,���A�P9 ��RP|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��_  B��yRHd �,n|,���A�P9 ��RT|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��_  C�yRHd �,n|,���A�P9 ��RT|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��_  C�yRHd �,n|,���A�P9 ��RT|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��_  C�yRHd �,n|,���A�P9 ��RT|ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��_  C�yRHd �,n|,���A�P9 ��RX{ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��_  C�yRHd �,n|,���A�P9 ��RX{ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��_  C�yRHd �,n|,���A�P9 ��RX{ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��_  C�yRHd �,n|,���A�P9 ��RX{ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ��_  C�yRHd �,n|,���A�P9 ��R\{ZcTT0 k� ��:��:��d  e1�t B  ��H    �  ���  E�� 1�����|,��F �\�.�'��ÑZ3� T0 k� ��������d  e1�t B  ��3   �  ���  E�� 1�����|,��F �^�-�/��ˑZ3� T0 k� �������d  e1�t B  ��3   �  ���  E� 1�����|,��E��`�,�7��ӑZ3� T0 k� ������d  e1�t B  ��3   �  �Æ  E� 1�����|,��E��a�,�?��ۑZ3� T0 k� ������d  e1�t B  ��3   �  �Æ  E� 1�����|,���E��c�+�G���Z3� T0 k� �#��'���d  e1�t B  �3   �  �Æ  E�A�����|,���E��e� *�S���Z3� T0 k� �;��?���d  e1�t B  ��?   �  �Æ  B�'�A�����|,���E��f�$*�[���Z3� T0 k� �O��S���d  e1�t B ��?   �  �Ǉ  B�7�A�����|,���B��j((�k���Z3��T0 k� �w��{���d  e1�t B ��?   �  ��Ǉ  B�?�A�����|,���B��k,'�s���Z3��T0 k� ��������d  e1�t B ��?   �  ��ˇ  B�G�A�����|,���B��m0&�{���Z3��T0 k� ��������d  e1�t B ��?   �  ��ˇ  B�O�Q�����|,���B��n4%�����Z3��T0 k� ��������d  e1�t B ��?   �  ��χ  B�W�Q����|,���B��p8$����#�Z3��T0 k� ��������d  e1�t B ��?   �  ��χ  B�_�Q����|,���B��qr<#����+�Z3��T0 k� ��������d  e1�t B ��?   �  ��Ӈ  B�g�Q����|,���B�sr@"����/�Z3��T0 k� ��������d  e1�t B ��?   �  ��ӈ  B�o�Q����|,��B�trD!��� 7�Z3��T0 k� ������d  e1�t B ��?   �  ��׈  B�w�b��+�|,� B�vrH ��� ?�Z3��T0 k� �#��'���d  e1�t B ��?   �  ��׈  B��b��3�|,�B�wrL��� G�Z3��T0 k� �7��;���d  e1�t B ��?   �  ��ۈ  B���b��;�|,�B� xP��� O�^��T0 k� �O��S���d  e1�t B ��?   �  ��߈  B���b��C�|,�$B�$zTB�� W�^��T0 k� �c��g���d  e1�t B ��?   �  ���  B���b��K�|,�,E�,{XBü _�^��T0 k� �w��{���d  e1�t B ��?   �  ���  B���b#��S�|,4E�4|`B˽ g�^��T0 k� ��������d  e1�t B ��?   �  ���  B���b'��[�|,<E�<~dBӾ o�^��T0 k� ��������d  e1�t B ��?   �  ���  B���b/��c�|,DE�@hBۿ w�^��T0 k� ��������d  e1�t B ��?  �  ���  B���b3��o�|,LE�H�l"�� �^��T0 k� ��������d  e1�t B �?   �  ���  B���b7��w�|,T	E�P�p"�� ��^��T0 k� 3�������d  e1�t B ��?   �  ����  B���b?���|,\
E�X��x"����^��T0 k� 3�������d  e1�t B ��?   �  ����  B���bC�އ�|,dE�`�|"����^��T0 k� 3�������d  e1�t B ��?   �  ����  B���bG�ޏ�|,lE�d҈"����^��T0 k� 3�������d  e1�t B ��?   �  ���  B���bO�ޗ�|,�tE�lҐ#���^��T0 k� 3�������d  e1�t B ��?   �  ���  B���bS�ޟ�|,�|E�t~Ҙ
#���^��T0 k� ��������d  e1�t B ��?   �  ���  B���bW����|,��E�|~¤#���^��T0 k� ��������d  e1�t B ��?   �  ���  B���b[����|,��E��}¬���^��T0 k� ��������d  e1�t B ��?   �  ���  B��bc����|,��E��|´�Þ^��T0 k� ��������d  e1�t B ��?  �  ���  B��bg��ú|,ќE��|¼ '�˞^��T0 k� ��������d  e1�t B ��?   �  ���  B��bk��˺|,ѤE��{���/�ϟ^��T0 k� �������d  e1�t B ��?   �  ��#�  B��bo��ӹ|,ѬE��z���7�נ^��T0 k� �������d  e1�t B	 ��?   �  ��'�  B�'��s��۹|,ѴB�z���?� ߡ^��T0 k� �������d  e1�t B	 ��?   �  ��/�  B�/��{���|,��B�y���G� �^��T0 k� �������d  e1�t B	 ��?   �  ��3�  B�7�����|,��B�x���K� �^��T0 k� �������d  e1�t B
 ��?   �  ��7�  B�C�������|,��B��w���S� ��^��T0 k� C�������d  e1�t B
 ��?   �  ��?�  B�K�������|,��B��w���	[� ��^��T0 k� C�������d  e1�t B
 ��?   � 
 ��C�  B�S������|,��E�v��	c�!�^��T0 k� C�������d  e1�t B
 ��?   � 	 ��K�  B�[������|,��E�u��	g�!�^��T0 k� C�������d  e1�t B
 ��?   �  ��O�  B�c������|,��E�t��	o�!�^��T0 k� C������d  e1�t B ��?   �  ��W�  B�k�����#�|,��E�s��	w�!�^��T0 k� #{�����d  e1�t B ��?   �  ��[�  B�s�����+�|,�E�s�#�	{�!�^��T0 k� #w��{���d  e1�t B ��?   �  ��c�  B�{�����3�|,�E�r�'�	#��!'�^��T0 k� #s��w���d  e1�t B $�?   �  ��g�  B҃�����;�|,�Eq�/�	#���/�^��T0 k� #s��w���d  e1�t B ��?   �  ��s�  Bҗ�����O�|,�(Ep�?�	#���?�^��T0 k� �o��s���d  e1�t B ��?   �  ��{�  Bҟ�����W�|,�0B�o�C�	#���C�^��T0 k� �o��s���d  e1�t B ��?   �  �߃�  E������_�|,�8B�$n�K�$���K�Z3��T0 k� �o��s���d  e1�t B
 ��?   �  �߇�  E������g�|,�@B�,n�S�$���S�Z3��T0 k� �o��s���d  e1�t B
 ��?   �  ����  E������o�|,�HB�4msW�$���[�Z3��T0 k� �k��o���d  e1�t B
 ��?   �  ����  E�����{�|,rPB�<ms_�$���_�Z3��T0 k� �k��o���d  e1�t B
 ��?   �  ����  E����σ�|,r\IDlsg�$���g�Z3��T0 k� �k��o���d  e1�t B
 ��?   �  ����  E����ϋ�|,rdILlsk�$#���o�Z��T0 k� �k��o���d  e1�t B	 ��?   �  ����  E����ϓ�|,rlIPkss�$#���w�Z��T0 k� #k��o���d  e1�t B	 ��?   �  ����  E�������|,rtIXksw�$#���{�Z��T0 k� #g��k���d  e1�t B	 ��?   �  ����  E������|,|I`ks�$#����Z��T0 k� #g��k���d  e1�t B ��?   �  ����  E������|,�I"djs��$#����Z��T0 k� #g��k���d  e1�t B ��?   �  ��Ǎ  E�������|,�I"ljs��$#����Z��T0 k� #g��k���d  e1�t B ��?   �  ��ύ  E������|,�I"pjs������Z��T0 k� �g��k���d  e1�t B ��?   �  ��׍  E��'��Ǯ|,�I"tjs������Z��T0 k� �c��g���d  e1�t B ��?   �  ��ۍ  E���/��Ϯ|,�I"xjc������Z��T0 k� �c��g���d  e1�t B ��?   �  ���  E���3��ۭ|,�I�ic������Z��T0 k� �c��g���d  e1�t B ��?   �  ���  E�+��C���|,r�I�ic������Z��T0 k� �c��g���d  e1�t B ��?   �  ����  E�7��K���|,r�
I�ic������Z��T0 k� �_��c���d  e1�t B ��3   �  ����  E�?��S����|,r�	I�ic����ǾZ��T0 k� #g��k���d  e1�t B ��3  �  ���  E�G��[���|,r�I"�ic���ϿZ��T0 k� #o��s���d  e1�t B ��3   �  ���  E�O��c���|,r�I"�ic�����Z3��T0 k� #w��{���d  e1�t B ��3   �  ���  E�_��s���|,r�I"�ic������Z3��T0 k� #�������d  e1�t B ��3   �  �#�  Esg��{��'�|,r�I"�icî����Z3��T0 k� ��������d  e1�t B  ��3   �  �+�  Eso����3�|,r�I�icǬ�#���Z3��T0 k� ��������d  e1�t B  ,�3  �  �7�  Es�����C�|,sI�iS˨�/���Z��T0 k� ��������d  e1�t B  ��3   �  �?�  Es��s���K�|,s I�iSϦ�3��Z��T0 k� ��������d  e1�t B  ��3   �  �G�  Es��s���S�|,s�I�iSϤ�7��Z��T0 k� ��������d  e1�t B ��3   �  �O�  Es��s���_�|,s#�I"�iSϢ�;��Z��T0 k� ��������d  e1�t B �3   �  �[�  Es��s���o�|,s3�I"�iSӞ�G�"�Z��T0 k� #�������d  e1�t B ��?   �  �c�  Es������w�|,s7�I"�iSӜ�K�"#�Z��T0 k� #�������d  e1�t B ��?   �  �k�  Es�������|,s?�I"�iSӚ�O�"+�Z��T0 k� #�������d  e1�t B ��?   �  �o�  Es��������|,sC�I�iSӘtS�"3�Z��T0 k� #�������d  e1�t B ��?   �  �w�  Ec������|,sK�I�iSӖt[�"7�Z��T0 k� #�������d  e1�t B ��;   �  Ї�  Ec������|,sW�I�iSӒtc�"G�_s��T0 k� C�������d  e1�t B �;   �  Ћ�  Ec������|,s_�I�iSӐtg�"K�_s��T0 k� C�������d  e1�t B ��;   �  Г�  Ec����� ��|,sc�I"�iSώto��S�_s��T0 k� C�������d  e1�t B ��;   �  Л�  Ec����� ��|,ck�I"�iCύts��[�_s��T0 k� C�������d  e1�t B ��;   �  Ч�  Ec����� Ϯ|,cw�I"�iCˉt{��g�_s��T0 k� ��������d  e1�t B ��;   �  Я�  Ec����� ׯ|,c{�I"�iCˈt��k�_s��T0 k� ��������d  e1�t B ��;   �  ���  Ec����� ߯|,c�I�iCǆt���s�_t�T0 k� ��������d  e1�t B ��;   �  ���  Ec����� �|,c��I�i�ǅt���{�_t�T0 k� ��������d  e1�t B ��;   �  �Ǐ  ES����� �|,c��I�i�Ät����_t�T0 k� ��������d  e1�t B ��;   �  �ˏ  ES����� ��|,c��I�i�Ât�����_t�T0 k� ��������d  e1�t B ��;   �  �ۏ  ES������|,c��@b�i���d�����_t�T0 k� ��������d  e1�t B  ��;   �  ��  ES������|,c��@b�i���d�����_��T0 k� ��������d  e1�t B  ��;   �  ��  C�������|,S��@b�i���d�����_��T0 k� ��������d  e1�t B  �;   �  ��  C������'�|,S��@b�i���d�����_��T0 k� 3�������d  e1�t B  /�;   �  ���  C������/�|,S��@b�i���d�����_��T0 k� 3�������d  e1�t B  ��;   �  ���  C������7�|,S��@��i���d�����_��T0 k� 3�������d  e1�t B  ��;   �  ��  OS������G�|,S��@��i���d�����_��T0 k� 3�������d  e1�t B  ��;   �  ��  OS������O�|,S��@��i���d�����_��T0 k� #�������d  e1�t B  ��;   �  ��  OS������W�|,S��@��i���d�����_��T0 k� #�������d  e1�t B  ��;   �  ��  OS������c�|,c��A�i���d�����_��T0 k� #�������d  e1�t B  ��;   �  ��'�  OS������k�|,c��A�i���d��B��_��T0 k� #�������d  e1�t B  ��;   �  ��/�  OS������s�|,c��A�i���T��B��_��T0 k� #�������d  e1�t B  ��;   �  ��7�  OS������{�|,c��A�i���T��B��_���T0 k� ��������d  e1�t B  ��;   �  ��;�  OS��������|,c��A�i��T�B��_���T0 k� ��������d  e1�t B  ��;   �  ��C�  OS��������|,c��C��i�{�T{�B��_���T0 k� ��������d  e1�t B  ��;   �  ��K�  OS��������|,c��C��i�w�T{����_���T0 k� ��������d  e1�t B  ��;   �  ��S�  OS��������|,s��C��i�o�Tw����_���T0 k� �������d  e1�t B  ��;   �  ��_�  OS��������|,s��C�i�g�To����_���T0 k� �������d  e1�t B  ��;   �  ��g�  OS��������|,s��C�i�_��k���_���T0 k� �������d  e1�t B  ��;   �  ��o�  OS��������|,s��C�i�[��g���_���T0 k� �������d  e1�t B  ��;   �  ��s�  OS��������|,s��C�i�S��c���_���T0 k� �������d  e1�t B  ��;  �  ��{�  OS��������|,s��C�i�O��[�� _���T0 k� �������d  e1�t B  ��;   �  ��  OS��������|,s��C�i�G��W��_���T0 k� �������d  e1�t B  ��;   �  ��  OS��������|,s��C�i�?�TS��_���T0 k� �������d  e1�t B  ��K   �  ��  OS��������|,s��C�i�3�TG�� _���T0 k� �������d  e1�t B  ��K   �  ���  OS��������|,s��C�i�/�TC��$_���T0 k� �������d  e1�t B  ��K   �  ���  C��������|,s��C�i�'�T?��(
_���T0 k� �������d  e1�t B  ��K   �  ���  C��������|,s��C�i��T7��,_���T0 k� �������d  e1�t B  ��K   �  ���  C�������|,s��C�i��T+��4_���T0 k� �������d  e1�t B  ��K   �  ���  C�������|,s��C�i��T'��4_���T0 k� �������d  e1�t B  ��K   �  �Ǚ  C�������|,s��C�i��T��8_���T0 k� �������d  e1�t B  ��K   �  �˙  C�������|,s��C�i���D��<_���T0 k� �������d  e1�t B  ��K   �  �Ӛ  C�������|,s��D|i���D��<_���T0 k� �������d  e1�t B  ��K   �  �ߛ  C������'�|,s��Dpi��D��@_���T0 k� �������d  e1�t B  ��K   �  ��  C�����2+�|,s��Dli�ߡC���D_���T0 k� �������d  e1�t B  ��K   �  ��  C�����2/�|,s��Ddi�ףC���D_���T0 k� �������d  e1�t B  ��K   �  ��  C�����23�|,s��D`i�ϤC��D_���T0 k� �������d  e1�t B  �K   �  ��  C�����2?�|,s��DPi���C��H!_���T0 k� �����d  e1�t B  ��O   �  ��  C�����2C�|,s��EBLi���CۓSH#[���T0 k� �����d  e1�t B  ��O   �  ��  C�����2G�|,s��EBDi���CӒSH$[���T0 k� �����d  e1�t B  ��O   �  ��  C�����2K�|,s��EB<i���CӒSH&[���T0 k� �����d  e1�t B  ��O   �  ��  C�����2O�|,s��EB4i���CϑSH'[���T0 k� �����d  e1�t B  ��O   �  �'�  C�w����2W�|,s��EB(h���3ǏCH*[���T0 k� �����d  e1�t B  ��O  �  �"/�  C�o����B[�|,s��EB h���3ǏCH,[���T0 k� �|����d  e1�t B  ��O   �  �"7�  C�k����B_�|,s��EBg���3ÎCH.[���T0 k� �x�|��d  e1�t B  ��O   �  �";�  E�g����Bc�|,s��EBg�{�3��CH/[���T0 k� �p!�t!��d  e1�t B  ��O   �  �"G�  E�[���Bk�|,s��EBf�o�3��CH2[���T0 k� �h'�l'��d  e1�t B  ��O   �  �O�  E�W���Bo�|,s�EA�f�g�C���H4[���T0 k� �`*�d*��d  e1�t B  ��O   �  �W�  E�S��{�Bs�|,s{�E1�e�_�C���D6[���T0 k� �\-�`-��d  e1�t B  ��O   �  �[�  E�K��{�Bw�|,s{�E1�d�W�C���D7[���T0 k� �X0�\0��d  e1�t B  ��O   �  �c�  E�G��w�B{�|,sw�E1�d�O�C���D9[���T0 k� �D4�H4��d  e1�t B  ��J   �  �o�  E�;��w�B�!�,so�E1�b�?�C���@;[���T0 k� �87�<7��d  e1�t B  ��J   �  �w�  E�7��s�B�!�,so�E1�a�;�C���<=[���T0 k� �08�48��d  e1�t B  ��J   � 	 �{�  D3/��s�R�!�,sk�E��`�3�C���<>[���T0 k� �(:�,:��d  e1�t B  ��J   � 
 ���  D3+��o�R�!�,sk�E��`�+�C���8@[���T0 k� �$;�(;��d  e1�t B  ��J   �  ���  D3'��o�R�
!�,sg�E��_�#�C���4A[���T0 k� �=� =��d  e1�t B  ��J   �  ����  D3��k�R�!�,sc�E��]��C��c0D[���T0 k� �@�@��d  e1�t B  ��J   �  ����  ES��k�R�!�,s_�E��\��S��c,E[���T0 k� ��C��C��d  e1�t B  ��J   �  ����  ES��k� ��!�,s[�E��[��S��c(G[���T0 k� ��E��E��d  e1�t B  ��J   �  ����  ES��g� ��!�,s[�E��Y���S��c(H[���T0 k� ��F��F��d  e1�t B  ��J   �  ����  ER���g� ��|,sW�E��X���S��c$I[���T0 k� ��H��H��d  e1�t B  ��J   �  ���  ER���c� ��|,sW�E��W���S��C K[���T0 k� ��N��N��d  e1�t B  ��J   �  ���  ER���c� ��|,sS�C��V���S�CL[���T0 k� ��S��S��d  e1�t B  �J    �  �˲  E����_� ��|,sO�C�pT��� �{�CO[���T0 k� ��X��X��d  e1�t B  �J    �  �Ӳ  E����_� ��|,sK�C�hS��� �w�CP[���T0 k� ��\��\��d  e1�t B  ��J    �  ��۳  E����_� ��!|,sK�C�dR��� �w�CRZc��T0 k� ��^��^��d  e1�t B  ��J    �  ��ߴ  E����[�´"|,sG�A\Q��� �s�CSZc��T0 k� ��a��a��d  e1�t B  ��J    �  ���  E����[�¸&|,sC�ALNѳ� �o�C VZc��T0 k� ��e��e��d  e1�t B  ��J    �  ���  E���W�¼(|,sC�AHMѯ� �o��WZc��T0 k� ��f��f��d  e1�t B  ��J    �  ����  E���W�¼*!�,s?�A@Lѧ� �o��YZc��T0 k� ��h��h��d  e1�t B  ��J    �  ���  E���W���,!�,s?�A8KQ�� �k��[Zc��T0 k� ��i��i��d  e1�t B  ��J    �  ���  E���W���-!�,s;�A4JQ�� �k��\Zc��T0 k� �k��k��d  e1�t B  ��J    �  ���  E���S���/!�,s;�A,IQ�� �g��^Zc��T0 k� �l��l��d  e1�t B  ��J   �  ���  E���S���1!�,s7�A(IQ�� �g���_Zc��T0 k� �i��i��d  e1�t B  ��J    �  ���  E���S���3!�,s7�A HQ�� �c���`Zc��T0 k� �g��g��d  e1�t B  ��J    �  ��#�  E���O���5!�,s3�AGQ� �c���bZc��T0 k� �f��f��d  e1�t B  ��J    �  ��+�  E���O���8!�,s/�AFQ{� �_���cZc��T0 k� �e��e��d  e1�t B  ��J    �  ��/�  E�w��O���;!�,s/�AEQs� �_���eZc��T0 k� �d��d��d  e1�t B  �J    �  ��7�  E�s��O���>!�,s+�ADQo� �[���fZc��T0 k� �b��b��d  e1�t B ��O    �  ��?�  E�k��K���A!�,s+�ACQg� �[���gZc��T0 k� �a��a��d  e1�t B ��O    �  ��C�  E�c��K���D|,s'�A �BQc� �W���iZc��T0 k� �_��_��d  e1�t B ��O    �  ��K�  E�_��K���G|,s'�A �AQ_� �W���jZc��T0 k� �t]�x]��d  e1�t B ��O    �  ��O�  D�W��K���J|,s'�A �AQW� �W�¼kZc��T0 k� �h\�l\��d  e1�t B ��O   �  ��W�  D�O��G���L|,s#�A �@QS� �S�´lZc��T0 k� �\Z�`Z��d  e1�t B ��O    �  �C[�  D�K��G���O|,s#�A �?QO� �S�ҰnZc��T0 k� �PY�TY��d  e1�t B ��O    �  �Cc�  D�C��G���R|,s�A �>QG� �O�ҬoZc��T0 k� �DW�HW��d  e1�t B ��O    �  �Cg�  D�?��G���T|,s�A �=QC� �O�ҨpZc��T0 k� �8V�<V��d  e1�t B ��O    �  �Co�  D�7��C���W|,s�A �=Q?� �O�ҤqZc��T0 k� �,T�0T��d  e1�t B ��O    �  �Cs�  D�3��C���Y|,s�A �<Q7� �K�ҠrZc��T0 k� � S�$S��d  e1�t B ��O    �  ��w�  D�+��C���\|,s�A �;Q3� �K��sZc��T0 k� �Q�Q��d  e1�t B ��O   �  ���  D�'��C���^|,s�A �:Q/� �G��uZc��T0 k� �O�O��d  e1�t B ��O    �  ����  D���?���a|,s�A �:Q+� �G��vZc��T0 k� ��N� N��d  e1�t B ��O   �  ����  D���?���c|,s�A �9Q'� �G��wZc��T0 k� ��L��L��d  e1�t B ��O    �  ����  D���?���e|,s�A �8Q� �C��xZc��T0 k� ��K��K��d  e1�t B ��O    �  ����  D���?���h|,s�A �8Q� �C��yZc��T0 k� ��I��I��d  e1�t B ��O    �  �×�  D��s?���h|,s�A �7Q� �C��zZc��T0 k� ��H��H��d  e1�t B ��O    �  �Û�  D��s;�B�j|,s�A �6Q� �?��|Zc��T0 k� ��F��F��d  e1�t B  �O    �  �ß�  D�� s;�B�i|,s�A �6Q  �?��|~Zc��T0 k� �E��E��d  e1�t B ��O    �  �ã�  D��s;�B�i|,s�A �5Q �?��|Zc| T0 k� �C��C��d  e1�t B  �O    �  �ç�  LQ�s;�B|h|,s�A �4Q �;��xZc| T0 k� �A��A��d  e1�t B ��O    �  �ë�  LQ�s;�Bxh|,s�A �4Q  �;��t~Zc| T0 k� �@��@��d  e1�t B ��O    �  �ï�  LQ�s7�Bxh|,s�A �3P� �;��p~Zc| T0 k� �>��>��d  e1�t B ��O    �  �ó�  LQ�s7�Btg|,s�A �3P� �7��l~Zc| T0 k� �x=�|=��d  e1�t B ��O    �  �÷�  LQ�	s7�Bpg|,s�A �2P� �7��h}Zcx T0 k� �l;�p;��d  e1�t B ��O    �  �û�  LQ��7�Bpg|,s�A �1P� �7��h}Zcx T0 k� �`:�d:��d  e1�t B ��O    �  ����  LQ��7�Blf|,s�A �1P� �3��d}Zcx T0 k� �T8�X8��d  e1�t B ��O    �  ����  LQ��7�Bhf|,���A �0P� �3��`|Zcx T0 k� �H7�L7��d  e1�t B ��O    �  ����  LQ��3�Bhf|,���A �0P� �3��\|ZcxT0 k� �<5�@5��d  e1�t B ��O    �  ����  LQ��3�Bde|,���A �/P�	 �3��\|ZcxT0 k� �04�44��d  e1�t B ��O    �  ����  LQ�c3�Bde|,���A |/P�
 �/��X{ZctT0 k� �$2�(2��d  e1�t B ��O    �  ����  LQ�c3�B`e|,���A |.P�
 �/�RT{ZctT0 k� �0�0��d  e1�t B ��O    �  ����  LQ�c/�B\d|,���A x.P� �/�RP{ZctT0 k� �/�/��d  e1�t B ��O    �  ����  LQ�c/�B\d|,���A t-P� �/�RPzZctT0 k� � -�-��d  e1�t B ��O    �  ����  La�c+�BXd|,���A p-P� �+�RLzZctT0 k� ��,��,��d  e1�t B ��O    �  ����  La�S+�BXd|,���A l,P� �+�RHzZctT0 k� ��*��*��d  e1�t B ��O    �  ����  La�S'�BTc|,b��A h,P� �+�RHzZcpT0 k� ��)��)��d  e1�t B ��O    �  ����  La�S'�BTc|,b�A h+P� �+�RDyZcpT0 k� ��'��'��d  e1�t B ��O    �  ����  La�S#�BPc|,b�A d+P� �'�R@yZcpT0 k� ��&��&��d  e1�t B ��O    �  ����  La�S�BLb|,b�A `*P� �'�R@yZcpT0 k� �$��$��d  e1�t B ��O    �  ����  La�C�BLb|,b�A \*P� �'�R<xZcpT0 k� �"��"��d  e1�t B ��O    �  ����  La�C�BHb|,b�A \)P� �'�R<xZcpT0 k� �!��!��d  e1�t B ��O    �  ����  La�C�BHb|,b�A X)P� �#�R8xZcpT0 k� �����d  e1�t B ��O    �  ����  La� C�Da|,b�A T(P� �#�R4xZclT0 k� ������d  e1�t B ��O    �  ����  La�!C�Da|,b�A T(P� �#�R4wZclT0 k� �x�|��d  e1�t B ��O    �  ����  La�"C�@a|,��A P(P� �#�R0wZclT0 k� �l�p��d  e1�t B ��O    �  ����  La�#3�@a|,��A L'P� �#�R0wZclT0 k� �`�d��d  e1�t B  ��H    �  ����  La�$3�<`|,��A L'P� ��R,wZclT0 k� �`�d��d  e1�t B  -�H    �  ����  La�%3�B<`|,��A H&P� ��R,vZclT0 k� �\�`��d  e1�t B  ��H    �  ����  La�&3�B8`|,��A D&P� ��R(vZclT0 k� �X�\��d  e1�t B  ��H    �  ����  La|'2��B8`|,��A D&P� ��R(vZclT0 k� �X�\��d  e1�t B  ��H    �  ����  La|(B��B4`|,��A @%P� ��R$vZclT0 k� �T�X��d  e1�t B ��H    �  ����  Lax)B��B4`|,��A <%P� ��R$vZchT0 k� �P�T��d  e1�t B ��H    �  ����  Lat*B��20`|,��A <$P� ��R uZchT0 k� �P�T��d  e1�t B ��H    �  ���  Lat+B��20b|,��A 8$P� ��R uZchT0 k� �L�P��d  e1�t B ��H    �  ���  Lap,B��2,c|,��A 8$P� ��RuZchT0 k� �H�L��d  e1�t B ��H    �  ���  Lal-B��2(e|,��A 4#P� ��RuZchT0 k� �H�L��d  e1�t B ��H    �  ���  Lah.B��2(e|,��A 0#P� ��/�{ZchT0 k� �D�H��d  e1�t B �H    �  ���  Lah.B��4(f|,�ߧA 0#P� ��/�~ZchT0 k� �D�H��d  e1�t B ��H    �  ���	  Lad/B��4(g|,�ߧA ,"P� ��/��ZchT0 k� �@�D��d  e1�t B ��H    �  ���
  La`0B��4(h|,�ߧA ,"P� ��/��ZchT0 k� �@�D��d  e1�t B ��H    �  ���  La`1B��4(i|,�ߧA ("P� ��/��ZcdT0 k� �<�@��d  e1�t B ��H    �  ���  La\2R��4(j|,�ߧA (!P� ��/��ZcdT0 k� �8�<��d  e1�t B $�H    �  ���  LaX2R��4(j|,�ߧA $!P� ��/��ZcdT0 k�  <�@��d  e1�t B ��H    �  ��  LaX3R��4,k|,�ۧA $!P� ��/��ZcdT0 k�  8�<��d  e1�t B ��H    �  ��  LaT4R��4,l|,�ۧA   P| ��/��ZcdT0 k�  8�<��d  e1�t B ��H    �  ��  LaT5R��4,m|,�ۧA   P| ��/��ZcdT0 k�  4�8��d  e1�t B ��H    �  ��  LaP5R��4,m|,�ۧA  Px ��/��ZcdT0 k�  4�8��d  e1�t B ��H    �  ��  LaL6R��4,n|,�ۧA  Px ��/��ZcdT0 k�  0�4��d  e1�t B ��H    �  ��  LaL7R��4,o|,�ۨA Pt ��/��ZcdT0 k� �0 �4 ��d  e1�t B  ��H    �  ��  LaH7R�4,o|,�רA Pt  ��/��ZcdT0 k� �, �0 ��d  e1�t B  ��H    �  ��  LaH8R�4,p|,�רA Pp  ��/��ZcdT0 k� �,!�0!��d  e1�t B  ��H   �  ��  LaD9R�4,q|,�רA Pp  ��/��ZcdT0 k� �(!�,!��d  e1�t B  ��H    �  ��  LaD9b�4,q|,�רA Pl! ��/��Zc`T0 k� �(!�,!��d  e1�t B  /�H    �  ��   La@:b�4,r|,�רA Pl! ��/��Zc`T0 k� 0$"�("��d  e1�t B  ��H    �  ��!  LQ@;b�4,r|,�רA Pl! ��/��Zc`T0 k� 0$"�("��d  e1�t B  ��H    �  ��"  LQ<;b�4,r|,�ӨA Ph" ��/��Zc`T0 k� 0 "�$"��d  e1�t B  ��H    �  ��$  LQ<<b�
4,r|,�ӨA Ph" ��/��Zc`T0 k� 0 #�$#��d  e1�t B  ��H    �  ��%  LQ8=b�4,r|,�ӨA Pd# ��/��Zc`T0 k� 0 #�$#��d  e1�t B  ��H    �  ��&  LQ8=b�4,r|,�ӨA Pd# ��/��Zc`T0 k� �$� $��d  e1�t B  ��H    �  ��'  LQ4>b�4,r|,�ӨA P`# ��/��Zc`T0 k� �$� $��d  e1�t B  ��H   �  ��)  E�4>b�40r|,�ӨA P`$ ��/��Zc`T0 k� �$�$��d  e1�t B  ��H    �  �                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��N ]�%�%� � �� _��   ? ? 
   � �t     _�� �W           
         	 Z �          Р�    ���  
@				         ��         �  �    ��  �               ��     	 ���         ��       ���  0
 
          yͲ  0 0       V     y�` ֤    ���   
        > Z �         ���    ���   8
	           d:*     
	   �H     dL� ��    �{                	 Z �          �       ���   8          n�n       . �H�     n�� �$    �G)   
          0  Z �          ��     ���   P	          K  ��	      B��-     K��-                              ����               �  ���   P          ��ض        V �Q�    ��ض �Q�                       Z��          �     ��@   0

           Y�         j���     Z"���    ����              F ����          ��     ��B   (
           9��        ~ g�     9�U i�     U��                ����          �     ��H   8�         ��G          � �[�    ��G �[�                          �         	 ��     ��@   (            {K�        � ��     {wm ��\    �m�                     �         
 �  �  ��A   P
B 
          ���
	      � �)     � �)                              �� U             �  ��@    8		 1                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          :�  ��        ���yc     :�k��{�     U�� "                x                j  �       �                          :    ��        ���       :  ��           "                                                 �                          �    � �� ���  � � �������    	       
      
  =   ��� `%�I       $� �[� %� \� �d 0a� �� b@ �� �c@ �� d@ �D g`���X ���� ����  ����. ����< ����J ����X � (� `r@ )D  s  �� s@ 
�< V� 
�� V� 
�\ W  �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ 
�\ U� 
� V  
�| V ���� � 
�� V� 
�\ W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� �  ���l  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    B�j l �  B �
� �  �  
�  9    ��     �        n��  ��     � �       9    ��     �           � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �H��      �� �T ���        �'T ��        �        ��        �        ��        �  
  ��     ���Xm�        ��                         �$ ( �� �                                    �                  ����            9  ���%��    ��� F�2            �BUF y Yake rson     0:00                                                                        1  1     �C
� �K[ �C.Y � C6i �CJ � C"R �c�a � c�i �	B�E � 
B�U �cV � � c^ � �c� � � c� � �
k� � � k� � � k� � a	� � a	� � q� � q� �"�L "�^ �"�L � *�[ � *�[ �"�L � *�[ �"�L � *�["�M  "�_ �!"�M � *�\ #"�` �$"�N � *�] q&� �'"�O ("�a �)"�O � *�^{+�{ 
�"z 
�!r 
�j 
�g 
�d1� �d 
�_ 
�
 � 
�h � 
�j �6�[ � 
�j � 
�3 �  *K| �  *H| � ;*O| �  *H| �="L � >*O| �  *H|                                                                                                                                                                                                                         d� R `       �     @ 
        �     ] P E h  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��    ��� ��������������������������������������������������������   �4, ?  * ���@S���@�@��A	 ��|���                                                                                                                                                                                                                                                                                                                                z� ��                                                                                                                                                                                                                                         K    -    ��   D�J    	  4�  	                           ������������������������������������������������������                                                                     	                                                                  �      u      u               �  �          	  
 	 
 	 	 ������ �������������  ������������������ ����������� �����  ������� ���� ���������������� ����������� ���������������������� ��������������������������� �������� �� ������� ��� ����������� � �� �������� ����� ����������������� �� �����������������                         	     5          �  L�J                                     ������������������������������������������������������                                                                                                                                             �    ee      �      �          ��                 	 	 � ������������������� ������ ��������� � ���������������  �������������������������� ���� ������ � ����  ������������� ����������������  ��� �������������� ���� ������������������������������������� ������ ���� ��� ������� ��               �                                                                                                                                                                                                                                                                                    
                             �             


             �  }�                                                                                          ������������      ����������������������������  +9����������������������������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 4 H <               	                  � ;�� �\        �t�S$
�C$+TA                                                                                                                                                                                                                                                             )n)n�  E                m      f                              d                                                                                                                                                                                                                                                                                                                                                                                                               > �  	>�  (�  (�  
�  EZm� ��f�A��� =��������d�3��H�,�ɬ� �N ����r�                ����  � u
       	 	 �   &  AG� �   s                    �                                                                                                                                                                                                                                                                                                                                      p B I   j                       !��                                                                                                                                                                                                                            Y��   �� �� �      �� Z 	     ������ �������������  ������������������ ����������� �����  ������� ���� ���������������� ����������� ���������������������� ��������������������������� �������� �� ������� ��� ����������� � �� �������� ����� ����������������� �� ������������������ ������������������� ������ ��������� � ���������������  �������������������������� ���� ������ � ����  ������������� ����������������  ��� �������������� ���� ������������������������������������� ������ ���� ��� ������� ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      @      ,      :                       B     �   �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$ ^h  ��   p   	  ��     �           �� �   6   
���� ���    �����     �    ��������������J JNi   �    ���      $     � ��� �� � ��� �$  � �  �� �  �      �  ��   ����� e�����  g���        f ^�         ��        �      ��Nz���2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "! ""! " ""  "!  "! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "!  " ! " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "! ""! " ""  "!  "! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                          	��ˋ����۪��ۚ{Ƚ�g˽˖�-��"�� .� 
�8 
�� 
D> DC �D0 �D 
�C U@ �� 	�� ��" , " "/ "/� �� �   �                    �   ��  ��  w�  k�� g�� w�� ��� �۹ ��� ��� 3̰ �  >�" 2� 2"�DC �3  ��  ��  +   "   "   "/� ��     �                               �  �� �  �  �   �       �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                             �  �˰ ��� �wp ���                                                                                                                                                                 ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r`ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                            �������  ���    �        � ��                    ���� �                                                                                                                                                                                                      � � ̹ �� �� �� ��� ��� �̻ 9�� EJ� EJ� 4D� 3DJ 4Z 3D �E ɽˠ
� "" �"�"! �"��" ��   �            �  �˰ ̻� ��p �wp ��  ��  ��  ��  ��  �̰ ۻ� ݙ� ݪ� =�� 0�  �   �   �   �   �   �   �   �   �   "   "�    ��  �    �      �   �" �"� "������     �     �� �� ��
��׊��w٪�|��������            "   "   "       �         �        �   �     �       �   �   �   �   �      �                    ��� ���� ��    �     �                                       �   ���                            �   �                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                        � ��                  �  �˰ ��� �wp ���           �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                       �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                /���"/�  ��                    �                                                                            �               �  �  ��  �   �   �         �       �                        �   ��  ���  � �    �                                                                                                                                             �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �      �  �  �  �  �  �   �                                    �   �                                                                                                                                                                                                                        �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��     �   �  �  �  �  �   �                    �� �� �� w� m| ��  �  ��  ��  �   �                     "  ""  """"""
�                               	� ��  �  �  �   �                                                                                                                                                                                            �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �       /   �  �   ��                             �                        ���� ��� ����                      �  �� �� �� ��                         ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                        �          �   � � �  ��� ��  �                    �                        ���� ��� ����                �    ��                 !��� �                                                                                                                                                                                                       �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                {`  g`  w                      �  �  ��"� ��� "                               �                        ���� ��� ����                            �   ���      �  �  �   �   ��  �                            �   ���                            �   �                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��               �   �   �  �  �  �  �   �   �                                       �  ���                    �  �   ��                     �    � �  ��                  ���                              �   ���                            �   �                                                                                                          �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��           �   �                   �  ��  ��  ��  ��� ��� ��� ��˰ɜ˰��˻�̻���������3���DDD�                                                                                                                                                                                                             �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=""""��������AA�A    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ADA�LL��L�D����3333DDDD x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(XxLL����������D����3333DDDD w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""����������A������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(""""�������I�I������ �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�""""�������I��D���I������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`�D�M�D���M������3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(MD�M�A�����MD�����3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(�""""�����AMAD������ � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(�""""������������������ � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(�""""wwwwwwwGGD � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(�""""wwwwwwqwAqwAwA �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(�""""wwwwqwqAwAqAqAq = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=A�A�A�A��LD�����3333DDDD    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( �A�LDL�L�D�L�����3333DDDD x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx""""wwwwwwDGAD w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww""""wwwwqqDAAq  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(""""wwwwwwwGGwGGwGwGw �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((�UQUUQUUQUUQUUUDUUUUU3333DDDD ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`DEQQUUDUTEUUUU3333DDDD M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M""""������������������������ � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(�""""�������DAADAI � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(��A�AM�M�DM��M334CDDDD 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5DD����M��DM�����3333DDDD x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x""""wwwwwwDGqGq w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwwGwwDGwwwwwwww + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+ADAH�DJ�H�H�����3333DDDD � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(��H��J�AD�DH�D����3333DDDD � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(�""""�������DD����� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
� �K[ �C.Y � C6i �CJ � C"R �c�a � c�i �	B�E � 
B�U �cV � � c^ � �c� � � c� � �
k� � � k� � � k� � a	� � a	� � q� � q� �"�L "�^ �"�L � *�[ � *�[ �"�L � *�[ �"�L � *�["�M  "�_ �!"�M � *�\ #"�` �$"�N � *�] q&� �'"�O ("�a �)"�O � *�^{+�{ 
�"z 
�!r 
�j 
�g 
�d1� �d 
�_ 
�
 � 
�h � 
�j �6�[ � 
�j � 
�3 �  *K| �  *H| � ;*O| �  *H| �="L � >*O| �  *H|3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.����������������������������������������� ��=�K�X�X�_��B�G�Q�K� � � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������,�>�0�	�
�������������������� � � � � � �����������������������������������������%��������������������2�0�.� ��!������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            