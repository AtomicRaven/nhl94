GST@�                                                            \     �                                               ��� N     �  ��           ����e ����J�������ĸ��x�������        �g     #    ����                                d8<n    �  ?     h�����  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"    B�j�
�  B ��
  /                                                                               ����������������������������������       ��    =b= 0Q0 44 111  4            	 
                    ��� �� � � ��                 hE 
)         8�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             $F  ")          == �����������������������������������������������������������������������������                                �   ?       �   @  &   �   �                                                                                 '    
)hE  "$)F    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E l �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    �GA�   �Y|$ ~� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V 	  �  �u�GA�   �Y|$ ~� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V 	  �  �r�GA�   �Y|$ ~� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V 	  �  �p�GA�   �Y|$ ~� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V 	  �  �n�GA�   �Y|$ ~� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V 	  �  �l�GA�   �Y|$ ~� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V 
  �  �j�GA�   �Y|$ ~� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V 
  �  �g�GA�   �Y|$ �� @FF� �G  APT0 k� �t�xe1�t B	�1	�"?Q  ��V 
  �  �e�GA�   �Y|$ �� @FF� �G  APT0 k� �h�le1�t B	�1	�"?Q  ��V 
  �  �c�GA�   �Y|$ �� @FF� �G  APT0 k� �X�\e1�t B	�1	�"?Q  ��V 
  �  �`�GA�   �Y|$ �� @FF� �G  APT0 k� �P�Te1�t B	�1	�"?Q  ��V 
  �  �^�GA�   �Y|$ �� @FF� �G  APT0 k� �H�Le1�t B	�1	�"?Q  ��V 
  �  �\�GA�   �Y|$ �� @FF� �G  APT0 k� �@�De1�t B	�1	�"?Q  ��V 
  �  �Z�GA�   �Y|$ �� @FF� �G  APT0 k� �4�8e1�t B	�1	�"?Q  ��V 
  �  �W�GA�   �Y|$ �| @FF� �G  APT0 k� �,�0e1�t B	�1	�"?Q  ��V 
  �  �U�GA�   �Y|$ �t @FF� �G  APT0 k� �$�(e1�t B	�1	�"?Q  ��V 
  �  �S�GA�   �Y|$ �l @FF� �G  APT0 k� �� e1�t B	�1	�"?Q  ��V 
  �  �Q�GA�   �Y|$ �d @FF� �G  APT0 k� � � e1�t B	�1	�"?Q  ��V 
  �  �O�GA�   �Y|$ �\ @FF� �G  APT0 k� � � e1�t B	�1	�"?Q  ��V 
  �  �M�GA�   �Y|$ �T @FF� �G  APT0 k� � � e1�t B	�1	�"?Q  ��V 
  �  �K�GA�   �Y|$ �L @FF� �G  APT0 k� �� �  e1�t B	�1	�"?Q  ��V 
  �  �I�GA�   �Y|$ �D @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V 
  �  �G�GA�   �Y|$ �< @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V 
  �  �F�GA�   �Y|$ �, @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V 
  �  �E�GA�   �Y|$ �$ @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  �D�GA�   �Y|$ � @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  �C�GA�   �Y|$ � @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  �B�GA�   �Y|$ n @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  �A�GA�   �Y|$ n  @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  �@�GA�   �a�$ m� @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  �?�GA�   �a�$ m� @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  �>�GA�   �a�$ m� @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  �=�GA�   �a�$ m� @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  �<�GA�   �a�$ m� @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  �;�GA�   �a�$ m� @FF� �G  APT0 k� �t �x e1�t B	�1	�"?Q  ��V   �  �:�GA�   �a�$ m� @FF� �G  APT0 k� �l �p e1�t B	�1	�"?Q  ��V   �  �9�GA�   �a�$ m� @FF� �G  APT0 k� �d �h e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ m� @FF� �G  APT0 k� �\ �` e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ }� @FF� �G  APT0 k� �X�\e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ }� @FF� �G  APT0 k� �T�Xe1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ }� @FF� �G  APT0 k� �L�Pe1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ }� @FF� �G  APT0 k� �D�He1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ }� @FF� �G  APT0 k� �<�@e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ }| @FF� �G  APT0 k� �4�8e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ }l @FF� �G  APT0 k� �$�(e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ }d @FF� �G  APT0 k� �� e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ }\ @FF� �G  APT0 k� ��e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ }T @FF� �G  APT0 k� ��e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ �L @FF� �G  APT0 k� � �e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ �D @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ �< @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ �4 @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ �(@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ M @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ M@FF� �G  APT0 k� ��	��	e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ M@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ M @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ L�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �a�$ L�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ L�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ L�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ L�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ <�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Y|$ <�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Z�$ <�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Z�$ <�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Z�$ <�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Z�'�<�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �Z�'�<�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �]\'�<�@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �]\'�<�	@FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  �8�GA�   �]\'�<�	@FF� �G  APT0 k� �x�|e1�t B	�1	�"?Q  ��V   �  �8�GA�   �]\'�<|
@FF� �G  APT0 k� �t�xe1�t B	�1	�"?Q  ��V   �  �8�GA�   �]\'�,p@FF� �G  APT0 k� �l�pe1�t B	�1	�"?Q  ��V   �  �8�GA�   �]\'�,l@FF� �G  APT0 k� �l�pe1�t B	�1	�"?Q  ��V   �  �8�GA�   �]\'�,d@FF� �G  APT0 k� �h�le1�t B	�1	�"?Q  ��V   �  �8�GA�   �]\'�,`@FF� �G  APT0 k� �h�le1�t B	�1	�"?Q  ��V   �  �8�GA�   �]l'�,X@FF� �G  APT0 k� �`�de1�t B	�1	�"?Q  ��V   �  �8�GA�   �]l'��T@FF� �G  APT0 k� �d�he1�t B	�1	�"?Q  ��V   �  �8�GA�   �]l'��P@FF� �G  APT0 k� �h �l e1�t B	�1	�"?Q  ��V   �  �8�GA�   �]l'��H@FF� �G  APT0 k� �d!�h!e1�t B	�1	�"?Q  ��V   �  �8�GA�   �]l'��D@FF� �G  APT0 k� �d"�h"e1�t B	�1	�"?Q  ��V   �  �8�GA�   �]l'��@@FF� �G  APT0 k� �d#�h#e1�t B	�1	�"?Q  ��V   �  �8�GA�   �]l'��4@FF� �G  APT0 k� �P �T e1�t B	�1	�"?Q �V   �  �8�GA�   �]l'��0@FF� �G  APT0 k� �D�He1�t B	�1	�"?Q ��_   �  �8�GA�   �]l'��,@FF� �G  APT0 k� �<�@e1�t B	�1	�"?Q ��_   �  �8�GA�   �]l'��(@FF� �G  APT0 k� �0�4e1�t B	�1	�"?Q ��_   �  �8�GA�   �]l'��$@FF� �G  APT0 k� �(�,e1�t B	�1	�"?Q ��_   �  �8�GA�   �]l'��@FF� �G  APT0 k� �� e1�t B	�1	�"?Q ��_   �  �8�GA�   �]l'��@FF� �G  APT0 k� ��e1�t B	�1	�"?Q ��_   �  �8�GA�   �]l'��@FF� �G  APT0 k� ��e1�t B	�1	�"?Q ��_   �  �8�GA�   �]l'��@FF� �G  APT0 k� ��� e1�t B	�1	�"?Q ��_   �  �8�GA�   �]l'��@FF� �G  APT0 k� ����e1�t B	�1	�"?Q	 ��_   �  �8�GA�   �]l'��!@FF� �G  APT0 k� ��#;P e1�t B	�1	�"?Q  �_   �  �8�GA�   �]l'�� "@FF� �G  APT0 k� ��#;P e1�t B	�1	�"?Q�_   �  �8�GA�   �]l'���" FF� �G  APT0 k� ��#;P e1�t B	�1	�"?Q��_   �  �8�GA�   �]l'���# FF� �G  APT0 k� ��#;P e1�t B	�1	�"?Q��_   �  �8�GA�   �]l'���$ FF� �G  APT0 k� ��#;P e1�t B	�1	�"?Q��_   �  �8�GA�   �]l'���% FF� �G  APT0 k� ��#KP e1�t B	�1	�"?Q��_   �  �8�GA�   �]l'���&  F��G  D0T0 k� ��#KP e1�t B	�1	�"?Q��_   �  �8�GA�   �]l'���& ` F��G  D?�T0 k� ��#KP e1�t B	�1	�"?Q��_   �  �8�GA�   �]l'���' ` F��G  D?�T0 k� ��#KP e1�t B	�1	�"?Q��_   �  �8��2A��� � O8# o;�Y| P< �(2��# �+�  3� T0 k� �  � e1�t B	�1�"  ��/ 	  �   2��2A��� � O8# o;�Y| P< �(2��# �+�  3� T0 k� �  � e1�t B	�1�"  /�/ 	  �   4��2A��� � O8# o;�Y| P< �(2��# �+�  3� T0 k� � � e1�t B	�1�"  ��/ 	  �   2��2A��� � O8# o;�Y| �8 �(2��# �+�  3� T0 k� � � e1�t B	�1�"  ��& 	  �   0��2A��� � O8# o;�Y| �0 �(2��# �+�  3� T0 k� � � e1�t B	�1�"  ��& 	  �   .��1A��� � O8# o;�Y| �( �(2��# �+�  3� T0 k� �� �  e1�t B	�1�"  ��& 	  �   ,��1A��� � O8# o;�Y|  �$ �(2��# �+�  3� T0 k� �� �� e1�t B	�1�"  ��& 	  �   *��1A��� o� O8# o7�Y|  � �(2��# �+�  3� T0 k� �� �� e1�t B	�1�"  ��& 	  �   (��1BO�� o� o8#
7�Y|  � �(2��# `+�  3� T0 k� �� �� e1�t B	�1�"  ��& 	  �   &��0BO�� o� o8#
7�Y|$ � �(2@�# `+�  3� T0 k� �� �� e1�t B	�1�"  ��& 	  �   $��0BO�� o� o8#
7�Y|$ � �(2@�# `+�  3� T0 k� �� �� e1�t B	�1�"  ��& 	  �   "��/BO�� o� o8#
3�Y|$ � �(2@�# `+�  3� T0 k� �� �� e1�t B	�1�"  �& 	  �   !��/BO���� o8#
3�Y|( P �(2@�# `+�  3� T0 k� ����e1�t B	�1�"  ��& 	  �    ��.@���� 
4#
3�Y|( P �(2@�#�/�  3� T0 k� ����e1�t B	�1�"  ��& 	  �   ��.@���� 
4#
/�Y|( P �(2 �#�/�  3� T0 k� ����e1�t B	�1�"  ��& 	  �   ��-@���� 
4#
/�Y|( P P(2 �#�/�  3� T0 k� ����e1�t B	�1�"  ��& 	  �   ��,@���� 
0#/+�Y|( P P(2 �#�/�  3� T0 k� ����e1�t B	�1�"  ��& 	  �   ��+@��� 
0#/+�Y|( P  P(2 �#�3�  3� T0 k� ����e1�t B	�1�"  ��& 	  �   ��+@o��� 
,#/'�Y|( P  P(2 �#�3�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��*@o��� 
,#/'�Y|( _� P(2 `�#�3�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��)@o��� 
(#/#�Y|( _�  (2 `�#�7�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��(@o��� 
(#/�Y|( _�  (2 `�# 7�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��'@o��/� 
/$#/�Y|( _�  (2 `�# ;�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��&CO��/� 
/ #/�Y|( _�  $2 `�# ;�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��%CO��/� 
/#/�Y|( _�  $3@�# ?�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��#CO��/� 
/#/�Y|( _� �$3@�$ ?�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��"CO��/� 
/#
O�Y|( _� �$3@�$ C�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��!CO��/� 
/#
O�Y|( _� �$3@�$ G�  3� T0 k� ����e1�t B	�1�"  ��&   �   
�� CO��� #
O�Y|( _� � 4@�$�G�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��CO��� #
O�Y|( _� � 4@�%�K�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��CO��� #
O�Y|( _� � 4@�%�O�  3� T0 k� ����e1�t B	�1�"  ��&   �   ��CO���  #��Y|( _� �5@�&�O�  3� T0 k� ����e1�t B	�1�"  ��&   �   	��CO��� �#���Y|( _� �5@�&�S�  3� T0 k� ����e1�t B	�1�"  ��&   �    	��CO���� �#���Y|( _� �6@�'�S�  3� T0 k� ����e1�t B	�1�"  ��&   �  ��	��C_���� .�#���Y|( _� �6P�(�W�  3� T0 k� ����e1�t B	�1�"  ��&   �  ��	��C_���� .�#���Y|( _� �7P�(�W�  3� T0 k� ����e1�t B	�1�"  ��&   �  ��	��C_���� .�#���Y|( _� �8P�*�_�  3� T0 k� ����e1�t B	�1�"  ��&   �  ��	��C_���� .�#
��Y|( o� �8P�+@_�  3� T0 k� ����e1�t B	�1�"  ��&   �  ��	��C_���� .�#
��Y|( o� �9P�+@c�  3� T0 k� ����e1�t B	�1�"  ��&   �  ��	��C_���� ��"
��Y|( o� �:P�,@c�  3� T0 k� ����e1�t B	�1�"  ��&   �  ��	��C_���� ��"
��Y|( o� �;P�-@g�  3� T0 k� ����e1�t B	�1�"  ��&   �  ���E����� ��"
��Y|( o� �;P�.@g�  3� T0 k� ����e1�t B	�1�"  ��&   �  ���E�ۿ�� ��"���Y|( o� � <P�. k�  3� T0 k� ����e1�t B	�1�"  ��&   �  ���E�۾�� ��"���Y|( o� ��=P�/ o�  3� T0 k� ����e1�t B	�1�"  ��&   �  ���E�ۻ�� ��"���Y|( o� ��?`�0 s�  3� T0 k� ����e1�t B	�1�"  ��&   �  ��o�E�ۺ�� ��"���Y|( o����@`�1 w�  3� T0 k� �� �� e1�t B	�1�"  $�&   �  ��o�E�۸�� ��"���Y|( _����A`�1 w�  3� T0 k� ?� �� e1�t B	�1�"  ��&   �  ��o�E�۷�� 
�!���Y|( _����B`�2 {�  3� T0 k� ?�����e1�t B	�1�"  ��&   �  ��o�E�۵�� 
�!��Y|( _����C`�2��  3� T0 k� ?�����e1�t B	�1�"  ��&   �  ��o�E�۴�� 
�!��Y|( _����D`�2���  3� T0 k� ?�����e1�t B	�1�"  ��&   �  ��o�E�ײ�� 
�!��Y|( _����E0�3���  3� T0 k� ?�����e1�t B	�1�"  ��&   �  ��o�E�װ�� 
�!��Y|( _����F0�3���  3� T0 k� ������e1�t B	�1�"  ��&   �  ��o�E�ׯ�� 
x!��Y|( _����G0�4���  3� T0 k� ������e1�t B	�1�"  ��&   �  ��o�E�׫�� 
h!�Y|( _����I0�5	0��  3� T0 k� ������e1�t B	�1�"  ��&   �  ��o�E�תϘ 
`!w�Y|( �����J �5	0��  3� T0 k� ������e1�t B	�1�"  ��&   �  ��_�E�ӨϘ 
X!o�Y|( �����K �6	0��  3� T0 k� ������e1�t B	�1�"  ��&   �  ��_�E�ӦϘ 
P k�Y|( ���ϼM �6	0��  3� T0 k� ������e1�t B	�1�"  ��&   �  ��_�E�ӤϘ 
H c�Y|( ���ϸN �7	0��  3� T0 k� ������e1�t B	�1�"  ��&   �  ��_�E�ϢϘ 
.@ [�Y|, ���ϴO �7	@��  3� T0 k� ������e1�t B	�1�"  ��&   �  ����E�˟��
., 
K�Y|, ���ϨR0�8	@��  3� T0 k� ������e1�t B	�1�"  ��&   �  ����E�˝��
.$ 
G�Y|0 ���ϤS0�9	@��  3� T0 k� ������e1�t B	�1�"  ��&   �  ����E�Ǜ��
. 
?�Y|0 ���	�T0�9	@��  3� T0 k� ������e1�t B	�1�"  ��&   �  ����
E�Ù��
. 
7�Y|4 ���	�V0�: ��  3� T0 k� ������e1�t B	�1�"  ��&   �  ��_�
E߿�/��
. 
'�Y|8 ���	�X0�: �   3� T0 k� ������e1�t B	�1�"  ��&   �  ��_�
E߻�/��
-� 
�Y|8 ���	�Y0�; �  3� T0 k� ������e1�t B	�1�"  ��&   �  ��_�	E߷�/��
-� 
�Y|< ���	�Z0�; �  3� T0 k� ������e1�t B	�1�"  ��&   �  ��_�	E߳�/��
-�
�Y|< ���	��[0�; �  3� T0 k� ������e1�t B	�1�"  ��&   �  ��_�	E߯�/��
�
�Y|@ ���	��\0�;�  3� T0 k� ������e1�t B	�1�"  ��&   �  ��O�	E߫�/��
�
��Y|@ ���	�|]0�;�  3� T0 k� ������e1�t B	�1�"  ��&   �  ��O�	Eߧ�/��
�
��Y|@ ���	�x^0�;�  3� T0 k� ������e1�t B	�1�"  ��&   �  ��O�	Eߟ���
�
-��Y|D ���	�t_0�;�  3� T0 k� ������e1�t B	�1�"  ��&   �  ��O�	Eߛ���-�
-��Y|D ���	p`0�;�	  3� T0 k� ������e1�t B	�1�"  ��&   �  ��O�	Eߓ���-�
-��Y|D ���	la �;�
  3� T0 k� ������e1�t B	�1�"  ��&   �  ��O�	E��-�
-��Y|H ���	ha �;�  3� T0 k� ������e1�t B	�1�"  ��&   �  ��?�	E��-�
-��Y|H ���	hb �;�  3� T0 k� ������e1�t B	�1�"  ��&   �  ��?�
E���-�
-��Y|H ���	dc �;�  3� T0 k� ������e1�t B	�1�"  ��&   �  ��?�
E�����-�
-��Y|H ���	�dc �;�  3� T0 k� ������e1�t B	�1�"  ��&   �  ��?�
E�{����-�
-��Y|H ���	�`dP�;�  3� T0 k� ������e1�t B	�1�"  �&    �  ��?�E�o����-t
��Y|H ���	�\dP�;��  3� T0 k� ������e1�t B	�1�"  �&    �  ��?�E�g����
Ml
��Y|H ���	�\eP�;��  3� T0 k� ������e1�t B	�1�"  ��&    �  �� ��E�c����
Md
��Y|H ����XeP�;��  3� T0 k� ������e1�t B	�1�"  ��&    �  �� �|E�_����
M\
��Y|H ����Tf��;��  3� T0 k� ������e1�t B	�1�"  �&    �  �� �xE�W����
MT
�Y|H ����Tf��;��  3� T0 k� ������e1�t B	�1�" ��/    �  �� �xE�S����
ML
{�Y|H ����Pg��;��  3� T0 k� �s��w�e1�t B	�1�" ��/    �  �� �tE�O����
MD
s�Y|H ����Lg��;�   3� T0 k� �c��g�e1�t B	�1�" ��/   �  �� �pE�K����
M<
k�Y|H ����Hg��;�  3� T0 k� �O��S�e1�t B	�1�" ��/    �  �� �lA�C����
M4
c�Y|H ����Dh��;�  3� T0 k� �;��?�e1�t B	�1�" ��/    �  �� �hA�?����
M,
_�Y|H ����@h��;�  3� T0 k� �'��+�e1�t B	�1�" ��/    �  �� �hA�;����
M$
W�Y|H ����<h��;�  3� T0 k� ����e1�t B	�1�" ��/   �  �� �dA�7����
M 
O�Y|H ����8h��;�   3� T0 k� ����e1�t B	�1�" ��/    �  �� �`A�3����
M
K�Y|H ����4h��;�(  3� T0 k� ������e1�t B	�1�" ��/    �  �� �\A�/����
M
C�Y|H ����0h�;�,  3� T0 k� ������e1�t B	�1�" ��/    �  �� �\A�'����
M
;�Y|H ����,h�;�4  3� T0 k� ������e1�t B	�1�" ��/    �  �� �XA�#����
M
7�Y|H ����(h�;�8  3� T0 k� ������e1�t B	�1�" ��/    �  �� �TA�����
L�
/�Y|H ����(h�;�@  3� T0 k� ������e1�t B	�1�" ��/    �  �� �TA�����
L�
+�Y|H ����$h�;�H  3� T0 k� ������e1�t B	�1�" ��/    �  �� �PA�� ��
L�
#�Y|H ���� h�;�L   3� T0 k� �{���e1�t B	�1�"	 ��/    �  �� �LA�� ��
L�
�Y|H ����g�;�T!  3� T0 k� �g��k�e1�t B	�1�"	 ��/    �  �� �LA�� ��
L�
�Y|H ����g�;�\"  3� T0 k� �W��[�e1�t B	�1�"	 ��/    �  �� �HA�� ��
L�
�Y|H ���g�;�`#  3� T0 k� �C��G�e1�t B	�1�"
 ��/    �  �� �DA�� ��
L�
�Y|H ���f�;�h%  3� T0 k� �/��3�e1�t B	�1�"
 ��/    �  �� �DA�� ��
L�
�Y|H ���f �;�p&  3� T0 k� ����e1�t B	�1�"
 ��/   �  �� �@A��� ��
L�
�Y|H ���f �;�t'  3� T0 k� ����e1�t B	�1�"
 ��/    �  �� �@A��� ��
L�
��Y|H ���e �;�|(  3� T0 k� ������e1�t B	�1�"
 ��/    �  �� �<A��� ��
L�
��Y|H ���e �;��)  3� T0 k� ������e1�t B	�1�" ��/    �  �� �8A�� ��
L�
��Y|H ��� d �;��+  3� T0 k� ������e1�t B	�1�" ��/    �  �� �8A�� ��
L�
��Y|H ��� d �;��,  3� T0 k� ������e1�t B	�1�" ��/    �  �� �4A�� ��
L�
��Y|H ���~�d x;��-  3� T0 k� ������e1�t B	�1�" ��/    �  �� �4A�� ��
L�
��Y|H P�~�c t;��/  3� T0 k� ������e1�t B	�1�" ��/    �  �� �0A�� ��
L�
��Y|H P�~�c l;��0  3� T0 k� ������e1�t B	�1�" ��/    �  �� �0A�� ��
L�
��Y|H P�~�c h;��2  3� T0 k� �o��s�e1�t B	�1�" ��/    �  �� �,A�ߋ ��
L�
��Y|H P�~�b d;��3  3� T0 k� �[��_�e1�t B	�1�" ��/    �  �� �,A�ߋ ��
L�
��Y|H P�~�b\;��5  3� T0 k� �K��O�e1�t B	�1�" ��/    �  �� �(A�ۋ ��
L�
��Y|H P�~�bX;��6  3� T0 k� �7��;�e1�t B	�1�" ��/   �  �� �(A�׋ ��
L�
��Y|H P�~�aP;��7  3� T0 k� �#��'�e1�t B	�1�" ��/    �  �� �$A�Ӌ ��
L�
��Y|H P���aH<��9  3� T0 k� ����e1�t B	�1�" ��/    �  �� �$A�ό ��
L�
��Y|H P���aD<��;  3� T0 k� ������e1�t B	�1�"
 ��/    �  �� � A�ό ��
L�
��Y|H P���a@<<��<  3� T0 k� ������e1�t B	�1�"
 ��/    �  �� � A�ˌ ��
L|
��Y|H P���`@8<��>  3� T0 k� ������e1�t B	�1�"
 ��/    �  �� �A�ǌ ��
Lx
��Y|H P���`@0<��?  3� T0 k� ������e1�t B	�1�"
 ��/    �  �� �A�Ì ��
Lt
��Y|H P���`@,=��A  3� T0 k� ������e1�t B	�1�"
 ��/    �  �� �A�Í ��
Lp
��Y|H P���_@$=��B  3� T0 k� ������e1�t B	�1�"	 ��/    �  �� �A��� ��
Ll
��Y|H P���_@=��D  3� T0 k� ������e1�t B	�1�"	 ��/    �  �� �A��� �
Lh
��Y|H P���_�>��E  3� T0 k� �w��{�e1�t B	�1�"	 ��/    �  �� �A��� �
Ld
��Y|H P���_�>��G  3� T0 k� �c��g�e1�t B	�1�" ��/    �  �� �A��� �
L`
��Y|H P���^�?��H  3� T0 k� �O��S�e1�t B	�1�" ��/    �  �� �A��� �
L\
��Y|H P���^�?��I  3� T0 k� �?��C�e1�t B	�1�" ��/    �  �� �A��� �
LX
��Y|H P���^��@��K  3� T0 k� �+��/�e1�t B	�1�" ��/    �  �� �A��� �
LT
��Y|H P���]��@��L  3� T0 k� ����e1�t B	�1�" ��/    �  �� �A��� �
LP
��Y|H P���]��A��M  3� T0 k� ����e1�t B	�1�" ��/    �  �� �A��� �
LL
��Y|H P���]��A��O  3� T0 k� ������e1�t B	�1�" ��/    �  �� �A��� �
LH
��Y|H P���]��B��P  3� T0 k� ������e1�t B	�1�" ��/    �  �� �A��� �
LD
��Y|H P���]��B��Q  3� T0 k� ������e1�t B	�1�" ��/    �  �� �A��� �
LD
�Y|H P���\��C��S  3� T0 k� ������e1�t B	�1�" ��/    �  �� �A��� �
L@
�Y|H P���\��C��T  3� T0 k� ������e1�t B	�1�" ��/    �  �� �A��� �
L<
{�Y|H P���\��D��U  3� T0 k� ������e1�t B	�1�" ��/    �  �� �A��� �
L8
w�Y|H P���\��D��V  3� T0 k� �����e1�t B	�1�" ��/    �  �� � A��� �
L4
s�Y|H P���[��E��W  3� T0 k� �k��o�e1�t B	�1�" (�/    �  �� � A��� �
L0
s�Y|H P���[��E��Y  3� T0 k� ;o��s�e1�t B	�1�" ��/    �  �� ��A��� �
L0
o�Y|H P���[��F��Z  3� T0 k� ;s��w�e1�t B	�1�" ��/    �  �� ��A��� �
L,
k�Y|H P#���[��F��[  3� T0 k� ;w��{�e1�t B	�1�" ��/    �  �� ��A��� #�
L(
g�Y|H P#���[��G��\  3� T0 k� ;����e1�t B	�1�"  ��/    �  �� ��A��� #�
L$
g�Y|H P#���Z��G��]  3� T0 k� ;�����e1�t B	�1�"  ��/    �  �� ��A��� #�
L$
c�Y|H P#���Z��H��^  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A��� '�
L 
_�Y|H P#���Z�H��_  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A��� '�
L
_�Y|H P'���Z�I��`  3� T0 k� ������e1�t B	�1�"  /�/    �  �� ��A��� +�
L
[�Y|H P'���Z�I��a  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A��� +�
L
W�Y|H P'���Y�J��b  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A��� +�
L
W�Y|H P'���Y|J��c  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A��� /�
L
S�Y|H P'���YxK��d  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A��� /�
L
O�Y|H P'���YtK�e  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�� /�
L
O�Y|H P+���YpK�f  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�� 3�
L
K�Y|H P+���XhL�g  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�{� 3�
L
K�Y|H P+���XdL�h  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�{� 3�
L
G�Y|H P+���X`M�i  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�{� 7�
L
C�Y|H P+���X\M�j  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�w� 7�
L 
C�Y|H P+�~�XXM�k  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�w� 7�
K�
?�Y|H P+�~�XTN�l  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�s� ;�
K�
?�Y|H P/�~�XPN�l  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�s� ;�
K�
;�Y|H P/�~�WLN�m  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�s� ;�
K�
;�Y|H P/�~�WHO�n  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�o� ;�
K�
7�Y|H P/�~�W@O�o  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�o� ?�
K�
7�Y|H P/��W<O�p  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�k� ?�
K�
3�Y|H P/��W8P�p  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�k� ?�
K�
3�Y|H P/��V4P|q  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�k� C�
K�
/�Y|H P3��V0Pxr  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�g� C�
K�
/�Y|H P3��V0Qps  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�g� C�
K�
+�Y|H P3�~�U,Qls  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�g� C�
K�
+�Y|H P3�~�U(Qdt  3� T0 k� ������e1�t B	�1�"  ��/    �  �� ��A�c� G�
K�
'�Y|H P3�~�U$R`u  3� T0 k� �����e1�t B	�1�"  ��/    �  �� ��A�c� G�
K�
'�Y|H P3�~�T RXv  3� T0 k� ����e1�t B	�1�"  ��/    �  �� ��A�c� G�
K�
#�Y|H P3�~�TRTv  3� T0 k� ����e1�t B	�1�"  ��/    �  �� ��A�_� G�
K�
#�Y|H P3�~�TSLw  3� T0 k� ����e1�t B	�1�"  ��/    �  �� ��A�_� K�
K�
�Y|H P7�~�TS�Dx  3� T0 k� ����e1�t B	�1�"  ��/    �  �� ��A�_� K�
K�
�Y|H P7�~�SS�@x  3� T0 k� ����e1�t B	�1�"  ��/    �  �� ��A�_� K�
K�
�Y|H P7�~�SS�8y  3� T0 k� ����e1�t B	�1�"  ��/    �  �� ��A�[� K�
K�
�Y|H P7�~�ST�0z  3� T0 k� ���#�e1�t B	�1�"  ��/    �  �� ��A�[� O�
K�
�Y|H P7�~�RT�,z  3� T0 k� �#��'�e1�t B	�1�"  ��/    �  �� ��A�[� O�
K�
�Y|H P7�~�RT�${  3� T0 k� �'��+�e1�t B	�1�"  ��/    �  �� ��A�W� O�
K�
�Y|H P7�~�R U�{  3� T0 k� �/��3�e1�t B	�1�"  ��/    �  �� ��A�W� O�
K�
�Y|H P7�~�R U�|  3� T0 k� �?��C�e1�t B	�1�"  ��D    �  �� ��A�W� O�
K�
�Y|H P7���Q�U�}  3� T0 k� �C��G�e1�t B	�1�"  ��D    �  �� ��A�W� S�
K�
�Y|H ;���Q�U�}  3� T0 k� �G��K�e1�t B	�1�"  ��D    �  �� ��A�S� S�
K�
�Y|H ;���Q�V� ~  3� T0 k� �K��O�e1�t B	�1�"  ��D    �  �� ��A�S� S�
K�
�a�H ;���Q�V��~  "�� T0 k� �K��O�e1�t B	�1�"  ��D    �  �� ��A�S� S�
K�
�a�H ;���P��V��  "�� T0 k� �O��S�e1�t B	�1�"  ��D    �  �� ��A�S� S�
K�
�a�H ;���P��V��  "�� T0 k� �K��O�e1�t B	�1�"  ��D    �  �� ��A�O� W�
K�
�a�H ;���P��W���  "�� T0 k� �K��O�e1�t B	�1�"  ��D    �  �� ��A�O� W�
K�
�a�H ;���P��W�؀  "�� T0 k� �K��O�e1�t B	�1�"  ��D    �  �� ��A�O� W�
K�
�a�H ;���O��W��  "�� T0 k� �G��K�e1�t B	�1�"  ��D    �  �� ��A�O� W�
K�
�a�H ;���O��W��  "�� T0 k� �G��K�e1�t B	�1�"  ��D    �  �� ��A�K� W�
K�
�a�H ;���O��W�  "�� T0 k� �G��K�e1�t B	�1�"  ��D    �  �� ��A�K� [�
K�
�a�H  ?���O��X�  "�� T0 k� �C��G�e1�t B	�1�"  ��D    �  �� ��A�K� [�
K�
�a�H  ?���O��X�~  "�� T0 k� �C��G�e1�t B	�1�"  ��D    �  �� ��A�K� [�
K�
�a�H  ?���N��X�~  "�� T0 k� �C��G�e1�t B	�1�"  ��D    �  �� �� A�K� [�
K�
��Y|H  ?���N��Y�~  3� T0 k� �C��G�e1�t B	�1�"  ��D    �  �� �� A�G� [�
K�
��Y|H  ?���N��Y�~  3� T0 k� �?��C�e1�t B	�1�"  ��D    �  �� �� A�G� [�
K�
��Y|H  ?���N��Z�~  3� T0 k� �?��C�e1�t B	�1�"  ��D    �  �� �� A�G� _�
K�
��Y|H  ?���NN�Z�}  3� T0 k� �?��C�e1�t B	�1�"  ��D    �  �� �� A�G� _�
K�
��Y|H  ?���MN�[�}  3� T0 k� �;��?�e1�t B	�1�"  ��D    �  �� �� A�G� _�
K�
��Y|H  ?���MN�[|}  3� T0 k� �;��?�e1�t B	�1�"  ��D    �  �� �� A�C� _�
K�
��Y|H ?���MN�\t}  3� T0 k� �;��?�e1�t B	�1�"  ��D    �  �� �� A�C� _�
K�
��Y|H ?���MN�\l}  3� T0 k� �;��?�e1�t B	�1�"  ��D    �  �� �� A�C� _�
K�
��Y|H ?���MN�]d|  3� T0 k� �7��;�e1�t B	�1�"  ��D    �  �� �� A�C� c�
K�
��Y|H ?���LN�^`|  3� T0 k� �7��;�e1�t B	�1�"  ��D    �  �� �� A�C� c�
K�
��Y|H C���L>�^ X|  3� T0 k� �7��;�e1�t B	�1�"  ��D    �  �� �� A�?� c�
K�
��a�H C���L>�_ P|  "s� T0 k� �3��7�e1�t B	�1�"  ��D    �  �� �� A�?� c�
K�
��a�H C���L>�` L|  "s� T0 k� �3��7�e1�t B	�1�"  ��D    �  �� �� A�?� c�
K�
��a�H C���L>�a D{  "s� T0 k� �3��7�e1�t B	�1�"  ��D    �  �� �� A�?� c�
K�
��a�H C���L>�b @{  "s� T0 k� �3��7�e1�t B	�1�"  ��D    �  �� �� A�?� c�
K�
��a�H PC���K>�c 8{  "s� T0 k� �/��3�e1�t B	�1�"  ��D    �  �� �� A�?� g�
K�
��a�H PC���K>�d 4{  "s� T0 k� �/��3�e1�t B	�1�"  ��D    �  �� ��!A�;� g�
K� 
��a�H PC���K>�e ,{  "s� T0 k� �/��3�e1�t B	�1�"  ��D    �  �� ��!A�;� g�
K� 
��a�H PC���K>�f (z  "s� T0 k� �/��3�e1�t B	�1�"  ��D    �  �� ��!A�;� g�
K� 
��a�H PC���K>�g $z  "s� T0 k� �/��3�e1�t B	�1�"  ��D    �  �� ��!A�;� g�
K� 
��a�H PC���K>�h z  "s� T0 k� �+��/�e1�t B	�1�"  ��D    �  �� ��!A�;� g�
K� 
��a�H PC���J.�i z  "s� T0 k� �+��/�e1�t B	�1�"  ��D    �  �� ��!A�;� g�
K�!
��Y|H PC���J.�j z  3� T0 k� �+��/�e1�t B	�1�"  ��D    �  �� ��!A�;� k�
K�!
��Y|H PC���J.�k z  3� T0 k� �+��/�e1�t B	�1�"  ��D    �  �� ��!A�7� k�
K�!
��Y|H PG���J.�l y  3� T0 k� �'��+�e1�t B	�1�"  ��D    �  �� ��!A�7� k�
K�!
��Y|H PG���J.|n  y  3� T0 k� �'��+�e1�t B	�1�"  ��D    �  �� ��!A�7� k�
K�!
��Y|H PG���J.xo/�y  3� T0 k� �'��+�e1�t B	�1�"  ��D    �  �� ��!A�7� k�
K�"
��Y|H PG�~�J.tq/�y  3� T0 k� �'��+�e1�t B	�1�"  ��D    �  �� ��!A�7� k�
K�"
��Y|H PG�~�I.ts/�y  3� T0 k� �#��'�e1�t B	�1�"  ��D   �  �� ��!A�7� k�
K�"
��Y|H PG�~�I.tt/�y  3� T0 k� �#��'�e1�t B	�1�"  ��D    �  �� ��!A�3� k�
K�"
��Y|H PG�~�I.pu/�x  3� T0 k� �#��'�e1�t B	�1�"  ��D    �  �� ��!A�3� o�
K�"
��Y|H PG�~�Ipw/�x  3� T0 k� �#��'�e1�t B	�1�"  ��D    �  �� ��!A�3� o�
K�"
��Y|H PG� �Ipx/�x  3� T0 k� �#��'�e1�t B	�1�"  ��D    �  �� ��!A�3� o�
K�#
��Y|H PG� �Ipy/�x  3� T0 k� �#��'�e1�t B	�1�"  ��D    �  �� ��!A�3� o�
K�#
��Y|H PG� �Ip{/�x  3� T0 k� ���#�e1�t B	�1�"  ��D    �  �� ��!A�3� o�
K�#
��Y|H PG� �Ip|/�x  3� T0 k� ���#�e1�t B	�1�"  ��D    �  �� ��!A�3� o�
K�#
��Y|H PG� �Hp}/�x  3� T0 k� ���#�e1�t B	�1�"  ��D    �  �� ��!A�3� o�
K�#
��Y|H PG���Hp~/�x  3� T0 k� ���#�e1�t B	�1�"  ��D    �  �� ��"A�/� o�
K�#
��Y|H PG���Hp/�w  3� T0 k� ���#�e1�t B	�1�"  ��D    �  �� ��"A�/� o�
K�$
��Y|H PG���Hp�/�w  3� T0 k� ���#�e1�t B	�1�"  ��D   �  �� ��"A�/� o�
K�$
��Y|H PG���Hp�/�w  3� T0 k� ����e1�t B	�1�"  ��D    �  �� ��"A�/� s�
K�$
��Y|H PK���H�p�/�w  3� T0 k� ����e1�t B	�1�"  ��D    �  �� ��"A�/� s�
K�$
��Y|H PK���H�t�/�w  3� T0 k� ����e1�t B	�1�"  ��D    �  �� ��"A�/� s�
K�$
��Y|H PK���H�t/�w  3� T0 k� ����e1�t B	�1�"  ��D    �  �� ��"A�/� s�
K�$
��Y|H PK���H�t/�w  3� T0 k� ����e1�t B	�1�"  ��D    �  �� ��"A�/� s�
K�$
��Y|H PK���G�t/�w  3� T0 k� ����e1�t B	�1�"  ��D    �  �� ��"A�/� s�
K�%
��Y|H PK���G�t/�v  3� T0 k� ����e1�t B	�1�"  ��D    �  �� ��"A�/� s�
K�%
��Y|H PK���G�x~/�v  3� T0 k� ����e1�t B	�1�"  ��D    �  �� ��"A�+� s�
K�%
��Y|H PK���G�x~/�v  3� T0 k� ����e1�t B	�1�"  ��D    �  �� ��"A�+� s�
K�%
��Y|H PK���G�x~/�v  3� T0 k� ����e1�t B	�1�"  ��D    �  �� ��"A�+� s�
K�%
��Y|H PK���G�x~�v  3� T0 k� ����e1�t B	�1�"  ��D    �  ��\XA�Ǣp[�tY �tZ�� �L rO�� �H  A_�T0 k� �<b�@be1�t B�1	�"?Q  ��7   � <�8\XA�Ǣp\�xX �tZ�� �L$rO�� �L  A_�T0 k� �<b�@be1�t B�1	�"?Q  ��7   � <�8\YA�Ǣl\�|X �tb�� �L$rO�� �L  A_�T0 k� �@b�Dbe1�t B�1	�"?Q  ��7   � <�8\YA�Ǣl\��X �tb�� �L$rO�� �P  A_�T0 k� �@b�Dbe1�t B�1	�"?Q  ��7   � <�8\YA�Ǣl]��X �tb�� �L$rO�� �P  A_�T0 k� �@b�Dbe1�t B�1	�"?Q  ��7   � <�8\YA�Ǣl]��W �tb�� �L$rO�� �T  A_�T0 k� �@b�Dbe1�t B�1	�"?Q  ��7   � <�8\ZA�Ǣl^��W �tb�� �L$rO�� �T  A_߳T0 k� �@a�Dae1�t B�1	�"?Q  ��7   � <�8\ZA�Ǣl^��W �tb�� �L(rO�� �T  A_߳T0 k� �@a�Dae1�t B�1	�"?Q  ��7   � <�8\ZA�Ǣl^��W �tb�� �L(rO�� �X  A_߳T0 k� �Da�Hae1�t B�1	�"?Q  ��7   � <�8\ZA�Ǣl_��V �tb�� �L(rO�� �X  A_۳T0 k� �Da�Hae1�t B�1	�"?Q  ��7   � <�8\[A�Ǣl_��V �tb�� �L(rO�� �X  A_۳T0 k� �Da�Hae1�t B�1	�"?Q  ��7   � <�8\[A�Ǣl`��V �tb�� �L(rO�� �\  A_۴T0 k� �Da�Hae1�t B�1	�"?Q  ��7   � <�8\ [A�Ǣl`��V �tb�� �L(rO�� �\  A_״T0 k� �Da�Hae1�t B�1	�"?Q  ��7   � <�8\ [A�Ǣl`��U �tZ�� ��(rO�� �`  A_״T0 k� �@`�D`e1�t B�1	�"?Q  ��7   � <�8\ [A�Ǣla��U �tZ�� ��,rO�� �`  A_ӴT0 k� �<`�@`e1�t B�1	�"?Q  ��7   � <�8\ \A�Ǣla��U �tZ�� ��,rO�� �`  A_ӴT0 k� �<`�@`e1�t B�1	�"?Q  ��7   � <�8\ \A�Ǣla��U �tZ�� ��,rO�� �d  A_ӴT0 k� �<`�@`e1�t B�1	�"?Q  ��7   � <�8\ \A�Ǣlb��U �tZ�� ��,rO�� �d  A_ϴT0 k� �<`�@`e1�t B�1	�"?Q  ��7   � <�8\ \A�Ǣhb��T �tZ�� ��,rO�� �d  A_ϵT0 k� �<`�@`e1�t B�1	�"?Q  ��7   � <�8\ \A�Ǣhb �T �tZ�� ��,rO�� �h  A_ϵT0 k� �<`�@`e1�t B�1	�"?Q  ��   � <�8\ ]A�Ǣhc �T �tZ�� ��,qO�� �h  A_˵T0 k� �<_�@_e1�t B�1	�"?Q  ��   � <�8\ ]A�Ǣhc �T �tZ�� ��,q@� �h  A_˵T0 k� �<_�@_e1�t B�1	�"?Q  ��   � <�8\ ]A�Ǣhc �S �tZ�� ��0q@� �h  A_˵T0 k� �@_�D_e1�t B�1	�"?Q  ��   � <�8\ ]A�Ǣhd �S �tZ�� ��0q@� �l  A_ǵT0 k� �@_�D_e1�t B�1	�"?Q  ��   � <�8\ ]A�Ǣhd �S �tZ�� �	0q@� �l  A_ǶT0 k� �@_�D_e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhd S �tZ�� �	0q@� �l  A_ǶT0 k� �@_�D_e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhe S �tZ�� �	0q@� �p  A_ǶT0 k� �@_�D_e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhe S �tZ�� �	0q@#� �p  A_öT0 k� �@_�D_e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhe R �tZ�� �	0q@+� �p  A_öT0 k� �@_�D_e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhe R �tZ�� �	0q@/� �t  A_öT0 k� �@_�D_e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhf  R �tZ�� �	0q@3� �t  A_��T0 k� �@_�D_e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhf $R �tZ�� �	4q@7� �t  A_��T0 k� �D_�H_e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhf (R �tZ�� �	4q@?� �t  A_��T0 k� �D_�H_e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhg 0Q �tZ�� �	4q@C� �x  A_��T0 k� �D_�H_e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhg 4Q �tZ�� ��4q@G� �x  A_��T0 k� �D^�H^e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhg 8Q �tZ�� ��4q@K� �x  A_��T0 k� �D^�H^e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhg <Q �tZ�� ��4q@S� �x  A_��T0 k� �D^�H^e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhh DQ �tZ�� ��4q@W� �|  A_��T0 k� �D^�H^e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣhh HQ �tZ�� ��4q@[� �|  A_��T0 k� �D^�H^e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣdh LQ �tZ�� ��4q@_� �|  A_��T0 k� �D^�H^e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣdh PP �tZ�� ��4q@g� �|	  A_��T0 k� �D^�H^e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣdh TP �tZ�� ��8q@k� ��	  A_��T0 k� �H^�L^e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣdi \P �tZ�� ��8q@o� ��	  A_��T0 k� �H^�L^e1�t B�1	�"?Q  ��   � <�8� ]A�Ǣdi `P �tZ�� ��8q@s� ��	  A_��T0 k� �DZ�HZe1�t B�1	�"?Q  �   � <�8� ]A�Ǣdi dP �tZ�� ��8q@{� ��	  A_��T0 k� �@W�DWe1�t B�1	�"?Q ��   � <�8� ]A�Ǣdi hP �tZ�� ��8q@� ��	  A_��T0 k� �8S�<Se1�t B�1	�"?Q ��   � <�8� ]A�Ǣdj lP �tZ��  �8q@�� ��	  A_��T0 k� �4O�8Oe1�t B�1	�"?Q ��   � <�8� ]A�Ǣdj pO �tZ��  �8q@�� ��	  A_��T0 k� �0K�4Ke1�t B�1	�"?Q ��   � <�8� ]A�Ǣdj tO �tZ��  �8q@�� ��	  A_��T0 k� �,H�0He1�t B�1	�"?Q ��   � <�8� ]A�Ǣdj xO �tZ��  �8q@�� ��	  A_��T0 k� �(D�,De1�t B�1	�"?Q ��   � <�8� ]A�Ǣdj |O �tZ��  �8q@�� ��	  A_��T0 k� �$@�(@e1�t B�1	�"?Q ��   � <�8� ]A�Ǣdk �O �tZ��  �8q@�� ��	  A_��T0 k� � <�$<e1�t B�1	�"?Q ��   � <�8� ]A�Ǣdk �O �tZ��  �<q@�� ��	  A_��T0 k� �8� 8e1�t B�1	�"?Q ��   � <�8� ]A�Ǣdk �O �tZ��  �<q@�� ��	  A_��T0 k� �5�5e1�t B�1	�"?Q ��   � <�8� ]A�Ǣdk �O �tZ��  �<q@�� ��	  A_��T0 k� �1�1e1�t B�1	�"?Q ��   � <�8� ]A�Ǣdk �N �tZ��  �<q@�� ��	  A_��T0 k� �-�-e1�t B�1	�"?Q ��   � <�8�GA�   �Y|  `@ @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|  `@ @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|  `@ @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|  `< @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|  `< @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|  `8 @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|  `8 @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|  `4 @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|  `4 @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ `0 @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ p, @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ p( @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ p$ @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ p$ @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ p  @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ p @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ p @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ p @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ p @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ � @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �  @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �|��e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �t �x e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �p �t e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �h �l e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �d �h e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �\ �` e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �T �X e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �L �P e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �H �L e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �@ �D e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �8 �< e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ �� @FF� �G  APT0 k� �0 �4 e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ o| @FF� �G  APT0 k� �( �, e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ ot @FF� �G  APT0 k� �  �$ e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ ol @FF� �G  APT0 k� � � e1�t B	�1	�"?Q  ��V   �  ���GA�   �Y|$ o\ @FF� �G  APT0 k� � � e1�t B	�1	�"?Q  ��V 	  �  ���GA�   �Y|$ oT @FF� �G  APT0 k� �  � e1�t B	�1	�"?Q  ��V 	  �  ���GA�   �Y|$ oL @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V 	  �  ���GA�   �Y|$ oD @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V 	  �  ���GA�   �Y|$ o< @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V 	  �  ���GA�   �Y|$ o4 @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V 	  �  ���GA�   �Y|$ o, @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V 	  �  ���GA�   �Y|$ o$ @FF� �G  APT0 k� �� �� e1�t B	�1	�"?Q  ��V 	  �  �~�GA�   �Y|$  @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V 	  �  �|�GA�   �Y|$  @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V 	  �  �z�GA�   �Y|$  @FF� �G  APT0 k� ����e1�t B	�1	�"?Q  ��V 	  �  �x                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \���� ]�.. � � "{�          ���I�     "r���X)     ��'                �          �     ���   0

 	 	         ��*    	     �����    ��!f���b     ���                  �         �0     ���   (	          ��t             ݡ    ��t �P      A            � �         ��  �  ���   8�

          %��   � �
     ��Z�     %l���^6    ���                 �$          `
`     ���   (	          ����   � �        .��s    �������H    ����               ���$           p
`      ���   P
	B           � ��       B�<�      ��<�                              ���                �  ���    8		 1 	            �ɘ>    	   V i�    �ɣ3 ^�    �[ �             Z��         ��     ��H   8	           G��  + +      j���     G�����c    ���               Z��          O��  �  ��@  0	
		 	          ~#�  � �
     ~����     ~b.����    �S�              v	 Z��           �     ��`  0 
           v�  � � 
	   ���b�     v����@    �|��              B Z��         	 ���    ��` @
(         �!a        �  �q    �!a  �q               ��       	 � !         
 �        ��F   H	           l0 � �     � �1"      l0 �1"                            Z���             �  ��@    8

 '                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         �úa  ��        ��a�    �ú���;    ���� "                x                j  �       �                         ��    ��        ��      ��  �           "                                                �                         ���� ����� ������   ����� 	         
       
  �    v0> ���G       �D �r@ �� s� �d  q  ��  n� �� �r@ �� s@ � s` �$ s� �D s� �d s� � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0� ���� ����� � 
�| V  
�\ W� 
�� W� 
�| W����� � �$ a� �D @a� ��  w@ �� �w� �d  x� �$  }` �d  }����� � C� `t� Dd u� D� u� D� u� C� `^@ Dd _  D� _  D� _@  �o� >D ``� ? @a� ?� b  
�< U� 
� V  
� V  
�\ W� 
�� W� 
�| W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������  �� /  ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"    B�j
��  B �
� �  �  
� ��    ��     ���      ��    ��     ���      ����  ��     �           � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �DBB	      �� �T ��        �bT ���        �        ��        �        ��        �   �    �h���� e        ��                         �$ ( � �����                                     �                 ����            �������%��    ����                �BUF e Duchesne y    0:00                                                                        6  6      �C
2� � J� �8 J� �	c~sc�u �c�u �cj@ cr8 �	B� 
B�/ �c�j � c�r � c�e � c�h � c�n � c�p �cV � � c^ � �C � �"� � � "� � �� � � 
� � � 
� � � 
� � �� � � 
� � � 
� � � "� � �� � � 
� � � 
� � � 
� � � ""� � �#� � � 
� � � 
� � �&� � � 
� � �(� � � 
� � �*� � � 
� �,*l-)�t8 .*DL0/*
lP 0*CTX 1*G\X  *K<X  *K<X  *K<5*<d6*2t07*6t8 8*DLP 9*RTX :*K\X  *K<)  "@ |R  "J z � >*Kx  )�x                                                                                                                                                                                                                         \� P              @        �     W P E c  ���� S               �������������������������������������� ���������	�
��������                                                                                          ��    ��� '  ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, E� < !��� J��@�@��@ڃ�@����.��K������(���                                                                                                                                                                                                                                                                                                               �@@����                                                                                                                                                                                                                                  [  	  &    ��  L�J                                     ������������������������������������������������������                                                                       
                                                           	      �    �              �          �< J              	 	 ���  ���������������� ��������������������  ����� ������� ��������������� ��������������� ������  ���� ��������������������������� ��������� ��� � ������������ ��� ����� ���  ���������� ���� ��� ����� �� ������� ��� � ���������������������           3           
        .    ��  9<�J     ��  	                           ������������������������������������������������������                                                                                                                                     �  ��                  V     �BD                   � ������������������������������������������������������������� ��������� ������������ ����� ��������� ������������������� � ��� ������� ������� ������������������ ��������� �� � ���� ������ ����������� ������ ����������  ����������� �                                                                                                                                                                                                                                                                                                                      �             


           �   }�         ������������  R~��������������������������������    ��������������������  '�����������������������������        R�                                 R�                                     �ww�ww333wwwwwwww�ww�ww�ww�ww333wwww I @ 5 
                                � (�� �\                                                                                                                                                                                                                                                                                    
)hE  "$)F                l               W                   `                                      ��                                                                                                                                                                                                                                                                                                                                      j                               @ D  � ��  � ��  � #��  � #��  J`D  ���������}�����������������M���������������d        6   w � : 	 |	          �   & AG� �   �              �4�                                                                                                                                                                                                                                                                                                                                  p I G   �      ��  #             !��                                                                                                                                                                                                                            Y   �� �~ ���      �� 3      ���  ���������������� ��������������������  ����� ������� ��������������� ��������������� ������  ���� ��������������������������� ��������� ��� � ������������ ��� ����� ���  ���������� ���� ��� ����� �� ������� ��� � ���������������������� ������������������������������������������������������������� ��������� ������������ ����� ��������� ������������������� � ��� ������� ������� ������������������ ��������� �� � ���� ������ ����������� ������ ����������  ����������� �     �     $�l�������l����������������������l��������������f���f���f��ff���f������ffffflffffffffffffffffffff����ff��lfflffffffffffffffffffffl��l��̼���l����l��lf���ll��������l�����ll������l�����������������l���������������l��������������fff�lff�ll��l���li��f���l���f��ffffffffffff��������������������fffffff�ffl��̻�����������������f�l���l�llll�l�̦ll̜f�̊�l̊���l����������������������������������������������������������������f���f���f���f���f���f��ɜ�����������������������̺��ƹ��li��fiy��������������˩�ff��fl��fk��fj���f̈�f̈�f̈�f̈�fl�{ʜ�����������l����������������̼��������������������������������������̼̼��������j���ˊ��̗��̸���ʈ���Ɉ��i���������������������������y��fj���k���̨��̹��l���̹��lɹ��ʘ�����ɬ��ȼ�������l���̘��̈���������̼����̼������̼�����̼��������������̼���������̼���̼̼���k�̼̈��̈��ˈ��˘̼����˘��̘�Ɉ����������������ˈ�����������k��ɫ��ɫ����ff��ɶ��ɻ�ll���������̉��ˈ��̈��̙��ˈ�̼���l�����������������̼����˼�̶���̻�������������˨̩��������������������ʈ����������|����i����Ʒi��i��������������������������j���f��������̹�̼���̘�fʘ��ɉ����̊�̼��ȸ�{�Ɉ��h�����l���j���h��fȹ����̈xx�������������f���l��l�������    1      >   � ��                       4     �   ���������J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��     �� p���� ���� p���� �$��   `d     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@       �      �     ��     3� � ��� �� � ��� � �2v �2��v  �      �  ��   ���� e�����  g���        f ^�         �� �              ���8���2�������J��e���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 " ""   "" "!  "" "  """ !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                   " ""   "" "!  "" "  """ !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                        "!  "! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                      �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                             �� ��������p��}`     �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                                    � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                   �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                      �  ������� ��       �  �  �   �   ��  �                            �   ���                            �   �                                                                                                    �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �    �   ��  �  ��  �             �  �   �   ��  �                �   �   �   �      �  �                         �  ���               �������  ���    �                    ��  ��  ���  �  �  �   �   ��  �                            �   ���                            �   �                                                                                                        �   �   �   � 
�w ��� ș����	���
���	������ ݼ� ݼ� �� �� 	�� �� 3E 34 D@ ��  ��  ʢ  ""� "/  ��� �      �    �   ��  ��  �p  �p  w   ��  ��� ��� ��� ˻� ̼˰��ː�۹�̽��̽����˸� "��@ DJ� EZ� DU� EZ  DL̘ 	�������" �""�"/��"� ��                    � ��� "  �         �    �  �       �   �   ��  �   �   �   �           �   �       ��  � �                    ��  ��  ��                          ��  ��  ���                                                                                                                                                                                                       �   �   �   �   w  �� ɪ�̚��ə���̚���ɭ�̼��̻��̻���+���(�� H� �C3 UC3
TDCTD0�C 	�� 
�� ���� ���"/� ��   ���   ��  ��  ��  w�  wp  ��� ��� ��̰��̀�͹���ڀ��ذ��� �̰ �̰ ̸� ��� ��3 333�3330�C3: TD3�C��ݸ�	��  ����̲����"/����     � �  �  ��  �  �   �   �      	  *  ,  +   "   ��   �   ��  �   �   �   �                             ��  ��  �          ��                           � ��                    ���� �                                                                                                                                                                                                          �� �����ݼڜ��ک��ک��z�	��� 
�� 
�� 	�� ̘ ɪ  ��  �  �� �� ������������ ���  � � � �� �� ������ ��                      �   ��  ��  �̰ ��� ��˰�̻��̻���������ˉ�U��EP�ET �I� ٕ  �D� �L� ��� ��" ����/�"�"�""�����                             �   �   �   �   z�  ��  ��  ���������  ��  ̿� ��� ��  ��� ��  ���  �  � �                     ��� ����                                �   �                                                                                                                                                                                                                	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  �   �   �   �   �       �     �"  "  �   "                                    �   �   �            �� �� �� g} �� vw                     �    � �  ��                  ���                              �   ���                            �   �                                                                                                        �   �   �   �  
� 	�� �� ���	���
���	������+�ݼ� �  
C  �U  �T 
UC 
UT ED  �D  ��  �  �   " �"  �     �        �   ��  ��  ��  w�  ��  ��� ��� ̻� ̻���˩�̽��̽� ˉ� ��  340 UT0 DD0 330 33  C  C  
�  �  ,�  ""  "  �� ��     �      �   ��  �  ��  �             �  �   �   ��  �                         �                             ���                         �  ��                    �����                                  �  �˰ ��� �wp ���                    �   ���                            �   �    ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                             "  "(��ȩ�ܚ��ۊ����� ��  �   �   �   �   �� ��� ̻� ˽� ��� �w� �������������������������� �̻ ���         �   �       �   �   "" �+� Ȼ� ɫ� ɨ� ��                �� �I��3 ��D 
UD 
UD TD  T�  ˸  ��  �� ̰ �+ ��"/ �"/  ����  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �         �                                           � ��                  �  �˰ ��� �wp ���                                                                                                                                                                      �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��                     �    � �  ��                  ���                                                                                                                                                                           ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r`     �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����        �   �  ���� �   �             �   ��  ��  ��  �  �   ��  ��                                                                                                                                                                 "  " �" ��" ��- �ۼ w۽��ݹ����� ��� ��  ˼  ��  ˼  ��  H�  �D  J�  J�  �  �  �  �  
�  �  �  �  ,�  " "" �" �"�   ˰  ��  wp ��ډ�v���r�̸��˰��� ��  ��  ��  ��  ̸  ��  ��  DC  C4@ T4@ T40 T30 T30 S;� H�  ��  ��  ��  ""  "  �""� "�/��        �   �   �      �  �   �   �   �   �              �   �   �   �             ���� �                        " "" """ �"  �   �   �                              � ��                  �  �˰ ��� �wp ���                                                                                                                                                                             �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""������������������""""������������������������""""������������������������""""������ADAIA�A""""�������I�A�A�A""""�����DD�I""""�������DAADAI""""������IDA��""""��������DD��I�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD������������������������3333DDDD�A�AM�M�DM��M334CDDDD�A�AM�M�DDM����3333DDDDDM����DD�����3333DDDDMAM��D�DDM�����3333DDDDDD����M��DM�����3333DDDD������������DD������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
2� � J� �8 J� �	c~sc�u �c�u �cj@	 cr8 �	B� 
B�/ �c�m � c�} � c�e � c�h � c�n � c�p �cV � � c^ � �C � �"� � � "� � �� � � 
� � � 
� � � 
� � �� � � 
� � � 
� � � "� � �� � � 
� � � 
� � � 
� � � ""� � �#� � � 
� � � 
� � �&� � � 
� � �(� � � 
� � �*� � � 
� �,*l-)�t8 .*DL0/*
lP 0*CTX 1*G\X  *K<X  *K<X  *K<5*<d6*2t07*6t8 8*DLP 9*RTX :*K\X  *K<)  "@ |R  "J z � >*Kx  )�x3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������$��7�O�Q�K��;�O�I�I�O� � � � � � � � � � �:�>�/����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0�����������������������������������������#��<�Z�K�\�K��.�[�I�N�K�Y�T�K� � � � � � �:�>�/�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������:�>�/� ��!�������������������������������������,�>�0�	�
�������������������� � � � � � �����������������������������������������%��������������������,�>�0� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $������������������������     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %������������������������ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                