GST@�                                                            \     �                                               7���      �     )         �������J���J�����������x�������        i      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    
 �j,� B ��
  4�                                                                              ����������������������������������      ��    bb= QQ0 4 111 44              		 

                     ��� �   � �                 nn ))
         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                   +       �   @  &   �   �                                                                                 '     )n)n
  �    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE + �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    @w� �@c\9@�AM�|(B��L���L� JD�0,sw�3�T0 k� ��� %�0e  51D Q  ��    � 
 �@w� �@c`9@�AM�|(B��L���L� KD�0-sw�3�T0 k� ����%�0e  51D Q  ��    � 
 �@{� ��@c`9@�AM�|(B��L���L�LD�0.s{�3�T0 k� ����%�0e  51D Q  ��    � 
 �@{� ��@cd9@�AM�|(B��L���L�LD�0/s�3�T0 k� ����%�0e  51D Q  ��    � 
 �@{� ��@cd9@�AM�|(���L���L�MD�0/s�3�T0 k� ����%�0e  51D Q  ��    � 
 �@� ��@ch:@�AM�|(���L���L�ND�00s��3�T0 k� ����%�0e  51D Q  ��    � 
 �@� ��@cl:@�AM�|(��L���L�OD�01s��3�T0 k� ��	��	%�0e  51D Q  ��    � 
 �@� ��@cl:@�AM�|(��L���L�PD�02s��3�T0 k� ��	��	%�0e  51D Q  ��    � 
 �@�� ��@cp:@�AM�|(��L���L�QD�03s��3�T0 k� ��	��	%�0e  51D Q  ��    � 
 �@�� ��@ct;@�AM�|(��L���L�RD�44���3�T0 k� ��	��	%�0e  51D Q  ��    � 
 �@�� ��@ct;@�AM�|(��L�� L�RD�45���3�T0 k� ��
��
%�0e  51D Q  ��    � 
 �@�� ��@cx;@�AM�|(��	L�� L�SD�46���3�T0 k� ����%�0e  51D Q  ��    � 
 �@�� ��@c|;@�AM�|(��L��L�TD�47���3�T0 k� ����%�0e  51D Q  ��    � 
 �@�� ��@c|;@�AM�|(��L��L�UD�48���3�T0 k� ����%�0e  51D Q  ��    � 
 �@�� ��@c�<@�@M�|(��L��L�UD�8:���3�T0 k� ����%�0e  51D Q  ��    � 
 �@�� ��@c�<@�@M�|(��L��L� VD�8;���3�T0 k� ����%�0e  51D Q  ��    � 
 �@�� ��@c�<@�@M�|(��L��L� WD�8<���3�T0 k� ����%�0e  51D Q  ��    � 
 �@�� ��@c�<@�@M�|(��L��L�$XD�8=���3�T0 k� ����%�0e  51D Q  ��    � 
 �@�� ��@c�<@�@M�|(��L��L�$XD�8?���3�T0 k� ����%�0e  51D Q  ��    � 
 �@�� ��@c�=@�@M�|(��L��L�(YD�8@���3�T0 k� ��� %�0e  51D Q  ��    � 
 �@�� ��@c�=@�@M�|(� L��L�(ZD�8A���3�T0 k� ��� %�0e  51D Q  ��    � 
 �@�� ��@c�=@�@M�|(� L��L�,ZD�8B���3�T0 k� � �%�0e  51D Q  ��    � 
 �@�� ��@c�=@�@M�|(�L� L�,[I�8C���3�T0 k� � �%�0e  51D Q  ��    � 
 �@�� ��@c�=@�@M�|(�L�L�0\I�8D���3�T0 k� ��%�0e  51D Q  ��    � 
 �@�� ��@c�>@�@M�|(�L�L�0\I�8E���3�T0 k� ��%�0e  51D Q  ��    � 
 �@�� ��@c�>@�@M�|(�L�L�0]I�8F���3�T0 k� ��%�0e  51D Q  ��    � 
 �@�� ��@c�>@�@M�|(�L�L�4^I�8G���3�T0 k� ��%�0e  51D Q  ��    � 
 �@�� ��@c�>@�@M�|(� L�L�4^I�8H���3�T0 k� ��%�0e  51D Q  ��    � 
 �@�� ��@c�>@�@M�|(�!L�L�8_I�8I���3�T0 k� �!�!%�0e  51D Q  ��    � 
 �@�� ��@c�?@�@M�|(�"L� L�8_I�8J���3�T0 k� �"�"%�0e  51D Q  ��    � 
 �@�� ��@c�?@�@M�|(�#L�$Ls8`I�8J���3�T0 k� �#�#%�0e  51D Q  ��    � 
 �@�� ��@c�?@�@M�|(�%L�(Ls<aI�8K���3�T0 k� �$�$%�0e  51D Q  ��    � 
 �@�� ��@c�?@�@M�|(�&L�(	Ls<aI�8K���3�T0 k� �&�&%�0e  51D Q  ��    � 
 �@�� ��@c�?@�@M�|(�'Lq,	Ls<bI�8L���3�T0 k� �'�'%�0e  51D Q  ��    � 
 �@�� ��@c�?@�@M�|(�(Lq0	Ls@bI�8L���3�T0 k� �(�(%�0e  51D Q  ��    � 
 �@�� ��@c�@@�@M�|(�)Lq4
Ls@cI�8M���3�T0 k� �)� )%�0e  51D Q  ��    � 
 �@�� ��@c�@@�@M�|(� *Lq8
D�DcI�8M���3�T0 k� �*� *%�0e  51D Q  ��    � 
 �@�� ��@c�@@�@M�|(� +Lq<
D�DdI�8N���3�T0 k� � +�$+%�0e  51D Q  ��    � 
 �@�� ��@c�@@�@M�|(�$,Lq@D�DeI�8N���3�T0 k� � ,�$,%�0e  51D Q  ��    � 
 �@�� ��@c�@@�@M�|(�$-D�DD�HeI�8N���3�T0 k� �$-�(-%�0e  51D Q  ��    � 
 �@�� ��@c�@@�@M�|(�$.D�HD�LfI�8N���3�T0 k� �$.�(.%�0e  51D Q  ��    � 
 �@�� ��@c�@@�@M�|(�(/D�LD�LgI�8O���3�T0 k� �$/�(/%�0e  51D Q  ��    � 
 �@�� ��@c�A@�@M�|(�(0D�PD�PgI�8O���3�T0 k� �(0�,0%�0e  51D Q  ��    � 
 �@�� ��@c�A@�@M�|(�,2D�XD�TiI�8O���3�T0 k� �,2�02%�0e  51D Q  ��    � 
 �@�� ��@c�A@�@M�|(�,3D�\D�TiI�8O���3�T0 k� �,3�03%�0e  51D Q  ��    � 
 �@�� ��@c�A@�@M�|(�04D�`D�XjI�8O���3�T0 k� �,4�04%�0e  51D Q  ��    � 
 �@�� ��@c�A@�@M�|(�05D�dD�XkI�8O���3�T0 k� �05�45%�0e  51D Q  ��    � 
 �@�� ��@c�A@�@M�|(�46D�hD�XkI�8O���3�T0 k� �06�46%�0e  51D Q  ��    � 
 �@�� ��@c�B@�@M�|(�47D�pD�\lI�8O���3�T0 k� �47�87%�0e  51D Q  ��    � 
 �@�� ��@c�B@�@M�|(�48D�tD�\lI�8Os��3�T0 k� �48�88%�0e  51D Q  ��    � 
 �@�� ��@c�B@�@M�|(�89D�xD�\lI�8Os��3�T0 k� �49�89%�0e  51D Q  ��    � 
 �@�� ��@c�B@�@M�|(�8:D�|D�\mA�8Os��3�T0 k� �8:�<:%�0e  51D Q  ��    � 
 �@�� ��@c�B@�@M�|(�8:D�D�`mA�8Os��3�T0 k� �8:�<:%�0e  51D Q  ��    � 
 �@�� ��@c�B@�@M�|(�<;D�D�`mA�8Os��3�T0 k� �8;�<;%�0e  51D Q  ��    � 
 �@�� ��@c�B@�@M�|(�<<D�D�`nA�8Os��3�T0 k� �<<�@<%�0e  51D Q  ��    � 
 �@�� ��@c�B@�@M�|(�<=D�D�`nA�8Os��3�T0 k� �<=�@=%�0e  51D Q  ��    � 
 �@�� ��@c�B@�@M�|(�@>D�D�`nA�8Os��3�T0 k� �<>�@>%�0e  51D Q  ��    � 
 �@�� ��@c�C@�@M�|(�@>D�D�`nA�8Os��3�T0 k� �@>�D>%�0e  51D Q  ��    � 
 �@�� ��@c�C@�@M�|(�@?D�D�`nA�8Os��3�T0 k� �@>�D>%�0e  51D Q  ��    � 
 �@�� ��@c�C@�@M�|(�@?D�D�`nA�8Os��3�T0 k� �@?�D?%�0e  51D Q  ��    � 
 �@�� ��@c�C@�@M�|(�@?D�D�`nA�8P ��3�T0 k� �@?�D?%�0e  51D Q  ��    � 
 �@�� ��@c�C@�@M�|( �@@D�D�`nA�8P ��3�T0 k� �<D�@D%�0e  51D Q  ��    � 
 �@�� ��@c�C@�@M�|( �D@D�D�`nA�8P ��3�T0 k� �8G�<G%�0e  51D Q  ��    � 
 �@�� ��@c�C@�@M�|( �D@D��@`nA�8P ��3�T0 k� �8J�<J%�0e  51D Q  ��    � 
 �@�� ��@c�C@�@M�|( �D@D�� @`nA�8P ��3�T0 k� �8K�<K%�0e  51D Q  ��    � 
 �@�� ��@c�C@�@M�|( �H@D��!@`nA�8P c��3�T0 k� �8L�<L%�0e  51D Q  ��    � 
 �@�� ��@c�DA @M�|( �H@Lq�#@`nL38P c��3�T0 k� �<M�@M%�0e  51D Q  ��    � 
 �@�� ��@c�DA @M�|( �H@Lq�$@`nL38Q c��3�T0 k� �<N�@N%�0e  51D Q  ��    � 
 �@�� ��@c�DA @M�|( �HALq�%@c`nL38Q c��3�T0 k� �<O�@O%�0e  51D Q  ��    � 
 �@�� ��@c�DA @M�|( �LALq�&@c`nL38Q c��3�T0 k� �<O�@O%�0e  51D Q  ��    � 
 �@�� ��@c�DA @M�|( �LALq�'@c`nL38Q ���3�T0 k� �@O�DO%�0e  51D Q  ��    � 
 �@�� ��@c�DA @M�|( �LALq�(@c`nL38Q ���3�T0 k� �@O�DO%�0e  51D Q  ��    � 
 �@�� ��@c�DA @M�|( �PALq�)@c`nL38Q ���3�T0 k� �@P�DP%�0e  51D Q  ��   � 
 �@�� ��@c�DA @M�|( �PBLq�*@�`nL38Q ���3�T0 k� �DP�HP%�0e  51D Q  ��    � 
 �@�� ��@c�DA@M�|( �PBLr +@�`nL38Q ���3�T0 k� �DP�HP%�0e  51D Q  ��    � 
 �@�� ��@c�DA@M�|( �PBLr,@�`nL38Q���3�T0 k� �DP�HP%�0e  51D Q  ��    � 
 �@�� ��@c�DA@M�|( �TBLr-@�`nL38R���3�T0 k� �DP�HP%�0e  51D Q  ��    � 
 �@�� ��@c�EA@M�|( �TBLr.@�`nL38R���3�T0 k� �HQ�LQ%�0e  51D Q  ��    � 
 �@�� ��@c�EA@M�|( �TCLr/C�`nL38R���3�T0 k� �HQ�LQ%�0e  51D Q  ��    � 
 �@�� ��@c�EA@M�|( �TCL�0C�`nL38R���3�T0 k� �HQ�LQ%�0e  51D Q  ��    � 
 �@�� ��@c�EA@M�|( �XCL� 1C�`nLC8R���3�T0 k� �HQ�LQ%�0e  51D Q  ��    � 
 �@�� ��@c�EA@M�|( �XCL�$2C�\nLC8R���3�T0 k� �LQ�PQ%�0e  51D Q  ��    � 
 �@�� ��@c�EA@M�|( �XCL�(3C�\mLC8R���3�T0 k� �LR�PR%�0e  51D Q  ��    � 
 �@�� ��@c�EA@M�|( �XDL�04C�\mLC8R���3�T0 k� �LR�PR%�0e  51D Q  ��    � 
 �@�� ï@c�EA@M�|( �\DL�45C�\mLC8R���3�T0 k� �LR�PR%�0e  51D Q  ��    � 
 �@�� ï@c�EA@M�|( �\DL�85C�XmLC8R���3�T0 k� �PR�TR%�0e  51D Q  ��    � 
 �@�� ï@c�EA@M�|( �\DL�<6C�XlLC8S�� 3�T0 k� �PR�TR%�0e  51D Q  ��    � 
 �@�� ï@c�EA@M�|( �\DL�@7C�XlLC8S��3�T0 k� �PR�TR%�0e  51D Q  ��    � 
 �@�� ï@c�EA@M�|( �\DL�D8C�TkLC8S��3�T0 k� �PS�TS%�0e  51D Q  ��    � 
 �@�� ï@c�FA@M�|( �`EL�H9C�TkLC8S��3�T0 k� �TS�XS%�0e  51D Q  ��    � 
 �@�� ï@c�FA@M�|( �`EL�L9C�PkLC8S��"s�T0 k� �TS�XS%�0e  51D Q  ��    � 
 �@�� ï@c�FA@M�|( �`EL�P:C�PjLC8S3�"s�T0 k� �TS�XS%�0e  51D Q  ��   � 
 �@�� ï@c�FA@M�|( �`EL�T;C�PjLC8S3�"s�T0 k� �TS�XS%�0e  51D Q  ��   � 
 �@�� ï@c�FA@M�|( �`EL�X<C�PjLC8S3�"s�T0 k� �TS�XS%�0e  51D Q  ��    � 
 �@�� î@c�FA@M�|( �dEL�\<C�LiLC8S3�"s�T0 k� �XT�\T%�0e  51D Q  ��    � 
 �@�� Ǯ@c�FA@M�|( �dEL�`=C�LiLC8S3�"s�T0 k� �XT�\T%�0e  51D Q  ��    � 
 �@�� Ǯ@c�FA@M�|( �dFL�d>C�LiLC8S3�"s�T0 k� �XT�\T%�0e  51D Q  ��    � 
 �@�� Ǯ@c�FA@M�|( �dFL�h?C�LiLC8S3�	"s�T0 k� �XT�\T%�0e  51D Q  ��    � 
 �@�� Ǯ@c�FA@M�|( �dFL�l?C�LiLC8T3�
"s�T0 k� �XT�\T%�0e  51D Q  ��    � 
 �@�� Ǯ@c�FA@M�|( �hFL�p@C�LiLC8T3|"s�T0 k� �XT�\T%�0e  51D Q  ��    � 
 �@�� Ǯ@c�FA@M�|( �hFL�tAC�LiLC8T3x"s�T0 k� �\T�`T%�0e  51D Q  ��    � 
 �@�� Ǯ@c�FA@M�|( �hFL�xAALiLC8TCx3�T0 k� �\T�`T%�0e  51D Q  ��    � 
 �@�� Ǯ@c�FA@M�|( �hFL�xBALiLC8TCt3�T0 k� �\U�`U%�0e  51D Q  ��    � 
 �@ù Ǯ@c�FA@M�|( �hGL�|CALiLC8TCt3�T0 k� �\U�`U%�0e  51D Q  ��    � 
 �@ù Ǯ@c�FA@M�|( �hGL��CALiLC8TCp3�T0 k� �\U�`U%�0e  51D Q  ��    � 
 �@ù Ǯ@c�GA@M�|( �lGL��DALiLC8TCl4 T0 k� �`U�dU%�0e  51D Q  ��    � 
 �@ù Ǯ@c�GA@M�|( �lGL��ECCLhLC8TCl4 T0 k� �`U�dU%�0e  51D Q  ��    � 
 �@ù Ǯ@c�GA@M�|( �lGL��ECCLhLC8TCh4 T0 k� �`U�dU%�0e  51D Q  ��    � 
 �@ù ˮ@c�GA@M�|( �lGL��FCCLhLC8TCh4 T0 k� �`U�dU%�0e  51D Q  ��    � 
 �@ù ˮ@c�GA@M�|( �lGL��FCCLgLC8TCd4 T0 k� �`V�dV%�0e  51D Q  ��    � 
 �@ù ˮ@c�GA@M�|( �lGL��GCCLgLC8TCd4 T0 k� �`V�dV%�0e  51D Q  ��    � 
 �@ù ˮ@c�GA@M�|( �pHL��GK�LgLC8TC`4 T0 k� �dV�hV%�0e  51D Q  ��    � 
 �@ù ˮ@c�GA@M�|( �pHL��HK�LgLC8TC`"� T0 k� �dV�hV%�0e  51D Q  ��    � 
 �@ù ˮ@c�GA@M�|( �pHL��IK�LfLC8US\!"� T0 k� �dV�hV%�0e  51D Q  ��    � 
 �@ù ˮ@c�GA@M�|( �pHL��IK�LfLC8US\#"� T0 k� �dV�hV%�0e  51D Q  ��    � 
 �@ù ˮ@c�GA@M�|( �pHL��JK�LfLC8USX%"� T0 k� �dV�hV%�0e  51D Q  ��    � 
 �@ø ˮ@c�GA@M�|( �pHL��JK�LfLC8USX&"� T0 k� �dV�hV%�0e  51D Q  ��    � 
 �@Ǹ ˮ@c�GA@M�|( �pHL��KK�LeLC8UST("� T0 k� �dV�hV%�0e  51D Q  ��    � 
 �@Ǹ ˮ@c�GA@M�|( �tHL��KK�LeLC8UST*"� T0 k� �hW�lW%�0e  51D Q  ��    � 
 �@Ǹ ˮ@c�GA@M�|( �tHL��LK�LeLC8USP,"� T0 k� �hW�lW%�0e  51D Q  ��    � 
 �@Ǹ ˮ@c�GA@M�|( �tHLr�LK�LeLC8USP."� T0 k� �hW�lW%�0e  51D Q  ��    � 
 �@Ǹ ˮ@c�GA@M�|( �tILr�MK�LeL38USL0"� T0 k� �hW�lW%�0e  51D Q  ��    � 
 �@Ǹ ˮ@c�GA@M�|( �tILr�MK�LeL38USL3"� T0 k� �hW�lW%�0e  51D Q  ��    � 
 �@Ǹ ˭@c�GA@M�|( �tILr�NK�LeL38USL54T0 k� �hW�lW%�0e  51D Q  ��    � 
 �@Ǹ ϭ@c�HA@M�|( �tILr�NK�LeL38UcH74T0 k� �hW�lW%�0e  51D Q  ��    � 
 �@Ǹ ϭ@c�HA@M�|( �xILr�OK�LeL38UcH94T0 k� �hW�lW%�0e  51D Q  ��    � 
 �@Ǹ ϭ@c�HA@M�|( �xID��OK�LeL38UcD;4T0 k� �lW�pW%�0e  51D Q  ��    � 
 �@Ǹ ϭ@c�HA@M�|( �xID��PK�LeL38UcD=4T0 k� �lW�pW%�0e  51D Q  ��    � 
 �@Ǹ ϭ@c�HA@M�|( �xID��PK�LeL38UcD?4T0 k� �lW�pW%�0e  51D Q  ��    � 
 �@Ǹ ϭ@c�HA@M�|( �xID��QK�LeA�8U	S@A4T0 k� �lX�pX%�0e  51D Q  ��    � 
 �D���m��B�\d%<��%��k�|{�E��KD��E��̿�3� T0 k� ������%�0e  51D Q  ��Z    ����8D���m��B�`d%<��%��k�|{�E��JD��E��̿�3� T0 k� ������%�0e  51D Q  ��Z    ����8D���m��B�`d%<��
��k�|w�E��HD��E��̻�3� T0 k� ������%�0e  51D Q  ��Z    ����8D��m��B�`d%<��
��k�|w�E��GD��E��̻�3� T0 k� ������%�0e  51D Q  ��Z    ����8D��m��B�dd%<��
��k�|w�E��ED��E��̻�3� T0 k� ������%�0e  51D Q  ��Z    ����8D��m��B�hd%<��
���k�|w�E��BD��E��̷�3� T0 k� ������%�0e  51D Q  $�Z    ����8D��m��B�hd%<��
���k�|s�C��AE�E�{�̳�3� T0 k� <�����%�0e  51D Q  ��_    ����8D��m��B�hd%<��
���k�|s�C��?E�E�s�̳�3� T0 k� <�����%�0e  51D Q  ��_    ����8D��m��B�hd%<��
���o�|s�C��>E�E�k�ܯ�3� T0 k� <�����%�0e  51D Q  ��_    ����8D��}��B�ld%<��
���o�|s�C��<E�E�c�ܯ�3� T0 k� <�����%�0e  51D Q  ��_    ����8D��}��B�ld%<��
���k�|o�C��:E�E�[�ܯ�3� T0 k� <�����%�0e  51D Q  ��_    ����8D��}��B�ld%<������g�|o�E��7BM�E�[�ܯ�3� T0 k� ������%�0e  51D Q  ��_    ����8D��}��B�ld%<�����|g�|o�E��5BM�E�W�ܫ�3� T0 k� ������%�0e  51D Q  ��_    ����8D��}��B�ld%<�����|` |k�E��4BM�E�W�ܫ�3� T0 k� ������%�0e  51D Q  ��_    ����8D��}��B�ld%<�����|`|k�E��2BM�E�S�ܫ�3� T0 k� ������%�0e  51D Q  ��_    ����8D��}��@ld%<�����|\|k�E��0BM�E�O�ܤ 3� T0 k� ������%�0e  51D Q  ��_    ����8D��}��@ld%<�����|\|k�E��.A��FK�ܤ3� T0 k� ������%�0e  51D Q  ��_    ����8D��}��@ld������|X|k�E��-A��FG�ܠ3� T0 k� ������%�0e  51D Q  ��_    ����8D��}��@ld������|T|g�E��)A��FC�ܠ3� T0 k� �� �� %�0e  51D Q  ��_    ����8D��M��@mld������|P|g�E��'A��FC�ܘ3� T0 k� �� �� %�0e  51D Q  ��_    ����8D��M��@mld������|L	|g�E��&A��F?�ܔ3� T0 k� �� �� %�0e  51D Q  ��_    ����8D��M��@mld������|H
|g�E��$A��F?�ܐ3� T0 k� �� �� %�0e  51D Q  ��_    ����8D��M��@mld�����|D|c�E��"A��F;�܌	3� T0 k� �� �� %�0e  51D Q  ��_    ����8D��M��@mld�����|@|c�E�� A��D�;�\�
3� T0 k� �� �� %�0e  51D Q  ��_    ����8D��	]��@mld�����|<|c�E��A��D�7�\�3� T0 k� ����%�0e  51D Q  ��_    ����8D��	]��@mld�����|8|c�E��A��D�7�\�3� T0 k� ����%�0e  51D Q  ��_    ����8I��	]��@mld�����|0|_�E��A]�D�7�\x3� T0 k� ����%�0e  51D Q  ��_    ����8I��	]��@mld�����|,|_�E��A]�D�7�\t3� T0 k� ����%�0e  51D Q  ��_    ����8I��	m��@mld�#����|(|_�E��A]�F3�\p3� T0 k� ����%�0e  51D Q  ��_    ����8I��	m��@mld�'����|$|_�E��A]�F3�\l3� T0 k� ����%�0e  51D Q  ��_    ����8I��	m��@mld�+����| |_�E��A]�F3�\h3� T0 k� ��� %�0e  51D Q  ��_    ����8I��	m��@mld�/����| |_�E��C��F3�\d3� T0 k� � �%�0e  51D Q  ��_    ����8I��	m��@mldM3����| |[�E��C��F3�\`3� T0 k� � �%�0e  51D Q  ��_    ����8I��	]�@mldM;����| |[�E��C��F3�\`3� T0 k� ��%�0e  51D Q  ��_    ����8I��	]�@mldM?����||[�E��C��F7�\`3� T0 k� ��%�0e  51D Q  ��_    ����8I��	]�@�ldMC����||[�E��C��E�7�\`3� T0 k� ��%�0e  51D Q  ��_    ����8I��	]�@�ldMG����||[�D<�C��E�7�\\3� T0 k� ��%�0e  51D Q  ��_    ����8I��	]�@�ldMK����||W�D<�C��E�7�\\3� T0 k� ��%�0e  51D Q  ��_    ����8I� 	m�@�ldMO����||W�D<�
C��E�;�\\3� T0 k� ��%�0e  51D Q  ��_    ����8I�	m�
CMld]W����||W�D<�C��E�?�\\3� T0 k� � �$%�0e  51D Q  ��_    ����8I�	m�CMlc][����||W�E�C��E�?�\\3� T0 k� �$�(%�0e  51D Q  ��_    ����8I�	m�CMlc][����|�W�E�C��E�C�\\3� T0 k� �$�(%�0e  51D Q  ��_    ����8I�	]�CMlc]_����|�W�E�C��E�C��\3� T0 k� �(�,%�0e  51D Q  ��_    ����8I�	]�CMlb�g����|�S�E�C��E�K��\3� T0 k� �0�4%�0e  51D Q  ��_    ����8I�	]�CMla�k����|�S�E�C��E�K��\3� T0 k� �4�8%�0e  51D Q  ��_    ����8I�	]�CMl`�o����|�S�E�C��E�O��\3� T0 k� �4�8%�0e  51D Q  ��_    ����8I�	m�C]l`�s����|�S�E�C��E�S��\3� T0 k� �8�<%�0e  51D Q  ��_    ����8I�
	m�C]l^�w���|�S�E�D�E�W��\3� T0 k� �@�D%�0e  51D Q  ��_    ����9I�
	m�C]l^�{���|lO�E�xD�E�[��\3� T0 k� �L�P%�0e  51D Q  ��3    ����:I�	m�C]l]=���|lO�E�tD�E�_��\3� T0 k� �X�\%�0e  51D Q  ��3    ����;I�	]�C]l[=����| lO�E�lD�E�g��`3� T0 k� �h�l%�0e  51D Q  ��3    ����<I�	]�C]lZ=����| lO�E�hE]�E�k��`3� T0 k� �p�t%�0e  51D Q  ��3    ����=I�	]�C]lX=���'�| lK�E�`E]�E�s��`3� T0 k� �x	�|	%�0e  51D Q  �3    ����=I�	]�C]lW=���+�| lG�E�\E]�E�w��`3� T0 k� �x	�|	%�0e  51D Q  ��3    ����=I�	m�CmlV=���3�| lG�E�XE]|E�w��`3� T0 k� �x�|%�0e  51D Q  ��3    ����=BN	m�CmlT=���;�|$�C�E�PE]pE.��d3� T0 k� �x	�|	%�0e  51D Q  ��3    ����>BN	m�CmlS-���C�!�$�?�E�PE]lE.��d3� T0 k� ����%�0e  51D Q  �3    ����?BNM�E-lP-���O�!� �;�R�PE�`E.��h3� T0 k� ����%�0e  51D Q  ��3    ����@BNM�E-lO-���S�!� �;�R�PE�X	E.��h3� T0 k� ����%�0e  51D Q  ��3    ����AFM�E-pM���_�!� �3�R�TE�L
E.��l3� T0 k� ����%�0e  51D Q  ��3    ����BFM�E-pK���g�!� �3�R�TE�DE.���p3� T0 k� ��	��	%�0e  51D Q  ��3    ����CFM�E-tJ���o�!� �/�R�TE�<E.���t3� T0 k� ��
��
%�0e  51D Q  ��3    ����DFM�E-tI���s�!� �/�R�TE�8E���t3� T0 k� ����%�0e  51D Q  ��3    ����EE� M� E-xF-����!� �+�R�X I�(E���|3� T0 k� ����%�0e  51D Q  ��3    ����FE� ]�!E-xE-�����| '�R�X I� E����3� T0 k� ����%�0e  51D Q  ��3    ����GE�$]�"E|C-� ���| '�R�[�I�E����3� T0 k� ����%�0e  51D Q  ��3    ����IE�(]�$E�A-����|$#�R�[�I�B�����3� T0 k� ����%�0e  51D Q  ��3    ����KB�,]�%E�?-����|$
#�R�_�I�B�����3� T0 k� ����%�0e  51D Q  ��3    ����MB�0]�'E�>-����|$
#�R�_�I�B�����3� T0 k� ����%�0e  51D Q  ��3    ����OB�4]�(E�=-����|$
#�R�_�I��B�����3� T0 k� ����%�0e  51D Q  ��3    ����QB�8]�+E�=-�	���|$	#�R�_�I��B�����3� T0 k� ����%�0e  51D Q  ��3    ����TB�<]�+E�=-�
���|$	�#�R�c�I��B�����3� T0 k� ����%�0e  51D Q  ��3    ����WB�@]�+E�>-����|$	�#�R�c�E\�B�����3� T0 k� ����%�0e  51D Q  ��3    ����ZB�Dm�+E�>-����!�$	�#�R�c�E\�B�����3� T0 k� ����%�0e  51D Q  ��3    ����]B�Hm�,E��>����!�$�#�R�c�E\�B�����3� T0 k� ����%�0e  51D Q  ��3    ����`B�Tm�-E��?����!�$�#�R�c�E\�B����3� T0 k� ����%�0e  51D Q  ��3    ����cB�Xm�-E��?�L��!�$'�R�g�A\�B����3� T0 k� ����%�0e  51D Q  ��3    ����fB�\m�.E��@�L��!�$'�R�g�A\�B����3� T0 k� ����%�0e  51D Q  ��3    ����iB�`m�.E��@�L��!�$'�R�g�A\�B�#���3� T0 k� ����%�0e  51D Q  ��3    ����lB�hm�/E��@�L��!�$+�R�g�A\�B�+���3� T0 k� ����%�0e  51D Q  ��3    ����oB�lm�0E��A�M�!�$+�R�g�A\�B�3���3� T0 k� ����%�0e  51D Q  ��3    ����sB�xm�1E��B�M�!�$/�R�k�A�B�C���3� T0 k� ����%�0e  51D Q  ��3    ����wB�|}�2E}�C�M�|$3�R�k�A�B�K�̨3� T0 k� ����%�0e  51D Q  ��3    ����{B΀}�3E}�C�M�|$3�R�k�A�B�S�̨3� T0 k� ����%�0e  51D Q  ��3    ����BΈ }�4E}�D�M#�|$7�R�k�A�B�[�̨3� T0 k� ����%�0e  51D Q  ��3    �����Bΐ }�5E}�E�M'�|$7�R�k�A�B�c�̬3� T0 k� � �%�0e  51D Q  �3    �����BΜ!��7E}�FM�!M3�|$�?�R�o�@��Es�̬3� T0 k� � �$%�0e  51D Q  ��?    �����BΠ!��8E}�GM�"]7�|$�C�R�o�@��E{�̬
3� T0 k� �0�4%�0e  51D Q  ��?    �����BΨ"��:D��HM�#]?�|$�C�R�o�@��E��̬
3� T0 k� �@�D%�0e  51D Q  ��?    �����Bά"��;D��IM�$]C�|$�G�R�o�@��E��̰	3� T0 k� �P�T%�0e  51D Q  ��?    �����Bδ"��<D��JN %]G�|$�K�R�o�@��E��̴	3� T0 k� �`�d%�0e  51D Q  ��?    �����Bθ#͘=D��KN&]O�|$�O�R�o�@l�E��̴3� T0 k� �p�t%�0e  51D Q  ��?    �����B��#͘?D��L^'�S�|$�S�R�s�@l�E��ܸ3� T0 k� ����%�0e  51D Q  ��?    �����B��$͘@D��M^(�W�|$�W�R�s�@l�E��ܼ3� T0 k� ����%�0e  51D Q  ��?    �����B��$͘AF�O^)�[�|$�_�R�s�@l�E��ܼ3� T0 k� ����%�0e  51D Q  ��?    �����B��$͘BF�P^*�_�|$�c�R�s�@m E����3� T0 k� �� �� %�0e  51D Q  ��?    �����B��%	}�CF�Q^+�g�|$�g�R�s�B�E�����3� T0 k� ��!��!%�0e  51D Q  ��?    �����B��%	}�EF�Rn ,�k�|$�k�R�s�B�E�����3� T0 k� ��"��"%�0e  51D Q  ��?    �����B��&	}�FF�Sn$-�o�|$�s�R�s�B�
E�����3� T0 k� ��"��"%�0e  51D Q  ��?    �����B��&	}�GF�Tn(.�s�|$�w�R�s�B�	E�����3� T0 k� ��#��#%�0e  51D Q  ��?    �����B��&	}�GF�Vn,/�w�|$�{�R�w�B�E�����3� T0 k� �$�$%�0e  51D Q  ��     �����E��'	��HF Wn00�{�|$���R�w�B� E�����3� T0 k� �$�$%�0e  51D Q  ��     �����E��'	��IFXn40��|$���R�w�B�(E�����3� T0 k� �%�%%�0e  51D Q  ��     �����E�'	��JFZn81��|$���R�w�B�,E�����3� T0 k� �%�%%�0e  51D Q  ��     �����E�(	��KF[n<2̓�|$���R�w�B�0E����3� T0 k� � %�$%%�0e  51D Q  ��     �  ��E�(	��KE�\n@3͇�|$���R�w�B�4E����3� T0 k� �(&�,&%�0e  51D Q  ��     �  ��E�)	}�LE�]nD4͋�|$���R�w�B�8D����3� T0 k� �,&�0&%�0e  51D Q  ��     � ��E�)	}�LE�_nH5͋�|$���R�w�B�@ D����3� T0 k� �4&�8&%�0e  51D Q  ��     � ��E�$)	}�ME� `nL5͏�|$���R�{�B�G�D�'�� 3� T0 k� �<'�@'%�0e  51D Q  ��     �  E�,*	}�ME�$anP6͏�|$���R�{�B�K�D�/��3� T0 k� �D$�H$%�0e  51D Q  ��     �  E�4*	}�NE�,bnT7͐ |$���R�{�B�O�D�7��3� T0 k� �L!�P!%�0e  51D Q  ��     �  E�8*	��NE�0dnX8ݐ|$�ëR�{�B�S�D�?��3� T0 k� �T �X %�0e  51D Q  ��     �  E�@*	��OE�4en\8ݔ|$�˪R�{�B�W�D�G��3� T0 k� �\�`%�0e  51D Q  ��     �  	E�H*	��OE�<fn\9ݔ|$�өR�{�B�_�D�O��3� T0 k� �d�h%�0e  51D Q  ��     �  EP+	��OB�@gn`:ݔ|$�רR�{�B�c�D�W�� 3� T0 k� �h"�l"%�0e  51D Q  ��     �  EX+	��OB�Hhnd;ݔ	|$�ߧR�{�B�g�D�_��$ 3� T0 k� �l%�p%%�0e  51D Q  ��     �  E\+	}�PB�Linh;ݔ
|$��R�{�B�k�D�g��( 3� T0 k� �p(�t(%�0e  51D Q  ��     �  Ed+	}�PB�Tjnl<ݔ|$��R�{�B�o�D�o��0 3� T0 k� �x*�|*%�0e  51D Q  ��     �  El+	}�PB�Xknl=ݔ|$���R��B�w�D�w��?�3� T0 k� ��+��+%�0e  51D Q  ��     �  Et,	}�PB�`lnp=ݔ|$���R��E-{�D���K�3� T0 k� ��,��,%�0e  51D Q  ��     �  E|,	}�PB�dmnt>ݔ|$��R��E-�D����K�3� T0 k� ��-��-%�0e  51D Q  ��     �  E�,	��PB�lnnt>�|$��R��E-��D����S�3� T0 k� ��/��/%�0e  51D Q  ��     �  @/�,	��PB�ponx?�|$��R��E-��D����_�3� T0 k� ��.��.%�0e  51D Q  ��     �  @/�,	��PB�xpnx?�|$��R��E-��D����k�3� T0 k� ��-��-%�0e  51D Q  ��     �  @/�-	��PB��qn|@�|$�#�R��E��D���s�3� T0 k� ��-��-%�0e  51D Q  ��     �  !@/�-	��PB��rn|@�|$�+�R��E��D����3� T0 k� ��-��-%�0e  51D Q  ��     �  #@/�-]�PB��sn�@݌|$�3�R��E��D�����3� T0 k� ��-��-%�0e  51D Q  ��     �  %@/�-]�PB��tn�@݌|$�7�R��E��F �����3� T0 k� � .�.%�0e  51D Q  ��     �  '@/�-]�PB��un�A݈|$�?�R��E��F �����3� T0 k� �.�.%�0e  51D Q  ��     �  )@/�-]�PB��vn�A݈|$�G�R���B���F �����3� T0 k� �.�.%�0e  51D Q  ��     �  +@/�.]�PB��wn�A݄ |$�O�R���B���F �����3�T0 k� �.� .%�0e  51D Q  ��     �  -@/�.��PB��xn�A݄!|$�W�R���B���F �����3�T0 k� �$.�(.%�0e  51D Q  ��     �  /@/�.��PB��xn�A݀#|$�_�R���B���F �����3�T0 k� �,.�0.%�0e  51D Q  ��     �  1@/�.��PB��yn�B݀$|$�g�R���B���F �����3�T0 k� �4/�8/%�0e  51D Q  ��     �  3@?�.��PB��zn�B�|%|$�o�R���B���F �����3�T0 k� �@/�D/%�0e  51D Q  ��     �  5@?�.��PB��{n�B�|'|$�w�R���B���F �����3�T0 k� �L/�P/%�0e  51D Q  ��     �  7@?�.��PB��|n�B�x(|$��R���B���F����3�T0 k� �X/�\/%�0e  51D Q  ��     �  9@?�/��PB��}n�B�x)|$݇�R���B���BA����3�T0 k� �`/�d/%�0e  51D Q  ��     �  ;@0/��PB��}n�B�t*|$݋�R���B���BA����3�T0 k� �h/�l/%�0e  51D Q  ��     �  =E/��PB��~n�C�t,|$���R���B���BA���3�T0 k� �\1�`1%�0e  51D Q  ��     �  ?E/��PB��n�C�t-|$���R���B���BA���3�T0 k� �T2�X2%�0e  51D Q  ��     �  AE/ݘPB� �n�C�p.|$���R���B��BA'���3�T0 k� �L2�P2%�0e  51D Q  ��     �  CE$/ݘOB�n�C�p/|$���R���B��BA+���3�T0 k� �L2�P2%�0e  51D Q  ��     �  EE,/ݘOB�n�C�l0|$���R���B��BA3��#�3�T0 k� �L2�P2%�0e  51D Q  ��     �  GE40ݜOB�n�C�l1|$���R���B��BA7��+�3�T0 k� �P3�T3%�0e  51D Q  ��     �  IE<0ݜOB� n�D�l2|$�ÑR���B�'�BA?��3�3�T0 k� �T3�X3%�0e  51D Q  ��     �  KE@0ݜNB�(~n�D�h3|(�ːR���B�/�BAG��;�3�T0 k� �X3�\3%�0e  51D Q  ��     �  MEH0ݜNB�0~n�D�h5|(�ӐR���B�7�BAK��C�3�T0 k� �\4�`4%�0e  51D Q  ��     �  O@ P0ݠNB�<~n�D�d6|(�ۏR���B�?�BAP �K�3�T0 k� �t3�x3%�0e  51D Q  ��     �  Q@ X0ݠMB�D~n�D�d7|(��R���B�G�BAT �S�3�T0 k� ��2��2%�0e  51D Q  ��     �  S@ `0ݤMB�L}n�D�d8|(��R���B�O�BAX�[�3�T0 k� ��1��1%�0e  51D Q  ��     �  U@ h0�LB�T}n�D�`9|(��R���B�W�BA`�c�3�T0 k� ��1��1%�0e  51D Q  ��     �  W@ p1�LB�\}n�E�`:|(���R���E_�BAd�o�3�T0 k� ��1��1%�0e  51D Q  ��     � 	 Y@ x1�KB�d}n�E�`;|(��R���Eg�BAl�w�3�T0 k� ��1��1%�0e  51D Q  ��     � 	 [@ �1�KB�l}n�E�\<|(��R���Eo�BAp��3�T0 k� ��1��1%�0e  51D Q  ��     � 	 ]@ �1�JB�t|n�E�\<|(��R���Es�BAt���3�T0 k� ��2��2%�0e  51D Q  ��     � 	 _@ �1�IB߀|n�E�\=|(��R���E{�BA|���3�T0 k� ��2��2%�0e  51D Q  ��     � 	 a@ �1�IB߈|n�E�X>|(�#�R���E��BA����3�T0 k� ��2��2%�0e  51D Q  ��     � 	 c@ �1�HBߐ|n�E�X?|(�+�R���E��BA����3�T0 k� ��2��2%�0e  51D Q  ��     � 	 e@ �1�GB��|n�E�X@|(�3�R���E��BA����3�T0 k� ��2��2%�0e  51D Q  ��     � 	 g@0�1�GB��{n�F�TA|(�;�R���E��BA����3�T0 k� �2�2%�0e  51D Q  ��     � 	 i@0�2��FB��{n�F�TB|(�C�R���E��BA����3�T0 k� �2�2%�0e  51D Q  ��     � 
 k@0�2��EB��{n�F�TC|(�K�R���E���BA����3�T0 k� �2� 2%�0e  51D Q  ��     � 
 m@0�2��DB��{n�F�PC|(�S�R���E���BA����3�T0 k� �(2�,2%�0e  51D Q  ��     � 
 o@0�2��CB��{n�F�PD|(�[�R���E���BA����3�T0 k� �03�43%�0e  51D Q  ��     � 
 qE��2��BB��zn�F�PE|(�c�R���E���BA����3�T0 k� �(/�,/%�0e  51D Q  ��     � 
 sE��2��AE��zn�F�LF|(�k�R���E���BA����3�T0 k� � ,�$,%�0e  51D Q  ��     � 
 uE��2��AE��zn�F�LG|(�s�R̋�E���BA�	���3�T0 k� �)� )%�0e  51D Q  ��     � 
 wE��2��@E��zn�F�LG|(�{�R̋�E���BA�	���3�T0 k� �'� '%�0e  51D Q  ��     � 
 yE��2��?E��zn�G�LH|(΃�R̋�E���BA�	��3�T0 k� � &�$&%�0e  51D Q  ��     � 
 {E��2��>E��zn�G�HI|(΋�R̋�E���BA�
��3�T0 k� � %�$%%�0e  51D Q  ��     � 
 }@q 2��<E� yn�G�HJ|(Γ�R̋�E���BA�
��3�T0 k� �(!�,!%�0e  51D Q  ��     � 
 @q2��;E�yn�G�HJ|(Λ�R̋�D���BA��#�3�T0 k� �0�4%�0e  51D Q  ��     � 
 �@q2�:E�yn�G�HK|(ޣ�R̋�D��BA��/�3�T0 k� �8�<%�0e  51D Q  ��     � 
 �@q1�9E�yn�G�DL|(ޫ�R̋�D��BA��7�3�T0 k� �@�D%�0e  51D Q  ��     � 
 �@q 1�8E� yn�G�DL|(޳�R̋�D��BA��?�3�T0 k� �H�L%�0e  51D Q  ��  
   � 
 �E�(1�7E�(yn�G�DM|(޻�U|��D�#�BA��G�3�T0 k� �L�P%�0e  51D Q  ��  
   � 
 �E�,1 6E�4xn�G�DN|(�ÂU|��D�+�BA��S�3�T0 k� �P�T%�0e  51D Q  ��  
   � 
 �E�404E�<xn�G�@N|(�˂U|��D�3�BA��[�3�T0 k� �X�\%�0e  51D Q  ��  
   � 
 �E�<03E�Dxn�H�@O|(�ӁU|��D�;�BA��c�3�T0 k� �`�d%�0e  51D Q  ��  
   � 
 �E�D02E�Lxn�H�@P|(�ہU|��D�C�BA��o�3�T0 k� �h�l%�0e  51D Q  ��  
   � 
 �E�L/1E�Twn�H�@P|(��U|��D�K�BA��w�3�T0 k� �p�t%�0e  51D Q  ��  
   � 
 �E�T//E�\wn�H�<Q|(��U|��D�S�BA���3�T0 k� �x�|%�0e  51D Q  ��  
   � 
 �E�\/.E�dwn�H�<R|(��U|��D�[�BA�ߋ�3�T0 k� �p�t%�0e  51D Q  ��  
   � 
 �E�d.�$-E�pv��H�<R|(���U|��D�c�BA�ߓ�3�T0 k� �p�t%�0e  51D Q  ��  
   � 
 �E�h.�(+E�xv��H�<S|(��A���D�o�BA�ߛ�3�T0 k� �p�t%�0e  51D Q  ��  
   � 
 �E�p-�,*B��u��H�8S|(��A���D�w�BA�ߣ�3�T0 k� �p�t%�0e  51D Q  ��  
   � 
 �E�x-�4)B��u��H�8T|(��A���D��BA�߯�3�T0 k� �t�x%�0e  51D Q  ��  
   � 
 �E1�,�8'B�t��H�4T|(��A���D��BA�߷�3�T0 k� �x�|%�0e  51D Q  ��  	   � 
 �E1�+�@&B�t��H�4U|(�#�A���E���BB ���3�T0 k� ����%�0e  51D Q  ��  	   � 
 �E1�+�D$B�s��H�0U|(�+�BL��E���BB���3�T0 k� ����%�0e  51D Q  ��  	   � 
 �E1�*�L#E�s��I�0V|(�3�BL��E���BB���3�T0 k� ����%�0e  51D Q  ��  	   � 
 �E1�)�P!E�r��I�,V|(�;�BL��E���BB���3�T0 k� ����%�0e  51D Q  ��  	   � 
 �E!�(�X E�r��I�,V|(�C�BL��E���BB���3�T0 k� ����%�0e  51D Q  ��  	   � 
 �E!�(�\E�q��I�(V|(�K�BL��E���BB���3�T0 k� ����%�0e  51D Q  ��  	   � 
 �E!�'�`E�q��I�(V|(�S�B���E���BB���3�T0 k� ����%�0e  51D Q  ��  	   � 
 �E!�&�hE�p��I�$V|(�[�B���E���BB���3�T0 k� ����%�0e  51D Q  ��  	   � 
 �E!�%�lE�p��I�$V|(�c�B���E���BB��3�T0 k� ����%�0e  51D Q  ��  	   � 
 �@q�$�tE�o��I� V|(�k�B���B���BB��3�T0 k� ����%�0e  51D Q  ��  	   � 
 �@q�#�xE�o��I V|(�s�B���B���BB��3�T0 k� ����%�0e  51D Q  ��  	   � 
 �@q�"�B��o��IV|(�{�B���B���BB �#�3�T0 k� ����%�0e  51D Q  ��  	   � 
 �@q�"�B��n��IV|(���B���B���BB$�/�3�T0 k� ����%�0e  51D Q  ��  	   � 
 �@q�!�B�n��IV|(���B���B���BB$�7�3�T0 k� ��
��
%�0e  51D Q  ��  	   � 
 �@q� �B�m��IV|(���B���E��BB(�?�3�T0 k� � 	�	%�0e  51D Q  ��  	   � 
 �@q��B�m��I�U|(���B���E��BB,�K�3�T0 k� ��%�0e  51D Q  ��  	   � 
 �@q��E� l��J�U|(���B���E��BB,�S�"��T0 k� ��%�0e  51D Q  ��  	   � 
 �@q��E�(l��J�U|(���B���E��BB0�[�"��T0 k� ��%�0e  51D Q  �  	   � 
 �@q��E�0k��J�T|(Ϸ�B���E�'�BB8�c�"��T0 k� ��%�0e  51D Q  ��  	   � 
 �@q��
E�8k��J�T|(Ͽ�B���E�/�BB<�o�"��T0 k� �� %�0e  51D Q  ��  	   � 
 �@q��E�@j��J�S|(�ǆB���E�7�BB@�w�"��T0 k� � �$%�0e  51D Q  ��  	   � 
 �@� �E�Hj� J�S|(�φB���D�?�BBD��"��T0 k� � �$%�0e  51D Q  ��  	   � 
 �@��E�Pi�J�R|(�׆B���D�G�BBH���"��T0 k� �$�(%�0e  51D Q  ��  	   � 
 �@���B�Xh�J�R|(�߇B���D�O�BBL���"��T0 k� �(�,%�0e  51D Q  ��  	   � 
 �@���B�`h�J�Q|(��B���D�W�BBP���"��T0 k� �,�0%�0e  51D Q  ��     � 
 �@���B�hg�J�Q|(��B���D�_�BBT���"��T0 k� �0�4%�0e  51D Q  ��     � 
 �@��� B�pf�J�P|(���B���D�g�BBX���"��T0 k� �4�8%�0e  51D Q  ��     � 
 �@����B�xf�$J�O|(���B���D�o�BB\���3�T0 k� �4�8%�0e  51D Q  ��     � 
 �@����B�e�(J�O|(��B���D�w�BBd���3�T0 k� �8�<%�0e  51D Q  ��     � 
 �@����B�d�0J�N|(��B���D��I�h���3�T0 k� �<�@%�0e  51D Q  ��     � 
 �@� ���B�c�8J�M|(��B���DЇ�I�l���3�T0 k� �@�D%�0e  51D Q  ��     � 
 �@�$���B�c�<J� L|(��B���DЏ�I�p���3�T0 k� �D�H%�0e  51D Q  ��     � 
 �@�(��B�b�DJ� L|(�'�B���DЗ�I�t���3�T0 k� �H �L %�0e  51D Q  ��     � 
 �@�,��B�a�LJ� K|(�/�B���D���I�t���3�T0 k� �O��S�%�0e  51D Q  ��     � 
 �@�0��B�`�TJ�$J|(�7�B���D��I�x���3�T0 k� �W��[�%�0e  51D Q  ��     � 
 �@�4��C�`�XJ�$I|(�?�B���D��J|���3�T0 k� �[��_�%�0e  51D Q  ��     � 
 �@�8��C�_�`J�(H|(�G�B��D��J���3�T0 k� �_��c�%�0e  51D Q  �     � 
 �@�@�'�C�^�hJM(G|(�O�B��D��J���3�T0 k� �c��g�%�0e  51D Q  �     � 
 �@�@ +�C�]�lIM,F|(�W�B��E���J���"s�T0 k� �g��k�%�0e  51D Q  ��     � 
 �@�D 3�C�\�tIM,F|(�_�B��E���J��#�"s�T0 k� �k��o�%�0e  51D Q  ��     � 
 �@�H 7�@a�\�|IM0E|(�g�B��E���I��/�"s�T0 k� �o��s�%�0e  51D Q  ��     � 
 �@�L ?�@a�[O�IM0D|(�o�B�'�E���I��7�"s�T0 k� �s��w�%�0e  51D Q  ��     � 
 �@�L G�@a�ZO�IM4C|(�w�B�+�E���I��?�"s�T0 k� �w��{�%�0e  51D Q  ��     � 
 �@�P K�@a�YO�IM4B|(��B�3�E���I��G�"s�T0 k� �s��w�%�0e  51D Q  ��     � 
 �@�T S�@a�YO�HM8A|(���B�;�E���I��S�"s�T0 k� �s��w�%�0e  51D Q  ��     � 
 �@�X W�@bXO�HM8A|(���B�C�E���J��[�"s�T0 k� �s��w�%�0e  51D Q  ��     � 
 �@�\
 _�@bWO�HM<@|(���B�K�E��J��c�"s�T0 k� �s��w�%�0e  51D Q  ��     � 
 �@�`	 c�@bVO�HM<?|(���B�S�D��J��o�"s�T0 k� �s��w�%�0e  51D Q  ��     � 
 �E"d k�@bVO�HM@>|(���B�[�D��J��w�"s�T0 k� �w��{�%�0e  51D Q  ��     � 
 �E"h o�@b UO�HM@>|(���B�c�D��J���3�T0 k� �{���%�0e  51D Q  ��     � 
 �E"l s�@b$TO�HMD=|(���B�k�D�#�I����3�T0 k� ������%�0e  51D Q  ��     � 
 �E"p {�@b,TO�GMD<|(�ËB�s�D�+�I���3�T0 k� ������%�0e  51D Q  ��     � 
 �E"t �@b0SO�GMD<|(�ˋB�{�D�3�I���3�T0 k� ������%�0e  51D Q  ��     � 
 �E"x ��@b8SO�GMH;|(�ӋB���D�;�I���3�T0 k� ������%�0e  51D Q  ��     � 
 �E"� ��@b@RO�GMH:|(�یB���D�C�I���3�T0 k� ������%�0e  51D Q  ��     � 
 �E"�  ��@bDQO�GML9|(��B���D�K�BB���3�T0 k� ������%�0e  51D Q  ��     � 
 �E"�� ��@bHQO�GML9|(��B���D�S�BB���3�T0 k� ������%�0e  51D Q  ��     � 
 �E�� ��@bPPO�GML8|(��B���D�[�BB����3�T0 k� ������%�0e  51D Q  ��     � 
 �E�� ��@bTPO�FMP8|(���B���D�c�BB����3�T0 k� ������%�0e  51D Q  ��     � 
 �E�� ��@b\OO�FMP7|(�B���D�g�BB����3�T0 k� ������%�0e  51D Q  ��     � 
 �E�� ��@b`NO�FMT6|(�B���D�o�Er����3�T0 k� ������%�0e  51D Q  ��     � 
 �E�� ��@bdNO�FMT6|(�B���D�w�Er����3�T0 k� ������%�0e  51D Q  ��     � 
 �FB�� ��@blMO�FMT5|(�B���D��Er����3�T0 k� ������%�0e  51D Q  ��     � 
 �FB�� ��@bpMO�FMX4|(#�B���D��Er�	1��3�T0 k� ������%�0e  51D Q  ��     � 
 �FB�� ��@btLO�FMX4|(+�B���D��Er�	2 3�T0 k� ������%�0e  51D Q  ��     � 
 �FB�� ��@b|L@ FMX3|(3�B���D��LR�	2 3�T0 k� ������%�0e  51D Q  ��     � 
 �FB�� ��@b�K@EM\3|(;�B���D��LR�	23�T0 k� ������%�0e  51D Q  ��     � 
 �FB�� ��@b�K@EM\2|(C�B��D��LR�	23�T0 k� ������%�0e  51D Q  ��     � 
 �FB�� ��@b�J@EM\2|(K�B��D��LR�	2 3�T0 k� ������%�0e  51D Q  �     � 
 �FR�� ��@b�J@EM`1|(O�B��D��LR�	B(3�T0 k� ������%�0e  51D Q ��    � 
 �FR�� ��@b�I@EM`1|(W�B�'�D��LR�	B03�T0 k� ����%�0e  51D Q ��    � 
 �FR�� ��@b�I@EM`0|(_�B�/�D���LR�	B43�T0 k� ����%�0e  51D Q ��    � 
 �FR�� ��@b�H@ EMd0|(g�B�7�D���LR�	B<3�T0 k� ����%�0e  51D Q ��   � 
 �FR�� ��@b�H@$EMd/!�(o�B�C�D���LR�	B@3�T0 k� �'��+�%�0e  51D Q ��    � 
 �Fb�� ��@b�G@(EMd/!�(w�B�K�D���LR�	2H3�T0 k� �3��7�%�0e  51D Q ��    � 
 �Fb�� ��@b�G@,EMh.!�(��B�W�D�� Lb�	2L3�T0 k� �?��C�%�0e  51D Q ��    � 
 �Fb�� ��@b�G@0DMh.!�(���B�_�D��Lb�	2P3�T0 k� �K��O�%�0e  51D Q ��    � 
 �Fb�� ��@b�F@4DMh-!�(���B�k�D��Lb�	2X3�T0 k� �T �X %�0e  51D Q ��    � 
 �Fb�� ��@b�F@4DMh-!�(���B�s�D��Lb�	2\3�T0 k� �`�d%�0e  51D Q ��    � 
 �Fb�� ��@b�E@8DMl,!�(���B�{�D��Lb�2`3�T0 k� �l�p%�0e  51D Q ��    � 
 �Fb�� ��@b�E@<DMl,!�(���B·�D� Lb�2d3�T0 k� �x�|%�0e  51D Q ��    � 
 �Fb�� ��@b�D@@DMl+!�(���BΏ�ELb�2l3�T0 k� ����%�0e  51D Q ��    � 
 �Fb�� ��@b�D@DDMl+!�(���BΛ�ELb�2p3�T0 k� ����%�0e  51D Q ��    � 
 �Fb�� �@b�D@HDMp*!�(���BΣ�E	Lb�2t3�T0 k� ����%�0e  51D Q $�    � 
 �Fb�� �@b�C@LDMp*|(�ÞBޯ�E
Lb�Bx3�T0 k� 3���%�0e  51D Q ��    � 
 �Fc� �@b�C@LDMp*|(�˟B޷�E$Lb�B|3�T0 k� 3���%�0e  51D Q ��    � 
 �Fc� �@b�C@PDMt)|(�ӠB޿�E(Lb�B�3�T0 k� 3���%�0e  51D Q ��    � 
 �Fc� �@b�B@TCMt)|(�סB���E0Lb�B�3�T0 k� 3���%�0e  51D Q ��    � 
 �Fc� �@b�B@XCMt(|(�ߢB���E8Lb�B�3�T0 k� 3���%�0e  51D Q ��    � 
 �Fc� �@b�A@XCMt(|(��E���E@Lb�B�3�T0 k� ����%�0e  51D Q ��    � 
 �Fc� �@b�A@\CMt(|(��E���EDLb�B�3�T0 k� ����%�0e  51D Q ��    � 
 �Fc� �@b�A@`CMx'|(��E���ELLb�B�3�T0 k� ����%�0e  51D Q ��    � 
 �Fc� �@b�@@dCMx'|(���E���D�TLb�2�3�T0 k� ����%�0e  51D Q ��    � 
 �Fc� #�@b�@@dCMx'|(A��E��D�XLb�2�3�T0 k� �|��%�0e  51D Q ��    � 
 �Fc� #�@b�@@hCMx&|(B�E��D�`Lb�2�3�T0 k� �|��%�0e  51D Q ��    � 
 �@� '�@b�?@lCM|&!�(B�D��D�hLb�2�3�T0 k� �x�|%�0e  51D Q ��    � 
 �@#� +�@b�?@pCM|%!�(B�D�#�D�pLb�2�3�T0 k� �t�x%�0e  51D Q ��    � 
 �@#� +�@b�?@pCM|%!�(B�D�+�E�tLb��3�T0 k� �p�t%�0e  51D Q ��   � 
 �@'� /�@b�>@tCM|%!�(B�D�3�E�|Lb� �3�T0 k� �p�t%�0e  51D Q ��    � 
 �@+� 3�@c >@xCM|$!�(B#�D�?�E��Lb� �3�T0 k� Cl�p%�0e  51D Q ��    � 
 �@+� 3�@c >@xCM�$!�(B+�D�G�E��Lb� �3�T0 k� Ch�l%�0e  51D Q ��    � 
 �@/� 7�@c>@|CM�$!�(B/�D�O�E��Lb� �3�T0 k� Ch�l%�0e  51D Q ��    � 
 �@3� ;�@c=@|BM�#!�(B3�D�[�E��Lb�!�3�T0 k� Cd�h%�0e  51D Q  ��    � 
 �@3� ;�@c=@�BM�#!�(B;�D�c�E�� Lb�!�3�T0 k� C`�d%�0e  51D Q  ��    � 
 �@7� ?�@c=@�BM�#!�(B?�D�o�E�� Lb�!�3�T0 k� #\	�`	%�0e  51D Q  -�    � 
 �@7� ?�@c<@�BM�#!�(RC�D�w�E��!Lb�!�3�T0 k� #\	�`	%�0e  51D Q  ��    � 
 �@;� C�@c<@�BM�"|(RK�D��Er�#Lb�!��3�T0 k� #X	�\	%�0e  51D Q  ��    � 
 �@?� G�@c<@�BM�"|(RO�D��Er�$Lb�"��3�T0 k� #T	�X	%�0e  51D Q  ��    � 
 �@?� G�@c<@�BM�"|(RS�D��Er�%Lb�"��3�T0 k� #T	�X	%�0e  51D Q  ��    � 
 �@C� K�@c;@�BM�!|(RW�D��Er�'Lb�"��3�T0 k� 3P	�T	%�0e  51D Q  ��    � 
 �@C� K�@c;@�BM�!|(R_�D��Er�(Lb�"��3�T0 k� 3L	�P	%�0e  51D Q ��    � 
 �@G� O�@c ;@�BM�!|(Rc�D��F�)Lb�"��3�T0 k� 3H
�L
%�0e  51D Q ��    � 
 �@G� O�@c ;@�BM�!|(Rg�D��F�+Lb�#� 3�T0 k� 3H
�L
%�0e  51D Q ��    � 
 �@K� S�@c$:@�BM� |(Rk�D���F�,Lb�#	�3�T0 k� 3D
�H
%�0e  51D Q ��    � 
 �@K� S�@c(:@�BM� |(Ro�D���F�-Lb�#	�3�T0 k� �@
�D
%�0e  51D Q ��    � 
 �@O� W�@c(:@�BM� |(Rs�D���F�/Lb�#	�3�T0 k� �@
�D
%�0e  51D Q ��    � 
 �@O� W�@c,:@�BM� |(bw�D���Lr�0LS #	�3�T0 k� �<
�@
%�0e  51D Q ��    � 
 �@S� [�@c,:@�BM�|(b�L��Lr�1LS#	� 3�T0 k� �8�<%�0e  51D Q ��   � 
 �@S� [�@c09@�BM�|(b��L��Lr�3LS$  3�T0 k� �4�8%�0e  51D Q ��    � 
 �@W� _�@c09@�BM�|(b��L��Lr�4LS$$ 3�T0 k� �4�8%�0e  51D Q  ��    � 
 �@W� _�@c49@�BM�|(b��L��Lr�5LS$, 3�T0 k� �0�4%�0e  51D Q  ��    � 
 �@[� c�@c49@�AM�|(b��Lp�Lr�7LS$3�3�T0 k� �,�0%�0e  51D Q  ��   � 
 �@[� c�@c88@�AM�|(b��Lp�Lr�8D�$7�3�T0 k� �,�0%�0e  51D Q  ��    � 
 �@_� g�@c88@�AM�|(b��Lp�Lr�9D�%	�?�3�T0 k� �(�,%�0e  51D Q  ��    � 
 �@_� g�@c<8@�AM�|(b��Lp#�Lr�:D�%	�C�3�T0 k� �$�(%�0e  51D Q  ��    � 
 �@c� g�@c<8@�AM�|(b��Lp+�Lr�;D�%	�G�3�T0 k� �$�(%�0e  51D Q  /�    � 
 �@c� k�@c@8@�AM�|(b��Lp3�Lr�<D�&	�K�3�T0 k� � �$%�0e  51D Q  ��    � 
 �@g� k�@c@7@�AM�|(r��Lp7�Lr�>D�&	�O�3�T0 k� #� %�0e  51D Q  ��    � 
 �@g� o�@cD7@�AM�|(r��Lp?�L��?D�'
S�3�T0 k� #�%�0e  51D Q  ��    � 
 �@g� o�@cD7@�AM�|(r��LpG�L��@D� '
W�3�T0 k� #�%�0e  51D Q  ��    � 
 �@k� s�@cH7@�AM�|(r��LpO�L��AD� (
[�3�T0 k� #�%�0e  51D Q  ��    � 
 �@k� s�@cH7@�AM�|(r��L�W�L��BD�$)
_�3�T0 k� #�%�0e  51D Q  ��    � 
 �@o� s�@cL7@�AM�|(r��L�_�L��CD�()
c�3�T0 k� ��%�0e  51D Q  ��    � 
 �@o� w�@cL7@�AM�|(r��L�c�L��DD�()	�g�3�T0 k� ��%�0e  51D Q  ��    � 
 �@o� w�@cP8@�AM�|(r��L�k�L��ED�()	�g�3�T0 k� ��%�0e  51D Q  ��   � 
 �@s� w�@cP8@�AM�|(r��L�s�L��FD�(*	�k�3�T0 k� ��%�0e  51D Q  ��    � 
 �@s� {�@cT8@�AM�|(r��L�{�L��GD�,*	�o�3�T0 k� ��%�0e  51D Q  ��    � 
 �@s� {�@cX8@�AM�|(r��L��L��HD�,+	�o�3�T0 k� � �%�0e  51D Q  ��    � 
 �@w� �@cX8@�AM�|(B��L���L��ID�,,ss�3�T0 k� � �%�0e  51D Q  ��    � 
 �                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��1b ]� z y � ����x�    
    � �R    ���� �    �| �   	            �   '             `     ���   0
%          ���    �	    � 3I�    ���� 3<m    �� �                    R �          
@     ���   0
 
          H=�         ���     H2� ���     ��   	               �         ��     ���   8

           @7�   $ $       Ej�     @7� E].       �                  A�$          ��      ���   8          K�   $ [     .�l�     O��l�+    �� X                  �$                ���   P
		          �Z  ��	     B�
[6     �Z�
[6                             ���K              L  ���    P              I�      V �}�     I�F �`    W�                 Z �         P      ��H   8
           Q� M M     j �V�     P�� ��S    �                W  Z �          ۀ�     ��@ 0	
           eN� � �	   ~ Ӌ�     ea� Ӂ�    �� �              T Z ��        ��     ��`   0	           U;�   
    � ΢R     U;� ΢R                       	 Z �         	 �     ��@  H
            A��  � �	   � �ݑ     ?�� �$�    ��h                	 Z �         
 �`�     ��@ 0
 		          � ��     �Q�     ��E�     P �                       �c             �  ��@    		 5                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          XT  ��        � �l�     W�I �N=    W� "                x                j  �       �                          X    ��        � �       W   �                                                               �                          � 3 � E�l�
 � � � � ��� � �                	 

     C ��  �o�C       �d �r@ �d s@ �$  t� �d `u  �$ u� �D 0u� �� v@ E� v`���. ����< ����J ����X � �� t  A$ b@ � �r@ � s@  _  /� _  /� _  0 _@ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π 
�< U� 
�� V  
�| V  
�\ V� 
�� V� 
�\ W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� �  
���4  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"     
�j,� B �
� �  �  
�  I    ��     � �      ��    ��     � �       I    ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �%      ��2T ���        � �T ���        �        ��        �        ��        �      ��      y p��        ��                         ��q < 		��� �                                    �                 ����            I ����%��   
 � 2 F��            16 Pat Verbeek ov n    0:01                                                                        4  4      �]C-m C"% �kj@ � krP �k�@ � k�P �c�( �	c�( � 	�> �
c�0 � c�@ � c�H �k~Z �k�R � k�Y �k�R �k�O � �J � �I �cV< � c^L �J� � �K5 �K% �c� � �c� �c� � � c� �	� � �	� � �� � � � �!"�3 � ""�E �#�/ �$
�> �%"� � � &"� � �'"� � �(*� � �)"�3 � *"�E �+�/ � 
�> �-�/ � 
�> � 
�> �0�. � 
�= t  *Q~ t  *Q~ t  *Q~ t  *Q~^  "O �\  "O �Z  "O �Y  "O �`  "H �^  "K �U <"C �] ="G �]  "K �U  "C �                                                                                                                                                                                                                         �� R @ �     �     @ 
         b     Q P E ]  ��                    	 �������������������������������������� ���������	�
��������                                                                                          ��    �@g�� ��������������������������������������������������������   �4, .  $ " L���*��@� @���A&�                                                                                                                                                                                                                                                                                                                                       �� ����"                                                                                                                                                                                                                                     O    0    ��   D�J    	  ��  	                           ������������������������������������������������������                                                                                                                                         �      �      �                �  �          	  
 	 
 	 	 ��������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� ���������������������             �                   �    (      �  K
�J      "a                             �������������������������������������������������������                                                                                                                                    �                    :�      � �� �          	 	 
  	 
 
 ������ ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ������            x                                                                                                                                                                                                                                                            
                                                 �             


             �  }�         ����������������  '|������������  '|����������������    ����������������  +����   ��������������������        +                                                    'v                  ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 0 I =               	                  � 2��� �\        �c�b7.P�1sc$                                                                                                                                                                                                                                                             )n)n
  �                        c                  `      l                                                                                                                                                                                                                                                                                                                                                                                                                            > �  >�  @�  (�  (�  J`�  ���������N�����#����� �����U����[�����[�                       ���         	�	�   & AG� U ��   	              �                                                                                                                                                                                                                                                                                                                                      p B F             -             !��                                                                                                                                                                                                                            Y��   �� �� �      �� @ 	     ��������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� ��������������������������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ������             $�������������������������������������������������������f��ff�fff�������Ƭffffffff�fff�fffffffffl�����̚�lfl��ffl�fffflffffffffff����������������ʺ��k���jY��f���������������������������������������������������������������������ff��ff�fff�ffU�ffU�fƪfffffffffffhffffʗuZUUXYUw��fffffffffff�zVffhVfffffffffffffkffffffffi�ffffk�fff�fffɖffjvffkfflfffffffff����������������������������ʫ����������������������������������ffffffffffff�f��f���kYk��{l��zff�jfƶfffl������������������y����lfff����˘���fff����x����f˘ffj�f�ff�l�fWf�f��li���j��f���f�UZ��j���ʫ������������������������������������������������������������lf���f���f�u����l��Yk���l���l�f�w��kW�fjww��W�������W���uw��x�f��w˘wWX�uww�xw�x���xx��wwx�wWxwZ̪{h��yŌ����X������U˙�u���W�������������������������������������������������������������������˪�Ǜʫņj�u�k�Z�ƫ�����W�������l���l��̨�������flˬ��l����k�̇wux��Uwwwww��Wx�����W������������U�Xʅ�zʨ��ʈ���W���u�̺u���YU������������������������̪���flƪ��������������f��ff�fff�fffffff���������fflffffffffffffffffffff�l���f���fk�lfffflffff�ffff�ffffww�����������ʫ�ffjWfkUz�U��������Y��u�xuX�wX��u�x�u�W�u�w�uwx�WZ�ffU�ffu��f�vvf�V�f�V�f�V�f�V�flI    B      8      W                       B     �   ����������      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$     $�   ���$� >�������� J  �� ��� ���� ��� �$ ^$   �   ����� ��  ����� �$ ^$  4  �  �� . 
e�     � ���   �� � ��� �� � ��� � �97 �9��7  �      �      )�����������J  g���        f ^�         �� � 
      )      ��1��������J���J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  "!    " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """""" "!   " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  "!    " ""  !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �           �  � ���� "            �  ��  �                                     �  �       �            "  �"     �                  ���� ��� ����                            �   O   T     ��                                 � ���� ��   � � �                                                                                                                                       0 0#0  03  10         �  �  � 
�� ��} ˚w
���	����+� �+� ��� ",  "�  ". 34 DC3 DD3 �DC ��  ��  
"   "  "  ""  "!    �                    �   �   �   w   m�  g�� z�� ����̹���˙�̼̰������������蜚��L��>\���" ""  ""  �+ "	��"� �����.�"��"! "  ��           /   ��  �   �    �  ���  ��� ��  �                        �   �   �                                           �    ���  ��                    ��  ��  ��� ���                                                                                                                                                                                                                   	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                       "   "  !�    ��                              �                        ���� ��� ����                      �  �� ��  �    � ���                                                                                                                                                                                                  �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �    �  ��  �                                     �  �       �            "  �"     �                       �������  ���    �                    ��  ��  ���                                                                                                                                                                                                                
  �  ̈ �� ,�  ""   "                       �������݅]̻�U�˅U3�U\�BU\�3 "��",�"��"��� ��  �             ݽ���۹����" ��" ��"��".�  �"  �/� .���" � ��              �   .   �   � � �� �� ��                    ��  ��  ���            � ˹ Y�����
�ڛ��٩ �� �̽���ݪ۽w�}�֪�vv���p���   �  ��"� ��� "                         �  �                         ���� ��� ����                � ��                    ���� �                                                                                                                                                                                              �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �      �  �  �  �  �  �   �                                              �   �                                                                                                                                                                                                                              �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                /���"/�  ��                    �                                                                            �               �  �  ��  �   �   �       ���                                                                                                                                                                                              ˰ ̻ ̻ �� {�  �� 
�� ��� ��� ������
���	��ܻ̍ݻ���"� 8"  8  �  D�  H�  X�  ��  �   �          "  "     �                        ��  ��� �̺�̻����ۻ�˽��̽��̝ ̙� �30 �EP �U@ �T0 EC0 T3  C:  K�  �"  �"/ ����˽� �"� "" �""� � �� ��      �   �� ��  �"  �                   
 "� ""� ""� "                       �                             ���                         �  ��                    �����                      ��  �  �  �   �                                                                                                                                                                                            � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �                          � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         �w
���̩ۚ,���+��   �   �   �   �  �  9  D3  D2 T2 DB DB �@ ��  ��  ��  �  "" ""�"!��" ��       �                w�  ��� ��� ��� ˼����ɀ�؊�˽ـ��˰��̰�̻@"���"+H�"$X�"$�@"E� U� E� D� ,˸  ��  ��  ,� "" �"" """�"!���� � �              �         �           �       �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                    �     �                         � ���� ��   � � �                                                                                                                                                �  ɪ ̹� ˫�ɫ��˙�̽ۻۻݽ���Xۼ"�C3"�T32�SD3UCDT0 3C  0  �   �  +  "  "   ����                     �� �� �� ��w ��& �vv ��p ̽  ̽  ��  ؠ  ��  (�  �"  �� 3"��3 �3  ��   �   �       "   "     ���                            
   Z   �  
�  
�  ��  ɍ ʠ "� "  ""� "� ��  ��                  �   �                        ���                         �  ��                    �����                                                                                                                                                                                                                                              �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                                               �         �  �� �  �� ��                                                                                                                                                   �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDD