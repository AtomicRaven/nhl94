GST@�                                                           �B     ��                                                        �� s ��  �         �������J���x������������������        *c     #    ����                                d8<n    �  ?    @�����  �
fD�
�L���"����D"� j   " B   J  jF�"    "�j* ,  �����
�"     �j@ �    ��
                                                                                  ����������������������������������     � ��    = a0 U1 210 .*  &  ӟ  � �  	  	           4� 4� 4� 4�                 �EE 1         =:;�����������������������������������������������������������������������������������������������������������������������������    UU  11  ..    &&   ��    ��  ��                  44  44  44  44                  n�  !!          :: �����������������������������������������������������������������������������                                �   N       �   @  &   �   �                                                                                 ' 1�EE  !n!�    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E N �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ^@&A]��@��\0` k�\��A 6L_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_\�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_\�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6K�_\�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6K�_\�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6K�_\�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6K�_\�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6K�_\�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6K�_\�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6K�_\�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6K�_l�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6K�_l�fL�P��W"s�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6K�_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6K�_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6K�_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6K�_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6K�_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6K�_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6K�_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6L_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6L_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6L_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6L_l�fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6L_l�fL�P��W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��L� 6L_l�fL�P��W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��L� 6L_l�fL�P��W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��L� 6L_l�fL�P\�W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��L� 6L_l�fL�P\�W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��L� 6L_l�f<�P\�W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��L� 6L_l�f<�P\�W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��L� 6L_l�f<�P\�W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_l�f<�P\�W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_l�f<�P\�W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_l�f<�P\�W"��T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_l�f��P\�W3�T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_l�f��P\�W3�T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_l�f��P\�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��P\�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��P\�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��P\�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_l�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_\�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_\�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_\�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_\�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_\�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_\�f��Pl�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6L_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��Pl�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P\�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P\�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P\�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P\�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P\�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P\�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��L� 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��L� 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��L� 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��L� 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��L� 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��L� 6A_��f<�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��L� 6A_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6A_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6A_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6A_��fL�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6A_��fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6A_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6A_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6A_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6A_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6A_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6K�_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6K�_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6K�_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6K�_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6K�_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\��A 6K�_\�fL�P��W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\"[��A 6K�_\�fL�P\�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\"[��A 6K�_\�fL�P\�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\"[��A 6K�_\�fL�P\�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\"[��A 6K�_l�fL�P\�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\"[��A 6K�_l�fL�P\�W3�T0 k� ������U8D"!U2d    %�O 	   � &�8^@&A]��@��\0` k�\"[��A 6K�_l�fL�P\�W3�T0 k� ������U8D"!U2d    ��O 	   � &�8^@&A]��@��\0` k�\"[��A 6K�_l�fL�P\�W3�T0 k� ������U8D"!U2d   ��O 	   � &�8^@&A]��@��\0` k�\"[��A 6K�_l�fL�P\�W3�T0 k� ������U8D"!U2d   ��O 	   � &�8VGAP@�P `|  A`@ A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|  A`@ A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|  A`@ A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|  A`< A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|  A`< A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|  A`8 A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|  A`4 A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|$ A`4 A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|$ Ap0 A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|$ Ap, A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|$ Ap( A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|$ Ap$ A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|$ E�  A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|$ E� A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|$ E� A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|$ E� A ���PT0 k� ������U8D"!T2d    ��V    �  ��VGAP@�P `|$ E� A ���PT0 k� ����U8D"!T2d    ��V    �  ��VGAP@�P `|$ E� A ���PT0 k� ����U8D"!T2d    ��V    �  ��VGAP@�P `|$ E�� A ���PT0 k� ����U8D"!T2d    ��V    �  ��VGAP@�P `|$ E�� A ���PT0 k� ����U8D"!T2d    ��V    �  ��VGAP@�P `|$ A�� A ���PT0 k� ����U8D"!T2d    ��V    �  ��VGAP@�P `|$ A��A ���PT0 k� ����U8D"!T2d    ��V    �  ��VGAP@�P `|$ A��A ���PT0 k� ����U8D"!T2d    ��V    �  ��VGAP@�P `|$ A��A ���PT0 k� ����U8D"!T2d    ��V    �  ��VGAP@�P `|$ A��A ���PT0 k� ����U8D"!T2d    ��V    �  ��VGAP@�P `|$ A��A ���PT0 k� ����U8D"!T2d    ��V    �  ��VGAP@�P `|$ E_�A ���PT0 k� ��
��
U8D"!T2d    ��V    �  ��VGAP@�P `|$ E_�A ���PT0 k� ����U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_�A ���PT0 k� ����U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_�A ���PT0 k� ����U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_�A ���PT0 k� �� �� U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_�A ���PT0 k� �� �� U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_�A ���PT0 k� ������U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_�A ���PT0 k� �w��{�U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_�A ���PT0 k� �o��s�U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_�A ���PT0 k� �g��k�U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_�A ���PT0 k� �_��c�U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_t	A ���PT0 k� �P �T U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_l	A ���PT0 k� �H �L U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_d
A ���PT0 k� �@ �D U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_\
A ���PT0 k� �8�<U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_T
A ���PT0 k� �0�4U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_DA ���PT0 k� � �$U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ E_<A ���PT0 k� ��U8D"!T2d    ��V 	   �  ��VGAP@�P `|$ EO4A ���PT0 k� � � U8D"!T2d    ��V 
   �  ��VGAP@�P `|$ EO,A ���PT0 k� ����U8D"!T2d    ��V 
   �  ��VGAP@�P `|$ EOA ���PT0 k� ������U8D"!T2d    ��V 
   �  ��VGAP@�P `|$ EOA ���PT0 k� ������U8D"!T2d    ��V 
   �  ��VGAP@�P `|$ EOA ���PT0 k� ������U8D"!T2d    ��V 
   �  �}VGAP@�P `|$ EN�A ���PT0 k� ������U8D"!T2d    ��V 
   �  �zVGAP@�P `|$ EN�A ���PT0 k� ������U8D"!T2d    ��V 
   �  �wVGAP@�P `|$ A�A ���PT0 k� ������U8D"!T2d    ��V 
   �  �tVGAP@�P `|$ A�A ���PT0 k� ������U8D"!T2d    ��V 
   �  �qVGAP@�P `|$ A�A ���PT0 k� ������U8D"!T2d    ��V 
   �  �nVGAP@�P `|$ A�A ���PT0 k� ������U8D"!T2d    ��V 
   �  �kVGAP@�P `|$ A�A ���PT0 k� ������U8D"!T2d    ��V 
   �  �iVGAP@�P `|$ A�A ���PT0 k� ������U8D"!T2d    ��V 
   �  �gVGAP@�P `|$ A�A ���PT0 k� �s��w�U8D"!T2d    ��V 
   �  �dVGAP@�P `|$ EޤA ���PT0 k� �s��w�U8D"!T2d    ��V 
   �  �aVGAP@�P `|$ EޜA ���PT0 k� �l�pU8D"!T2d    ��V 
   �  �_VGAP@�P `|$ EޔA ���PT0 k� �h�lU8D"!T2d    ��V 
   �  �\VGAP@�P `|$ EބA ���PT0 k� �\�`U8D"!T2d    ��V 
   �  �YVGAP@�P `|$ E�|A ���PT0 k� �T�XU8D"!T2d    ��V 
   �  �VVGAP@�P `|$ E�tA ���PT0 k� �L�PU8D"!T2d    ��V 
   �  �TVGAP@�P `|$ E�lA ���PT0 k� �D	�H	U8D"!T2d    ��V    �  �RVGAP@�P `|$ E�\A ���PT0 k� �4	�8	U8D"!T2d    ��V    �  �PVGAP@�P `|$ E�T
A ���PT0 k� �,	�0	U8D"!T2d    ��V    �  �NVGAP@�P `|$ E�L
A ���PT0 k� �$	�(	U8D"!T2d    ��V    �  �LVGAP@�P `|$ E�D
A ���PT0 k� �	� 	U8D"!T2d    ��V    �  �JVGAP@�P `|$ E�4
A ���PT0 k� �	�	U8D"!T2d    ��V    �  �HVGAP@�P `|$ E�,
A ���PT0 k� �	�	U8D"!T2d    ��V    �  �GVGAP@�P `|$ E�$
A ���PT0 k� ��	� 	U8D"!T2d    ��V    �  �FVGAP@�P `|$ E�
A ���PT0 k� ��	��	U8D"!T2d    ��V    �  �EVGAP@�P `|$ E�	A ���PT0 k� ��	��	U8D"!T2d    ��V    �  �DVGAP@�P `|$ E�	A ���PT0 k� ��	��	U8D"!T2d    ��V    �  �CVGAP@�P `|$ E]�	A ���PT0 k� ����U8D"!T2d    ��V    �  �BVGAP@�P `|$ E]�	A ���PT0 k� ����U8D"!T2d    ��V    �  �AVGAP@�P `|$ E]�	A ���PT0 k� ����U8D"!T2d    ��V    �  �@VGAP@�P `|$ E]�	A ���PT0 k� ����U8D"!T2d    ��V    �  �?VGAP@�P `|$ E]�	A ���PT0 k� �� �� U8D"!T2d    ��V    �  �>VGAP@�P `|$ E]�	A ���PT0 k� �� �� U8D"!T2d    ��V    �  �=VGAP@�P `|$ E]�A ���PT0 k� ������U8D"!T2d    ��V    �  �<VGAP@�P `|$ E]�A ���PT0 k� ������U8D"!T2d    ��V    �  �;VGAP@�P `|$ A]�A ���PT0 k� �� �� U8D"!T2d    ��V    �  �:VGAP@�P `|$ A]�A ���PT0 k� �p�tU8D"!T2d    ��V    �  �9VGAP@�P `|$ A]�A ���PT0 k� �d�hU8D"!T2d    ��V    �  �8VGAP@�P `|$ A]�A ���PT0 k� �P�TU8D"!T2d    ��V    �  �8VGAP@�P `|$ A]�A ���PT0 k� �H�LU8D"!T2d    ��V    �  �8VGAP@�P `|$ A]�A ���PT0 k� �@�DU8D"!T2d    ��V    �  �8VGAP@�P `|$ A]xA ���PT0 k� �8�<U8D"!T2d    ��V    �  �8VGAP@�P `|$ A]pA ���PT0 k� �0�4U8D"!T2d    ��V    �  �8VGAP@�P `|$ A]dA ���PT0 k� �$�(U8D"!T2d    ��V    �  �8VGAP@�P `|$ A]\A ���PT0 k� �� U8D"!T2d    ��V    �  �8VGAP@�P `|$ A]XA ���PT0 k� ��U8D"!T2d    ��V    �  �8VGAP@�P `|$ A]PA ���PT0 k� ��U8D"!T2d    ��V    �  �8VGAP@�P `|$ A]DA ���PT0 k� ��U8D"!T2d    ��V    �  �8VGAP@�P `|$ E�<A ���PT0 k� ��U8D"!T2d    ��V    �  �8VGAP@�P `|$ E�4A ���PT0 k� � �U8D"!T2d    ��V    �  �8VGAP@�P `|$ E�0A ���PT0 k� � �U8D"!T2d    ��V    �  �8VGAP@�P `|$ E� A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `|$ E�A ���PT0 k� ��
��
U8D"!T2d    ��V    �  �8VGAP@�P `|$ E�A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `|$ E�A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `|$ E��A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `|$ E��A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `|$ E��A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��	A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��	A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��
A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��A ���PT0 k� ����U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��A ���PT0 k� �� �� U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��A ���PT0 k� �� �� U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��A ���PT0 k� ��"��"U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��A ���PT0 k� ��#��#U8D"!T2d    ��V    �  �8VGAP@�P `�$ E��A ���PT0 k� ��#��#U8D"!T2d    ��V    �  �8VGAP@�P `�$ E�|A ���PT0 k� ��$��$U8D"!T2d    ��V    �  �8VGAP@�P `�$ H�pA ���PT0 k� �t%�x%U8D"!T2d    ��V    �  �8VGAP@�P `�$ H�lA ���PT0 k� �d%�h%U8D"!T2d    ��V    �  �8VGAP@�P `�$ H�dA ���PT0 k� �T%�X%U8D"!T2d    ��V    �  �8VGAP@�P `�$ H�`A ���PT0 k� �L&�P&U8D"!T2d    ��V    �  �8VGAP@�P `�$ H|TA ���PT0 k� �<#�@#U8D"!T2d    �V    �  �8VGAP@�P `�$ H|LA ���PT0 k� �4!�8!U8D"!T2d    ��_    �  �8VGAP@�P `�$ H|HA ���PT0 k� �, �0 U8D"!T2d    ��_    �  �8VGAP@�P `�$ H|@A ���PT0 k� �(�,U8D"!T2d    ��_    �  �8VGAP@�P `�$ Hl8A ���PT0 k� ��U8D"!T2d    ��_    �  �8VGAP@�P `�$ Hl0A ���PT0 k� ��U8D"!T2d    ��_    �  �8VGAP@�P `�$ Hl,A ���PT0 k� ��U8D"!T2d    ��_    �  �8VGAP@�P `�$ Hl$A ���PT0 k� � �U8D"!T2d    ��_    �  �8VGAP@�P `�$ HlA ���PT0 k� ����U8D"!T2d    ��_    �  �8VGAP@�P `�$ HlA ���PT0 k� ����U8D"!T2d     �_    �  �8VGAP@�P `$ Hl A ���PT0 k� ��#;P U8D"!T2d  �_    �  �8VGAP@�P `$ Hl!A ���PT0 k� ��#;P U8D"!T2d  ��_    �  �8VGAP@�P `$ Hl"A ���PT0 k� ��#;P U8D"!T2d  ��_    �  �8VGAP@�P `$ Hk�"A ���PT0 k� ��#;P U8D"!T2d  ��_    �  �8VGAP@�P `$ Hk�#A ���PT0 k� ��#;P U8D"!T2d  ��_    �  �8VGAP@�P `$ Hk�$AP���PT0 k� ��#KP U8D"!T2d  ��_    �  �8VGAP@�P `$ Hk�$AP�P0PT0 k� ��#KP U8D"!T2d  ��_    �  �8VGAP@�P `$ Hk�%AP0P0PT0 k� ��#KP U8D"!T2d  ��_    �  �8UcQAP@�P `$ BK�gL@��a��lAPT0 k� ��#kP U8D"!T2d   ��_    �  �8^@&A]��@��\0` k�\��A 6L_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O 
   � &�8^@&A]��@��\0` k�\��A 6L_��f\�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�f\�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�f\�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�f\�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�f\�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_\�f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_\�f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_\�f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_\�f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_\�f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_l�f��M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f��M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f��M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f��M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f��M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f��M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f��M��V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f��M��V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f��M��V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M��V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M��V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�M\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_l�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_\�f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��M 6A_��f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f�Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��L� 6A_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��L� 6A_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��L� 6A_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��L� 6A_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��L� 6A_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��L� 6A_��f��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��L� 6A_��f ��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��A 6A_��f ��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��A 6A_��f ��Ml�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��A 6A_��f ��Nl�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��A 6A_��f ��Nl�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"k��A 6A_��fL�Nl�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��fL�Nl�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��fL�Nl�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��fL�Nl�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��fL�O\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��fL�O\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��fL�O\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��fL�O\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f\�O\�V3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f\�P\�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f\�P\�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6A_��f\�P\�W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6A_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6A_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6A_��f ��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6A_��f ��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6A_��f ��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6K�_��f ��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6K�_��f ��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6K�_��f�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6K�_��f�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6K�_��f�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\"K��A 6K�_��f�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6K�_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f\�P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8^@&A]��@��\0` k�\��A 6L_��f��P��W3�T0 k� ������U8D"!U2d    ��O    � &�8                                                                                                                                                                            � � �  �  �  c A�  �J����  �     � \��z ]���-w � �  �          �X4�    �Q�X`F    ��q   ��          
    ��         !�       ��� (           �d         �  �-    ��d  �-                          	   �         �P  �  ���  8�            ��          %�    ���  %�                          � ��                 ��� 	@	            ��             $2    �  �d    ���   ��          A�$          �  �  ��� @ H$
           �j           .  �Q    ��  �    ���   ��         ��$          �  �  ���   H
	!           ��  ��
     B�	5�      ���	5�                              ���              �  ���      0              Z $ $     V��)�     gYE��)U                  Z�8          �`     �H   8            ʪ � �     j  �4    �W�  !f    ���   MM       Z�8        ڰ�    ��`   0
% 
            �i  : :    ~�6     a���6     ;     ��      	 Z�8         `�    ��@   0            ��  : �	   ���h    �XO���    p�?   ��        Z�8         	 ��    ��@   8           �  � �    ��Z�     A��[�    R�D   ��      S
 Z�8         
 	��    ��`   P
		           =&  �
     �  No    ��"  ơ    ���   	�	�               ���M                ��B    P                   ��      �                                                                           �                               ��        ���          ��                                                                 �                           ��  ��        ���Jk     ����Jk         "                 x                j     �   �                             � 66      ���   �x    ��   ��    s�                                      .        �                                                             	    
         
        ��  �W�       
�| V� 
� V� 
�\ W  
�< W� 
�� W� 
�\ W����J ����X � �D v` $ `o� � p�  p� �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� 
�< W� 
�� W� 
�\ W����� � 
�< V� 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����8��        ������  
�fD
��L���"����D" � j  "  B   J jF�"    "�j * , ����
��"     �j @�    �
� �  �  
�     ��     ��  �        ��     ��	            ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �_   0      �� T ���        �6T ���        �        ��        �        ��        �    ��
    ^�� �        ��                         �w� $ * ���                                    �                ����         
   � ���%��$    �8��          �    16 Verbeek  uk  on     5:17                                                                        2  5     �"(c�<"�DT
t"��*�D2X=2	P]2	
l}~D �" � � " � � " � � "M �  *NO �*P �  )�` � c�G*"� �* "�
"� �*� �@"�_@ "�q0�W0
�f@ "G x@  *G�X  *KxX  *HxH  *PxX  *HxH "*PxX  *HxH $*PxX  *Hx �&J� z � 'J� z �(B� � � )B� G*"�.G +"�@7,"�&7-*�53."�3 /"�#0� #1
� � 2*Oz � 3*BzH  *PRH  *PRH  *PRX  *KRX  *KRX  *KR � 
�	 z;"H �  *Hx �  *Hx �>b` � � b^ �                                                                                                                                                                                                                         4� � T                  %� �     G P E Z  ���� U               	�������������������������������������� ���������	�
��������                                                                                          ��    �*~���� ��������������������������������������������������������   �4X .  * $� ���� �	�)��@��ӂ��,�                                                                                                                                                                                                                                                                                                                                ��+                                                                                                                                                                                                                                         
      I  	      ��  H�J      7�  	                           ������������������������������������������������������                                                                                                                                         �        �      �        �    p�           
 	  
	 
 	 	 ����������� ���� ������ � ����������� ��� � ���������� ������������������������ �������� ��������������� ������������������������������������������ ������������� ��� ���������� ����������������������������� ��������������� ����                                  =    *        D�J    	 wu                             ������������������������������������������������������                                                                   
                                                                     �     �      �        �        �  �          	  
 	 
 	 	 ��� ������� ������ �  ��� �� ����� ������������������������������������������������ ��� �����  ���� ������������� ������������������� ����������� ����  ���������� ������������������  ������������������� �� ����� ��� ���������� �            �                                                                                                                                                                                                                                               
                                                            �             


             �`  }�          �#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 6 F 8                	                 � CPŷ �\                                                                                                                                                                                                                                                                                  �  1�EE  !n!�              k                              k                                                                                                                                                                                                                                                                                                                                                                                                    j   'M
  . .7 2 5 ?Lpj   u�  �����^�����$�����q�����D�����[����UE����ˣ        <  ���@ : / z        	  	�   & AG� �   �   
           �Z�                                                                                                                                                                                                                                                                                                                                    p C B   �      ��               !��                                                                                                                                                                                                                            Y   �� �� Ѱ       �� ?      ����������� ���� ������ � ����������� ��� � ���������� ������������������������ �������� ��������������� ������������������������������������������ ������������� ��� ���������� ����������������������������� ��������������� ������� ������� ������ �  ��� �� ����� ������������������������������������������������ ��� �����  ���� ������������� ������������������� ����������� ����  ���������� ������������������  ������������������� �� ����� ��� ���������� �   ��      $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    4      >   �                         f     �  �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f      �� |���� ���� |���� �$     �f ��     �f �$ ^$ �@       �       �     �   z 
� � v           
  �   ��  
  �   �$ ^$ x      ���  �  ��   ��   s ������J
  ����� c ���� ^�       ��   s    �   �       ���� 
�*�����������     �  �   �      ���v��� 
�*���� 1| r� ^  ��  yf  y<  ��������������������������������GvdDGw6wGwcfGwsfGwv6Gww6GwwcGwwcDDDDwwwwffffffffffffffffUUUUttttDDDDwwwwffffffffffffffffUUUUtttwN���t���wN��wt��wwN�wwt�wwwNwwwtGwweGwwU�tvf�wff�Fff�Fff��df��ffwwwwUUUUffffftDDft33gt5egt6Vgt5gwwwwUUUUffffDDDD3333eeeeVVVVwwwwwwwwUUUUffffDDFF35FfefDDVVFUufGfwwwwGwwwGwwwUUUUffffDDDDUUUUffffwwwwwwwuwwwuUUUUffffDDDDUUUUffffwwwwUUUUffffddDDfd33DD6VUd5eft6WwwwwUUUUffffDDGf35GfVVGvefGv6VGvwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwN�Fft�FfwN�dwt�fwwNGwwtGwwwDwwwtwt6Wwt5gwt6Wwt5gwt6Wwt5gtt6Wwt5gDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD6VGd5fGd6VGd5fGd6VGd5fGd6VGd5fGdFt5gFt6WFt5gFt6WFt5gFt6WFt5gFt6W5fGw6VGw5fGw6VGw5fGw6VGw5fGG6VGwgwwwvwwwwgwwwvwwwwgwwwvwwwwgwwwvGt6WGt5gDt6WDt5gND6WNt5gNt6WNt5g6VGd5fGf6VGw5fDD6VGU5fGf6VGf5fGfDDDDffffwwwwDDDDUUUUffffffffffffFt5gft6Wwt5gDD6WUt5gft6Wft5gft6W5fGt6VGt5fGD6VGD5fD�6VG�5fG�6VG�GwwwDwww�Gww�Dww~�Gww�Dww�DGw~�DNt6SNt5fNt6VNteeNwFVNwteNwwFfffd3333ffffVVVVeeeeVVVVeeeeffffDDDD333DffcDVVSDeecDVVSDeecDfVSDFecDUUUUDDDDDDDDDDDDDDDDDDDDDDDDDDDDD333D6ffD6VVD5fdD6VDD5fDD6VDD5fD3333ffffVVVVDDDD33335UUU5Vff5VDD3333ffffVVVVDDDD3333UUUUffffDDDD6VGfefGfVVGwDDDD3333UUUUffffDDDDffffffffwwwwDDDD3333UUUUffffDDDDft5cft6Vwt5eDDDD3333UUUUffffDDDD3333ffffeeeeDDDD3333UUUVffeVDD5V333DffcDeecDF6SDD5cDD6SDD5cDD6SDD333D6ffD5eeD6VVD5eeD6VVD5ffD6Vd5fG�fVG�efG�VVG�edw�VGw�dww�Ffffffffwwwwwwww����DDDDNNDD��������gwwwwwwwwwww��wwDDGwDDDw��DG���Dwwwwwwwwwwwww~��wwn�wwvwwwwgwwwvFfffFfffCeeeCVVVCeeeCVVVCeeeCVVVfDDDfDDDfDDDVDDDfDDDVDDDfDDDVDDDDfSDD5cDD6SDD5cDD6SDD5cDD6SDD5cDD6VDD5fDD6VDD5fDD6VDD5fDD6VDD5fD5VDD5VDD5VDD5VDD5VDD5VDD5VDD5VDDDDDDDDDADDDADDDDDDDDDDDADDDADDDDDDDDDDDDDDwDDDDDDDDDDDDDwDDDDD5VDD5VDD5VDD5VDD5VDD5VDD5VDD5VD5cDD6SDD5cDD6SDD5cDD6SDD5cDD6SDDDDfDDDfDDD5DDD6DDD5DDD6DDD5DDD6fffdfffdeeedVVVdeeedVVVdeeedVVVdCeeeCVVVCeeeCVVVCeeeCVVVCeeeCVVVfDDDVDDDfDDDVDDDfDDDVDDDfDDDVDDDD6SDD5c3D6VfD5eeD6VVDVffDDDDDDDDDDDD3333ffffeeeeVVVVffffDDDDDDDDD6VD35fDffVDeefDVVVDfffDDDDDDDDD5VDD5VDD5V335UUU5UUU5UUUVfffDDDDDDDDDDDD3333UUUUUUUUUUUUffffDDDDDD5VDD5V335VUUUVUUUVUUUVffffDDDDD5cDD6S3D5ffD6VVD5eeD6ffDDDDDDDDD5fD36VDfefDVVVDeefDfffDDDDDDDDDDDD5DDD6DDD5DDD6DDD5DDD6DDD5DDD6eeedVVVdeeedVVVdeeedVVVdeeedVVVdwwww�twwww~ww�w�wtwwtwwww~w�wwwwDDDDDDDDDADDDDDADDDDDDDDDDDtDD4DDqt4DDDD4DDsDDDDDDDDDDDD7AtCADADDADADDDDDDDADDDADDADqDADqDDDDDADDDADDDAADAADqADDAGADDDDwwwywww�www�www�www�www�www�www�������������������������www�www�www�www�www�www�www�www����������������������!�����!�-����������!-�����������!�����wwwwwwwtwwwOwww�wwt�ww�wwOGww�D��������������-��������������������������!����������-������NNNNNNNNNNNNN���FfwfDDDDDDDDDDDDNNNDNNNDNNND����gvftDDDDDDDDDDDDwts"wwB2ww22ws#Cws#4ww2twws�www�www�www�www�www�www�www�wwwywwww��������wwww������!��������wwwwww��w��w2��w���w��t���(�wy���������y���w�����y��Gwwwwt33Dt343CeeeCVVVEeeetVVVvEee�DVVzDFf�DDDfDDDVDDDe333VfffeeeeVVVVffffDDDDDDDDDDDD3333ffffeeeeVVVVffffDDDDDDD5DDD6333efffVeeeeVVVVffffDDDDeeedVVVdeeedVVVGeedgVVDzfdD�DDD�Df��NvDGN�DNN�DND~DGD��NDNt�DDDN#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFw"GC42wsDCwt�Cwt��ws�DGt�T7DfEGt{�Gwz��w���wt�Gw��wt�Gw�wtw�{�Gww��w��w2��w���w��w���x�wy����wwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wt3Gwt4wCGGttwG4�twO�wGt�GwE��wTfNw~D�����������������DD��ww�N��D�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wfuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGy�wwy�wtw�wOw�w�w�D�w2?�wCOGww�Dwwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGww23ws""wr22w244w#tD�t3~�}�ww}O3#�w""7w##'wCC#wDG2w3G~������wwwwVtwwUvwwenwwvWwwv�wwtwwtGww�3#�w""7w##'wCC#wDG2w3G~��7���wwww}�ww}�ww}�www�www}www}wwwwwwwr��ww��ww���w4��w��ww��www}ww'r'ww"GCw2wswCwtwCwtw�wswDGtwB'tww"w#w�2w�3w�3wG4wtGDwww"wr!r'wrwuUUG4wwD4wwCtwwCtww7tww7twwGtww8�3�3�3�8�3�3�33333"2#333"33UUUUwwwtwwwtwwwtwwwtwwwtwwwtwwwt��33�?33�?33�?333333#23323#3UUUUwwwwwwwwwwwwwfgvwwwwwwwwwwwwUUUUwwwtwwwtwwwtfwfdwwwtwwwtwwwtUUUUwwwwwwwwwwwwwwwwwwuwwwWwwwwwUUUUwwwWwwwWwwwWwwuwwwuwwUuwwwUwC�38C838C�38C833C332C"33C2#3UUUUwww~www~www~www~www~www~www~UUUUwfwnwvw~wfw~wvw~www~wfw~wgw~UUUUuwwwuwwwuwwwwWwwwWwwwWuwWUwwUUUUwwwwwwwwwwwwwwwwWwwwwwwwwwwwUUUUwwwdwwwdwwwdwwwdwwwdwwwdwwwdUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwUUUVwwwvwwwvwwwvwwwvwwwvwwwvwwwvGtwwGtwwGtwwGtwwGtwwGtwwGtwwGtwwwwwtwwwtwwwtwwwtwwwtwwwtwwwtwwwtww�www�www�www�www�www�www�www�w�www�www�www�www�www�www�www�wwwwwwdwwwdwwwdwwwdwwwdwwwdwwwdwwwdwwwvwwwvwwwvwwwvwwwvwwwvwwwvwwwvGtUUGTffGTffEdffEdffFdffFdffFdffUUUUfffffffffffffffffffffffff���UUUUffffffffffffffffffffffff����UU�Uff�eff�Vff�Vff�fff�fff�fʦ�f�UUU�fff�fff�fff�fff�fff�fff�fffUUUUffffffffffffffffffffffffffffwwwdwwwdd333d333d333d333d333dwwwwwwww33333333333333333333wwwvwwwv33363336333633363336FdffFdffAC333C333C333C333C333��������33333333333333333333�f�f�fFf�33�333�333�333�333�3�fff�fff33333333333333333333ffffffff33333333333333333333333d333d333d333d333d3333����wwww333333333333333333333333����wwww333633363336333633363333����wwwwC333C333C333C333C3333333����wwww33�333�333�333�333�33333����wwww�����<��5UUU5UUSU553SS2#33"532 5�����<��5UUU5UUUU555SSSS33333��������UUUUUUUU5555SSSS3333��������UUU�UU_�55=�SS]�33;������l���eUUUUUUSU552SS2#S3"3S2 0�����<��5UUU5UUSU552SS2#33"332 0����ȩ��S�UUU��US:�U59��38��009������<��UUUUUUUU5555SSSS33333������ÓUUX�UUS�SSX�553�338�003�����3���UUUU5UUUU555SSSS33333�����̚�Ue�5UX�U5Y�5X��S9��3����������UUUUUUUSU5523S2#"302 0�����<��5UUU5UUSU552SS2#33"302 0�����<��5UUV5UUUU555SSSU33353��������UUUUUUUUU5553SSS33330����l���eUUSUUU3SSS%U3"5S2#3S" "#  %                     200            "          "                         0;�  ��  �� ��  ۰  ۰  ��  ��                          #                         P"R                         "#                       "#  "                    0"                                                    �  9                     �#�� ��� ��� ��  �       02(�" �  � ��0(�������� �����   �                    "                         205            "         R 20R                                                                                    ��  ��  �� �� �  �  �  �   �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��  �S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �   3       �  �3 3�=������<��̼��� �3 33==ƙ�<ə�ƙ�3ƙ��ƙ���i� 3= ��3=�l�ә��<��l<��l<��l<���<    �   3=  �30 ��� ���=��������                        +   3     0  �<  3� 3� =� =� 0� 0������������������3�33033�0�3�0��;f��;��̽�������3��3��<���<�f���̳=�=�������3303<�<00�<30�3����������������=��=��3�3�=�3�0  �=  �3  �3� ��0 ̳0 �0 �0  0� =� =� 3�  3�  �<  0  33�0�3�0�3�0�3303�303�303�303303��<���0<��0<033<033003300330033030�30�<00�<0330333033303330333033�0��<���0�03303303=03=03��0 ̳0 ��0 �3� �3� �=  0  3�     �                           <�03=��3=�� 3��  �=  �        033003300330�330��303= ��33    330333033303330333<��333ݰ    0=�0<3���;�3 �=  3�             �                           wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  ""   "! " ""                                                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  " ! " ""  "!    " ""                                                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  ""   "! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��     �                                 � ����                               �                        ���� ��� ����                            ��  ��  ���                        "  "  "                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��     �                         ���  +"  "" ���������                   �                        ���� ��� ����                            ��  ��  ���        �   �                        �   ��  �   ��   �       �                                                                                                                                               �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                             �� ��������p��}`         �  ��  �  �  ��  �                   �                        ���� ��� ����                            ��  ��  ��� �"�!/"�  �                                                                                                                                                                                  	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                        �          �   � � �  ��� ��  �                    �                        ���� ��� ����          �   �   �   �  �  �  �  �                                                                                                                                                                                                                         	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                                   ��          ��                                ��                                      ��  ��  ���                                                                                                                                                                                                                   �� ̻ ��˛��  �� �˚̻���ۚ����I���䘼�^���^�٘�:�^�� ^�� D�( �) �) �) ��) ˹� ț�+��,��,����  �𫝝 ��� �ɍ ��ݨ��ډ�݊�� ��D@ �D�  J�� ݩ� ��� �ۻ �ک �ڹ�ɻ��̸���������� ����������            �   ��  ��  ��  ��  ��                                          �� ��� ��� ��  �                         �   �    � � �     �   �                   �  �� Ș ��  ��  �                �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                         �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �       /�      �                           �   �   �   �   �   �                      �   �                      �������  ���    �       �  �  �  �                                 ���                              �   ���                            �   �                                                                                                   "  " �" ��" ��- �ۼ w۽��ݹ����� ��� ��  ˼  ��  ˼  ��  H�  �D  J�  J�  �  �  �  �  
�  �  �  �  ,�  " "" �" �"�   ˰  ��  wp ��ډ�v���r�̸��˰��� ��  ��  ��  ��  ̸  ��  ��  DC  C4@ T4@ T40 T30 T30 S;� H�  ��  ��  ��  ""  "  �""� "�/��        �   �   �      �  �   �   �   �   �              �   �   �   �             ���� �                        " "" """ �"  �   �   �                              � ��                  �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                                 � �� �������ۛ˽���� �ͼ ��+ �""�B.�R#Z�C U�D �T Z� �; � �� ��� ��  ��� ˽� �wp ��� �vp �w� ��� ˙� ̻� �۰ �ِ ��� Ш� �� >�" 3��.30" ��  �   �                �"/ "" ""  ��  ��                       �  �  ��  �   �       �   �   ��  �"" �""  ""   "                 �   ��   �                            � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                     �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                            �  �˰ ��� �wp ���                                                                                                                                                                 "  " �" ��" ��- �ۼ w۽��ݹ����� ��� ��  ˼  ��  ˼  ��  H�  �D  J�  J�  �  �  �  �  
�  �  �  �  ,�  " "" �" �"�   ˰  ��  wp ��ډ�v���r�̸��˰��� ��  ��  ��  ��  ̸  ��  ��  DC  C4@ T4@ T40 T30 T30 S;� H�  ��  ��  ��  ""  "  �""� "�/��        �   �   �      �  �   �   �   �   �              �   �   �   �             ���� �                        " "" """ �"  �   �   �                              � ��                  �  �˰ ��� �wp ���                                                                                                                                                                                  �� ̻ ��˛��  �� �˚̻���ۚ����I���䘼�^���^�٘�:�^�� ^�� D�( �) �) �) ��) ˹� ț�+��,��,����  �𫝝 ��� �ɍ ��ݨ��ډ�݊�� ��D@ �D�  J�� ݩ� ��� �ۻ �ک �ڹ�ɻ��̸���������� ����������            �   ��  ��  ��  ��  ��                                          �� ��� ��� ��  �                         �   �                           �   �                    �          �         �   �  �  �   �         �                                                                                                                                                                                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@       

 
� ��	�
�9 
Ð �� ��0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDDDN��DDN��DDN��DDDDDNDDDNDDDDDNvSV~DGefS5v~D�EfSs�~D3�fUS~NC3g�U3V�C3~S35ns31Wc3Sqe5gDvS3Uw�DD��ww���w����N���������ffEUUUA3333S3333333333333333333333333333333333333333333DDDDVfwwN��DvffUwvffwwvf�wwvwwwwffffUUUU333333333333333333333333333333333333333333333333DDDD����DDDDS5UUS3fUSffUSwvfUfffeUUUU333333333333333333333333333333333333333333333333DDDDwwvfDDDDffeSUffe5ffUfSVU3S3333333333333333333333333333333333333333333333333DDDDfUU3DDNN1U  SUPeSUfeSgve1UffU3UUf5V31533133333333313331333333333333333333333333DDDD35UDD��        P   UP  5f  fn` ge� ~G>`g�s�V~G>5g�qV~G5g�V~5n13W163U3533DDNvgwDD�NDN      �� 
��        
������� ��  �� 
�������                        �������         �����
�� 	�   ���������                          �  	�� 
�� ��� ����� ��  
�  	�   �   �                                                    �   �   �                       DD~DDDD�DDDNfnDDEV�D5TdDUdD5dDUF�DenDDDDDDDDDFNDDrDDvP530   �Nwg���eN��e��Nv�N�vGN~NFd�tFd~�F6G�v6TDc%ef#%RR521520       w�DNV~��1fwfSUQfS�eUVN���tDDD����DDDDffff23S%S!" 2# 3 0   #����uf~NQgt�3n�DV~NDf�dN�GdDD~dN~�dNNcfDeVVD%5bt25gSU % 0 3                               ~  nDDDDD DD ��! %          �w D~ w~ D~�w~�~��D�DDDDDDDDDDDDDDDDDDDDDDDDDDD0S"     ~DN~�DN�DDNDDDNDDDDDDDDDDDDDDDDDDDDDDDDDDDDNDDD�DD�b#R23       DDN�DD�DDNDDD�DNDDD�DD�eNDDUDD�d�D��fdNNbdND&D�RtDSVt %"   DDG�DDDNDDDD�f�DeTnDCUVDQ5VDQFDTUnD�V�DDDDD�DDDD�DGDDGe3%  N��vN�Nv��NvNN��N��GDt��DfNgDfG�Dfd~GeeDF!VVe%%Ue"P3"S%3"Q    w~�DUg��Sgve1UUfe1�fUUD���gDDD����DDDDffff!2RR223% # 0   ��~��Vg�ewN6��5g��fnFD��vDDG�Dw�fDD�SdfRb4RU&cRV"3Q                               0  � dD �D �D  n�           w  �G  ww G� ww����~DDD�DDDDDDDDDDDDDDDDDDD�DDDR%       w�D��DD��DD�DDD�DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDNDDN�52RR        �DD�DDNDDD�DDNDDDDDNDDNFD�DEDDNFNdNNFfD��&D�b5dNR"gDPP5g  0   DDG�DDDNDDDD�f�DeEnDSUVDA5FDQVDUEnD�V�DDDDD�DDDD�DGDDGcRR2   N��vN�Nv��NvNN��N��GDt��DfNgDfG�Dfd~GeeDFRVVe5bRPR%       w~�DUg��Sgve1UUfe1�fUUD���gDDD����DDDDffff2QRU2! %0     ��~��Vg�ewN6��5g��fnFD��vDDG�Dw�fDD�VdfUed2VgR""#Q%"                             0     �  dD0�D  �D  n�            w  �G  ww G� ww����~DDD�DDDDDDDDDDDDDDDDDDD�DDD"       w�D��DD��DD�DDD�DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDNDDN�"%Q        �DD�DDNDDD�DDNDDDDDNDDNFD�DEDDNFNdNNFfD��VD�aedNRQgD0R%g RP   �DDNDDDDDDDDD�f�NeEnFSUVEA5FFQVNUEn��V��DDDN�DDDD�DgDDGSS00    ���wNDfDNgQDD�eDFN�DDdNDD�DDeDD%DG&UDFb0DuV GbU2fP5UR    ~@  vt` Vv� U� g~� ��@ DN` 00    5S  "5  20  R5           N�DD�DDDDDDDDNfnD�EV�e5TDUU�d5��UFNNenNDDDD�DDtDNDStDD%RS    �N�wD�FaDD�uDDNv�Dd�dDFDdDFndDF �DFQDDveDDfQDGUeDv%%vaP%    w�  WgF gn QU^ fw� ��D DD� "   P   RR1 0 %  5R         N�DD�DDDDDDDDNfnD�UF�d5UDUU�e4��EVNNenNDDDD�DDtDNDStDDSSU    �N�wD�FaDD�uDDNv�Dd�dDFDdDFndDFQ�DFVDDveDDfRDGUeDvRRvbRR     w�  WgF gn QU^ fw� ��D DD�     ! QQ  %P Q U% PP                     �� ~DD 䪤 �IG j�� �i��� M��K��kK���K�w�G��{Ggw�                        	�  ��  �� �  ~� � ��� ���wDD�DDD�~DD              ~� �D J� �� �� ֚ m�`K���F���K���K�w�G��{Ggw�                @   @   p   �		  	�� 	�~ ��� ��������wDD�DDD�~DD              �  ~D  �J  �  j�  �n ��@���F���K���K�w�G��{Ggw�            �   D   �   �   �   � D  �~  �z�ݙw�ݖ��wDD�DDD�~DD              �  ~D  �D  ��  n�  �n ��@���F���K���K�w�G��{Ggw�            �   D   �   I   �   � D  G~  I|�j�|�5���wDD�DDD�~DD    `   �   `  s�  G>` �uu �GVP�Ne`~��pg�FpV�Fpg�Fp~Dg`DD~ �D@                                                                                          0                               1                            "S%3"Q                         # 0    0                  "3Q                            UU  Q  SV  UU  ff DD ��   �fNvQVN�ceD�eUdNvfdN�DDD��DD�D~�NNvffD�UU�E5tEfUnEUfvff  D   D Nu1gfffg�DDn�~�d�fgfGcVDGe6NvR"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��                                 � � �� � � � � ����l(�(a(�����������������                	 
   ��� � � � � �����y(�(�����������������   ������� ������� �� ������������   � � � � � � � �����((�l(=����������������   ��	�
��������    ��������������������   ��� � � � � �����((�(( ����������������        ����     ! " # # $! % &  ����  ' (����� � � �����(-(5(Xx���������������� ) * + , - .  �ܤ�  / 0 � 1 2�� 3 4  �֤� / 5 6+*) � � � ��� � �����(�xww����������������     7 8 9 : : : : : ; < = = = = = = > ?::::: @ A B     � � � � ��� �����ww�(���������������� C CC 7 8 DD  E F G H         DD  E F G H A B CCC �� � � ��� �� ����(+((�����������������    7 8                       A B   �� � � ��� � ����(W(�m(`����������������   Q 7 8                       A B(Q   � � � � ��� ���	B�(a((M���������������� V W X 7 8                       A B(XWV � � � ��� � ���	C�(-(� 
(����������������� V W \ 7 8                       A B(\WV� ���� � � ��	E	D�(( (-(����������������� V W ] ^ _ ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` a b(]WV��� � � � � ��	F ��(X((6(5���������������� V W c d e f g h i j V W  k h i d e f l V W(j m(h(g(f(e(dcWV � � � � � � � ��	G ��l((�x���������������� V W n o p q ] r s t V Wn ] r u o p q v V W(t(s(r(](q(p(onWV���������H������yxww���������������� V W w f g h i d e f V W x i d e f k h y V W(f(e(d(i(h(g(f(QWV � ��O�N�M�L�K�J�I������w(+�(���������������� V W z { ] r u o p q V W | u o p q ] r u V W(q(p(o(u(r(](q }WV�A�A�V�U�T�S�R�Q���P(�((5(U(,���������������� V W ~  � � � � � � � � � � � � � � � ���(��(��(�(�((~WV�]�]�\�[�Z�Y�X���P(N(,(U((=((+���������������� � � � � � � �  �   �  � �� �� �  � �� � � � ���U�U�b�a�`�_���P(U(V(=((( ((5���������������� �     � � � � � � � � � � � �����������    ��i�h�g�f�e���P)d((( ((,(U((=���������������� � � � � � � � � � � � � � � � � ����������� � � � ���u�t�s�r�p�p�-(,(N(,(U((=((( ���������������� � � � � � � � � � � � � � � � � � �� � � � � � ��� � � � ��!x!y!z!{!|!}!y!~ � � � � � � � ����������������� � � � ��� � � � � ��� � � �� � ���� � � � � ���� � �!!�!�!�!�!�!�!� � � � � � � � ����������������� � � � � � � � � � � � � � � � ��� � � � � � � � � � �� � � ��� � � � � � �����(W(�m(`���������������� � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �	
	
	
	
	@���(a((M���������������� � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � � �� � � � � � �����(-(� 
(����������������� � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �� � �� � � � �� ���(( (-(����������������� � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq"(c�<"�DT
t"��*�D2X=2	P]2	
l}~D �" � � " � � " � � "M �  *NO �*P �  )�` � c�G*"� �* "�
"� �*� �@"�_@ "�q0�W0
�f@ "G x@  *G�X  *KxX  *HxH  *PxX  *HxH "*PxX  *HxH $*PxX  *Hx �&J� z � 'J� z �(B� � � )B� G*"�.G +"�@7,"�&7-*�53."�3 /"�#0� #1
� � 2*Oz � 3*BzH  *PRH  *PRH  *PRX  *KRX  *KRX  *KR � 
�	 z;"H �  *Hx �  *Hx �>b` � � b^ �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� � � �m�n�|�}�c�d�v�w��� � � � � ������������������������������������������������� � � ������������������ � � � � ��������������������������������������������������!��?�K�X�H�K�K�Q��a��b� � � ������������������������������������������������� � � � � � � � � � � � � � � � � ������������������������������������������������� � � � � � � � � � � � � � � � � ������������������������������������������������� � � � � � � � � � � � � � � � � �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��$������������������2�0�.� �� �������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������/�.�7� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������/�^�O�Z��1�G�S�K�������������������������1�G�S�K��<�Z�G�Z�Y�����������������������9�R�G�_�K�X��<�Z�G�Z�Y��������������������<�I�U�X�O�T�M��<�[�S�S�G�X�_�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������/�+��2�U�I�Q�K�_��8�O�M�N�Z��������0�����������=�U�X�U�T�Z�U� � � � � � � � � � � � � � ��� ����������9�N�O�R�G�J�K�R�V�N�O�G� � � � � � � � � ��� ������������������������������������ 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                       	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                