GST@�                                                           �[�                                                      ��I                      ���2�����	 ʴ����������H�������        �g     #    ����                                d8<n    �  ?     �b����  �
fD�
�L���"����D"��   " `  J  jF��     �j  
 ���
��
��    "�j��" " ��
  y                                                                               ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������=o  0  4g  1                      �                         �  �  �  �                  n�  	          8 �����������������������������������������������������������������������������                                D              @  &   �   �                                                                                 '       )n)n1n  	n�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E 3 �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������     ��aA�S� o� �� o��hi o�p@.A�4m ��J�TsZ3��T0 k� ��^��^	E1 4#Q&�1D"3Q. ��    � <����xA�� �F  X �h�  ��@��xA]F�A]�XZ3� T0 k� ��F��F	E1 4#Q&�1D"3Q. ��/ 	   � �d��xA�� �F  X �h�  ��@��xA]F�A]�XZ3� T0 k� ��F��F	E1 4#Q&�1D"3Q  /�/ 	   � �f��xA�� �F  X �h�  ��@��xA]F�A]�XZ3� T0 k� ��F��F	E1 4#Q&�1D"3Q  ��/ 	   � �h��xA����F  X �h�  ��@��xA]F�A]�XZ3� T0 k� ��F��F	E1 4#Q&�1D"3Q  ��/    � �j��xA����F  X �h��@��xA�F�A��XZ3� T0 k� ��F��F	E1 4#Q&�1D"3Q  ��/    � �l��xA����F  X �h��@��xA�F�A��XZ3� T0 k� ��F��F	E1 4#Q&�1D"3Q  ��/    � �n��xA����F  X �h��@��xA�F�A��XZ3� T0 k� ��F��F	E1 4#Q&�1D"3Q  ��/    � �p��xA����F  X �h��@��wA�F�A��XZ3� T0 k� ��F��F	E1 4#Q&�1D"3Q  ��/    � �qL�xDܤ��F  X lh��CL�wA�F��A��XZ3� T0 k� ��F��F	E1 4#Q&�1D"3Q  ��/    � �rL�xDܤ��FL X lh�\�CL�wA�F��A��XZ3� T0 k� ��F��F	E1 4#Q&�1D"3Q  ��/    � �sL�wDܤ��FL X lh�\�CL�vA�F��A��XZ3� T0 k� ��F� F	E1 4#Q&�1D"3Q  ��/    � �tL�wDܨ��FL X lh�\�CL�vA�F��A��XZ3� T0 k� � F�F	E1 4#Q&�1D"3Q  ��/    � �uL�wDܨ��FL X lh�\�CL�uA�F��A��XZ3� T0 k� �F�F	E1 4#Q&�1D"3Q  ��/    � �vܤwDܨ��FL X h�\�CL�uA�F��A��XZ3� T0 k� �F�F	E1 4#Q&�1D"3Q  ��/    � �xܤwDܬ��F�X h���CL�tP�F��BM�XZ3� T0 k� �F�F	E1 4#Q&�1D"3Q  ��/    � �yܤvDܬ��F�W h���CL�sP�F��BM�XZ3� T0 k� �F�F	E1 4#Q&�1D"3Q  ��/    � �zܨvDܰ��F�W h�	��C\�sP�F��BM�XZ3� T0 k� �F�F	E1 4#Q&�1D"3Q  ��/    � �{ܨvD���F�W h�	��C\�rP�F��BM�XZ3� T0 k� �F� F	E1 4#Q&�1D"3Q  ��/    � �|ܬuD���F�W�h�	��C\�qP�F��BM�XZ3� T0 k� � F�$F	E1 4#Q&�1D"3Q  ��/    � �}ܬuD���F�V�h�
��C\�pP�F��@m�XZ3� T0 k� �$F�(F	E1 4#Q&�1D"3Q  ��/    � �~ܰtD���F�U�l�
��C\�nP�$F=�@m�XZ3� T0 k� �,F�0F	E1 4#Q&�1D"3Q  ��/    � ��tD���F�U�l���C\�mP�(F=�@m�XZ3� T0 k� �0F�4F	E1 4#Q&�1D"3Q  ��/    � ��tD���F�T�l���C\�lP�,F=�@m�XZ3� T0 k� �,F�0F	E1 4#Q&�1D"3Q  $�"    � ��sD���F�T�p���C\�kP�,F=�@��XZ3� T0 k� -$G�(G	E1 4#Q&�1D"3Q  ��"    � ��rD����F�S�p���C\�iP�0F=�@��XZ3� T0 k� -$G�(G	E1 4#Q&�1D"3Q  ��"    � ��qD����F�R�t���C\�gP�8F-�@��XZ3� T0 k� -(G�,G	E1 4#Q&�1D"3Q  ��"    � ��qD�� ��FR�t���I\�eP�8F-�@��XZ3� T0 k� -(G�,G	E1 4#Q&�1D"3Q  ��"    � ��pD�� ��FQ�t���I\�dP�<F-�@m�XZ3� T0 k� �(G�,G	E1 4#Q&�1D"3Q  ��"    � ��pD��!��F P�x���I\�cP�@F-�@m�XZ3� T0 k� �(G�,G	E1 4#Q&�1D"3Q  ��"    � ���oD��"��F(O�x���I\�aE�DF-�!@m�XZ3� T0 k� �0G�4G	E1 4#Q&�1D"3Q  ��"    � ����nD��# F�(N�x���I\�`E�HF�"@m�XZ3� T0 k� �(E�,E	E1 4#Q&�1D"3Q  ��"    � ����nD��$F�,N�x���Il�_E�LG�#B��WZ3� T0 k� �$C�(C	E1 4#Q&�1D"3Q  ��"    � ����mD��%F�4M�|���	Il�]E�PG�%B��WZ3� T0 k� �(B�,B	E1 4#Q&�1D"3Q  ��"    � ����mD��%F�8L�|���Il�\FTH�%B��VZ3� T0 k� �(A�,A	E1 4#Q&�1D"3Q  ��"    � ����mD��%F�<L�|���Il�[FXH�&B��TZ3� T0 k� �(@�,@	E1 4#Q&�1D"3Q  ��"    � ����mE�&F�@K�|���I\�[FXH�'B�SZ3� T0 k� �,@�0@	E1 4#Q&�1D"3Q  ��"    � ����mE�&F�HJ�|���I\�ZF\I�(B�RZ3� T0 k� �0@�4@	E1 4#Q&�1D"3Q  ��"    � ����lE�'M G�PJ�|���I\�XFdJ��*B�OZ3� T0 k� �<@�@@	E1 4#Q&�1D"3Q  �"    � ��L�lE�'M$G�TI�|��� I\�WBMhK��+B�NZ3� T0 k� �D@�H@	E1 4#Q&�1D"3Q  �"    � ��L�lE�'M(G�XIL|���E,�WBMlK��+B��LZ3� T0 k� �L@�P@	E1 4#Q&�1D"3Q  ��"   � ��L�lE�(M,G�\HL|���E,�VBMpL��,B��KZ3� T0 k� �P@�T@	E1 4#Q&�1D"3Q  ��"    � ��L�lE�(M0G�\HL|���E,�UBMtL��-B��JZ3� T0 k� �T@�X@	E1 4#Q&�1D"3Q  ��"    � ��L�lE�)M4G�`GL|���E,�TBMxM��.B��IZ3� T0 k� �X@�\@	E1 4#Q&�1D"3Q  ��"    � �� �lE�*M4G�dGL|���E,�SBM|MM�.B��HZ3� T0 k� �\@�`@	E1 4#Q&�1D"3Q  ��"    � �� �lE�*M8G�hF |���E,�SBM�NM�/B��FZ3� T0 k� �`A�dA	E1 4#Q&�1D"3Q  ��"    � �� �lD��+M<G�lF |���@l�RBM�NM�0B��EZ3� T0 k� �dA�hA	E1 4#Q&�1D"3Q  ��"    � �� �lD��+M@G�pF |���@l�QBM�OM�0B��DZ3� T0 k� �hA�lA	E1 4#Q&�1D"3Q  ��"    � �� �lD��,MDG�tE |���@l�QBM�OM�1B��CZ3� T0 k� �x@�|@	E1 4#Q&�1D"3Q �"    � ����lD��-]HG�xE |���@l�PBM�OM�2B��BZ3� T0 k� ��?��?	E1 4#Q&�1D"3Q ��/    � ����kD��.]LG�|D�|���@l�OBM�PM�2B��BZ3� T0 k� ��?��?	E1 4#Q&�1D"3Q ��/    � ����kD��/]PG�|D�|���@l�NBM�PM�2B��BZ3� T0 k� ��>��>	E1 4#Q&�1D"3Q ��/    � ����kD��/]PG��D�|���@l�NBM�QM�2B��BZ3� T0 k� ��>��>	E1 4#Q&�1D"3Q ��/    � ����kD��0]TG��C�|���@l�MBM�QM�2B��BZ3� T0 k� ��=��=	E1 4#Q&�1D"3Q	 ��/    � ����kD��1mXG��C�����@l�LBM�RN 2B��BZ3� T0 k� ��=��=	E1 4#Q&�1D"3Q
 ��/    � ����kD��2m\G��C�����@l�LBM�RN 2B��BZ3� T0 k� ��<��<	E1 4#Q&�1D"3Q ��/    � ����kD��3m\G��B�����@l�KBM�RN2B��BZ3� T0 k� ��;��;	E1 4#Q&�1D"3Q �/    � ����kD� 4m`G��B�����@l�KBM�SN2Q]�BZ3� T0 k� ��;��;	E1 4#Q&�1D"3Q ��/    � ����kD�5mdG��B�����@l�JBM�SN2Q^ BZ3� T0 k� ��:��:	E1 4#Q&�1D"3Q ��/    � ����kD�6mhG��A�����@l�IBM�TN2Q^BZ3� T0 k� ��:��:	E1 4#Q&�1D"3Q ��/    � ����kD�8mhG��A����@l�IBM�TN2Q^AZ3� T0 k� ��:��:	E1 4#Q&�1D"3Q ��/    � ����kD�9mlG��A����@l�IBM�TN2Q^AZ3� T0 k� ��9��9	E1 4#Q&�1D"3Q ��/    � ����kD�9mpG��@����@l�IBM�UN1Q^AZ3� T0 k� ��9��9	E1 4#Q&�1D"3Q ��/    � ����kF:mpG��@����@l�IBM�U�1Q^AZ3� T0 k� ��8��8	E1 4#Q&�1D"3Q ��/    � ����kF :mtG��@����@l�IBM�V�1Q^AZ3� T0 k� ��8��8	E1 4#Q&�1D"3Q ��/    � ����kF$;mxG��?����@l�IBM�V�1QnAZ3� T0 k� ��7��7	E1 4#Q&�1D"3Q ��/    � ����jF,<mxG��?����@l�JBM�V�1QnAZ3� T0 k� ��7��7	E1 4#Q&�1D"3Q ��/    � ��� jF0<m|H��?����@l�JBM�W�1QnAZ3� T0 k� ��6��6	E1 4#Q&�1D"3Q ��/    � ���jF4=m�H��>����@l�JBM�W~0QnAZ3� T0 k� ��6��6	E1 4#Q&�1D"3Q ��/    � ���jF<>m�H��>����@l�JBM�W~0Qn AZ3� T0 k� ��5��5	E1 4#Q&�1D"3Q
 ��/    � ���jL}@?m�H��>����@l�JBM�X~0Qn$AZ3� T0 k� ��5��5	E1 4#Q&�1D"3Q
 ��/    � ���jL}H?m�H��>����@l�JBM�X~ /Qn$AZ3� T0 k� ��5��5	E1 4#Q&�1D"3Q	 ��/    � ���jL}L@m�H��=����@l�JBM�X~ /Q~(AZ3� T0 k� �4��4	E1 4#Q&�1D"3Q	 ��/    � ���$jL}L@m�H��=����@l�JBM�Y~$.Q~,AZ3� T0 k� �4��4	E1 4#Q&�1D"3Q	 ��/    � ���(jL}P@m�H��=����@l�JBM�Yn$-Q~,AZ3� T0 k� �3��3	E1 4#Q&�1D"3Q ��/    � ���0jL}TA �H��=����@l�JBM�Yn(-Q~0AZ3� T0 k� �3��3	E1 4#Q&�1D"3Q ��/    � ���8jL}XA �I��<����@l�JBM�Zn(,Q~0AZ3� T0 k� �2��2	E1 4#Q&�1D"3Q ��/    � ���<jL}\B �I��<����@l�JBM�Zn(,Q~4AZ3� T0 k� �2��2	E1 4#Q&�1D"3Q ��/    � ���DjL}`B �I��<����@l�JBM�Zn,+Q~8AZ3� T0 k� �1��1	E1 4#Q&�1D"3Q ��/    � ���LjL}`C �I��<����@l�JBM�Zn,*Q~8AZ3� T0 k� �1��1	E1 4#Q&�1D"3Q ��/    � ���PjL}dC �I��;� ���@l�JBM�[^,)Q~<AZ3� T0 k� �1��1	E1 4#Q&�1D"3Q ��/    � ���XjL}hD �J��;�!���@l�JBM�[^,)Q~<AZ3� T0 k� �0��0	E1 4#Q&�1D"3Q ��)    � ���`jL}lD �J��;,�"���@l�JBM�[^,(Q~@AZ3� T0 k� ��/��/	E1 4#Q&�1D"3Q ��)    � ���hjL}lD �J��;,�#���@l�KBM�\^,'Q~@AZ3� T0 k� ��/��/	E1 4#Q&�1D"3Q ��)    � ���pjL�pE �J��:,�$���@l�KBM�\^,'Q~DAZ3� T0 k� ��.� .	E1 4#Q&�1D"3Q ��)   � ���xjL�tE �J��:,�%���@l�KBM�\^,&Q~DAZ3� T0 k� � -�-	E1 4#Q&�1D"3Q ��)    � ���jL�xF �J��:,�&���@l�KBM�\N,%Q~HAZ3� T0 k� �/�/	E1 4#Q&�1D"3Q  ��)    � ���iL�xF �K��:,�'���@l�KBM�]N,%Q~HAZ3� T0 k� �0�0	E1 4#Q&�1D"3Q  ��)    � ���iL�|F �K��:,�)���@l�KBM�]N,$Q~LAZ3� T0 k� �1�1	E1 4#Q&�1D"3Q  ,�)    � ���iL��G �K��9,�)���@l�KBM�]N($Q~LAZ3� T0 k� �1�1	E1 4#Q&�1D"3Q  ��)    � ���iL��G �K��:,�)���@l�KBM�]N($Q~PAZ3� T0 k� �2�2	E1 4#Q&�1D"3Q  ��)    � ����iL��G �K��:,�*���@l�KBM�^N(#Q~PAZ3� T0 k� �2�2	E1 4#Q&�1D"3Q ��)    � ����hL��H �K��:,�+���@l�KBM�^N(#Q~TAZ3� T0 k� �2�2	E1 4#Q&�1D"3Q ��)    � ����hL��H �L��;��+���@l�KBM�^$#Q~TAZ3� T0 k� ��2��2	E1 4#Q&�1D"3Q ��)   � ����hL��H �L��;� ,���@l�KBM�^$"Q~XAZ3� T0 k� ��2��2	E1 4#Q&�1D"3Q ��)    � ����hL��I �L��;�-���@l�KBM�^ "Q~XAZ3� T0 k� ��1��1	E1 4#Q&�1D"3Q ��)    � ����hL��I �L��;�.���@l�KBN ^ "Q~\AZ3� T0 k� ��1��1	E1 4#Q&�1D"3Q ��)    � ����hL��I �L��;�/���@l�KBN^"Q~\AZ3� T0 k� ��1��1	E1 4#Q&�1D"3Q ��)    � ����hL��J �L��;�/���@l�LBN]"Q~`AZ3� T0 k� ��1��1	E1 4#Q&�1D"3Q ��)    � ����hL��J �M��;�0���@l�LBN]"Q~`AZ3� T0 k� ��1��1	E1 4#Q&�1D"3Q ��)    � ����hL��J �M��;�$1���@l�LBN]"Q~`AZ3� T0 k� ��1��1	E1 4#Q&�1D"3Q ��)    � ����hL��K �M��<�(2���@l�LBN]"Q~dAZ3� T0 k� ��1��1	E1 4#Q&�1D"3Q ��)    � ����hL��K �M��<�03���@l�LBN\"Q~dAZ3� T0 k� �1��1	E1 4#Q&�1D"3Q ��)   � ����hL��K �M��<�44���@l�MBN\"Q~hAZ3� T0 k� �1��1	E1 4#Q&�1D"3Q ��)    � ����hL��L �M��<�<5���@l�MBN\"Q~hAZ3� T0 k� �1��1	E1 4#Q&�1D"3Q ��)    � ����hL��L �M��<@6���@l�MBN [."Q~hAZ3� T0 k� �1��1	E1 4#Q&�1D"3Q ��)    � ����hL��L �N��<H7���@l�MBN$[.#Q~lAZ3� T0 k� �2��2	E1 4#Q&�1D"3Q ��)    � ��}�hL��L �N��<P8���@l�MBN([.#Q~lAZ3� T0 k� ��2��2	E1 4#Q&�1D"3Q ��)    � ��}�hL��M �N��<T9���@l�MBN,Z. #Q~lAZ3� T0 k� ��2��2	E1 4#Q&�1D"3Q ��)    � ��~hL��M �N��=\:���@l�NBN0Z-�#Q~pAZ3� T0 k� ��2��2	E1 4#Q&�1D"3Q ��)    � ��~gL��M �N��=`;���@l�NBN4Z��$Q~pAZ3� T0 k� ��.��.	E1 4#Q&�1D"3Q ��)    � ��~gL��N �N� =h<���@l�NBN8Y��$Q~pAZ3� T0 k� ��+��+	E1 4#Q&�1D"3Q ��)    � ��	�gL��N �N�=p>���@l�NBN<Y��$Q~tAZ3� T0 k� ��(��(	E1 4#Q&�1D"3Q ��)    � ��	�gL��N  N�=t?���@l�NBN@Y��$Q~tAZ3� T0 k� ��&��&	E1 4#Q&�1D"3Q ��)    � ��	�gL��N  O�=|@���@l�NBNDX��$Q~tAZ3� T0 k� ��%��%	E1 4#Q&�1D"3Q ��)    � ��	�gL��O O�=�A���@l�OBNHX��%Q~xAZ3� T0 k� ͼ$��$	E1 4#Q&�1D"3Q ��)    � ��	� gL��O O�=�B���@l�OBNLW��%Q~x@Z3� T0 k� ͸#��#	E1 4#Q&�1D"3Q ��)    � ��^$fL��O O�>�B���@l�OBNPW��%Q~x@Z3� T0 k� ����	E1 4#Q&�1D"3Q  ��)    � ��^(fL��P O�>�B���@l�OBNTW��%Q~|@Z3� T0 k� ����	E1 4#Q&�1D"3Q  ��)    � ��^(fL��Q O�>�C���@l�OBNXV��%Q~|@Z3� T0 k� ����	E1 4#Q&�1D"3Q  ��)    � ��^,fL��R O�$>�D���@l�OBNXV��%Q~|@Z3� T0 k� ����	E1 4#Q&�1D"3Q  .�)    � ��^0fL��R O�(>�E���@l�OBN\V��%Q~�@Z3� T0 k� ����	E1 4#Q&�1D"3Q  ��)    � ��^4fL��S O�,>��F���@l�PBN`V-�%Q~�@Z3� T0 k� ݜ��	E1 4#Q&�1D"3Q  ��)    � ��^8fL��S P�0>��F���@l�PBNdU-�&Q~�@Z3� T0 k� ݔ��	E1 4#Q&�1D"3Q  ��)    � ��^<fL��T�P�4>��G���@l�PBNhU-�&Q~�@Z3� T0 k� ݌��	E1 4#Q&�1D"3Q  ��)    � ��^<fL}�U�P�<>��H���@l�PBNhU-�&Q~�@Z3� T0 k� ݄��	E1 4#Q&�1D"3Q  ��)    � ��^@fL}�U�P�@>��H���@l�PBNlT-�&Q~�@Z3� T0 k� ݀��	E1 4#Q&�1D"3Q  ��)    � ��^DeL}�V�P�D?��H���@l�PBNpT=�&Q~�@Z3� T0 k� �|��	E1 4#Q&�1D"3Q  ��)    � ��nHeL}�W�P�L?��I���@l�PBNtT=�&Q~�@Z3� T0 k� �x�|	E1 4#Q&�1D"3Q  ��)    � ��nLeL}�X� P�P?��J���@l�PBNtT=�&Q~�@Z3� T0 k� �t�x	E1 4#Q&�1D"3Q  ��)    � ��nLeL}�Y� P�X?��J���@l�QBNxS=�&Q~�@Z3� T0 k� �l�p	E1 4#Q&�1D"3Q  ��)    � ��nPeF�Z�$P�\?��K���@l�QBN|S=�&Q~�@Z3� T0 k� �h�l	E1 4#Q&�1D"3Q  ��)    � ��nTeF�Z�$P�d?��L���@l�QBN|SM�&Q~�@Z3� T0 k� �d�h	E1 4#Q&�1D"3Q  ��)    � ��nXeF�[�(P�h?��L���@l�QBN�RM�&Q~�@Z3� T0 k� �`�d	E1 4#Q&�1D"3Q  ��)    � ��nXeF�\�(P�p?��M���@l�QBN�RM�&Q~�@Z3� T0 k� �\�`	E1 4#Q&�1D"3Q  ��)    � ��n\eF�]�,P�t@��M���@l�QBN�RM�&Q~�@Z3� T0 k� �X�\	E1 4#Q&�1D"3Q  ��)    � ��n`eE��^�,P�|@��N���@l�QBN�RM�&Q~�@Z3� T0 k� �T�X	E1 4#Q&�1D"3Q  ��)    � ��n`eE� ^�0P��@��O���@l�QBN�QM�&Q~�@Z3� T0 k� �T�X	E1 4#Q&�1D"3Q  ��)    � ��nddE�_�0P��@��O���@l�QBN�QM�&Q~�@Z3� T0 k� �P�T	E1 4#Q&�1D"3Q  ��)    � ��nhdE�`�4Q��A��P���@l�RBN�QM|&Q~�@Z3� T0 k� �L�P	E1 4#Q&�1D"3Q  ��)   � ��nhdE�a�4Q��A��P���@l�RBN�QMx&Q~�@Z3� T0 k� �H�L	E1 4#Q&�1D"3Q  ��)    � ��nldE�a�4Q��A��Q���@l�RBN�QMx&Q~�@Z3� T0 k� �D�H	E1 4#Q&�1D"3Q  ��)    � ��nldE�b�8Q��B��Q���@l�RBN�PMt'Q~�@Z3� T0 k� �@�D	E1 4#Q&�1D"3Q  ��)    � ��npdE� c�8Q��B��R���@l�RBN�PMp'Q~�@Z3� T0 k� �<�@	E1 4#Q&�1D"3Q  ��)    � ��ntdE�(c�<Q��C��S���@l�RBN�PMl'Q~�@Z3� T0 k� �8�<	E1 4#Q&�1D"3Q  ��)    � ��ntdE�,d�<Q��C��S���@l�RBN�PMh'Q~�@Z3� T0 k� �8�<	E1 4#Q&�1D"3Q  ��)    � ��nxdE�4e�<Q�D��T���@l�RBN�PMd'Q~�@Z3� T0 k� �4�8	E1 4#Q&�1D"3Q  ��)    � ��nxdE�8e�@Q�D��T���@l�RBN�P=d'Q~�@Z3� T0 k� �0�4	E1 4#Q&�1D"3Q  ��)    � ��n|dE�8e�@Q�E��U���@l�RBN�P=`'Q~�@Z3� T0 k� �,�0	E1 4#Q&�1D"3Q  ��)    � ��n�dE�<e�DQ�F� U���@l�RBN�P=\'Q~�@Z3� T0 k� �(�,	E1 4#Q&�1D"3Q  ��)    � ��n�dE�@e�DQ�F� U���@l�SBN�P=X'Q~�@Z3� T0 k� �(�,	E1 4#Q&�1D"3Q  ��)    � ��n�cE�Df�DQ��G�V���@l�SBN�P=X'Q~�@Z3� T0 k� �$�(	E1 4#Q&�1D"3Q  ��)    � ��n�cE�Hf HQ��G�W���@l�SBN�P-T'Q~�@Z3� T0 k� � �$	E1 4#Q&�1D"3Q  ��)    � ��n�cE�Lf HQ��G�W"��@l�SBN�P-P'Q~�@b�� T0 k� �� 	E1 4#Q&�1D"3Q  ��)   � ��n�cE�Pf HQ��H�W"��@l�SBN�P-L'Q~�@b�� T0 k� �� 	E1 4#Q&�1D"3Q  ��)    � ��n�cE�Pf LQ��H�X"��@l�SBN�P-L'Q~�@b�� T0 k� ��	E1 4#Q&�1D"3Q  ��)    � ��n�cE�Pf LQ��H�Y"��@l�SBN�O-H'Q~�@b�� T0 k� ��	E1 4#Q&�1D"3Q �)    � ��n�cE�Tf PQ� I�Y"��@l�SBN�OD'Q~�@b�� T0 k� ����	E1 4#Q&�1D"3Q ��/    � ��n�cE�Xf PQ�I�Z"��@l�SBN�OD'Q~�@b�� T0 k� ����	E1 4#Q&�1D"3Q ��/    � ��n�bE�\f PQ�I�["��@l�SBN�O@'Q~�?b�� T0 k� ����	E1 4#Q&�1D"3Q ��/    � ��n�bE�`f TQ�J�["��@l�SBN�O<'Q~�?b�� T0 k� ����	E1 4#Q&�1D"3Q ��/    � ��n�bE�de TQ�J�\"��@l�SBN�O<'Q~�?b�� T0 k� ����	E1 4#Q&�1D"3Q ��/    � ��n�bE�he TQ�J� \"��@l�TBN�O8'Q~�?b�� T0 k� ��
��
	E1 4#Q&�1D"3Q ��/    � ��n�bE�le XR�K�$]"��@l�TBN�O4'Q~�?b�� T0 k� �|��	E1 4#Q&�1D"3Q ��/    � ��n�bE�pd \R�K�$^���@l�TBN�O4'Q~�?Z3� T0 k� �h�l	E1 4#Q&�1D"3Q ��/    � ��n�bE�pd `R�K�(^���@l�TBN�O0'Q~�?Z3� T0 k� �T�X	E1 4#Q&�1D"3Q ��/    � ��n�bE�tc `R� K�,_���@l�TBN�O0'Q~�?Z3� T0 k� �@�D	E1 4#Q&�1D"3Q ��/    � ��n�bE�tc dS�$K�,_���@l�TBN�N,'Q~�?Z3� T0 k� �/��3�	E1 4#Q&�1D"3Q ��/    � ��n�aE�tc hR�$K�0`���@l�TBN�N('Q~�?Z3� T0 k� ����	E1 4#Q&�1D"3Q ��/    � ��^�aE�tc hR�(K�0a���@l�TBN�N((Q~�?Z3� T0 k� ����	E1 4#Q&�1D"3Q ��/    � ��^�aE�xc lR�,K�4a���@l�TBN�N$(Q~�?Z3� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aE�xc lR�0K�8b���@l�TBN�N$(Q~�?Z3� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aE�|c pR�0K�8b���@l�TBN�N (Q~�?Z3� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aE�|b tR�4K�<c���@l�TBN�N (Q��?Z3� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aC�|b tR�8L�<c���@l�TBN�N(Q��?Z3� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aC�|b xQ�8L�<c!���@l�TBN�N(Q��?bs� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aC�b xQ�8L�<c!���@l�UBN�N(Q��?bs� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aC�b |Q�<L�<d!���@l�UBN�N(Q��?bs� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aC�b |Q�<L�@d!���@l�UBN�N(Q��?bs� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aC�b �Q�@L�@e!���@l�UBN�N(Q��?bs� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aC�b �Q�@L�@e!���@l�UBN�M(Q��?bs� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aC�b �Q�DL�@e!���@l�UBN�M(Q��>bs� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�aC�b �Q�DL�@f!���@l�UBN�M(U.�>bs� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��~�aC��b �Q�HL�@f!���@l�UBN�M�(U.�>bs� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��~�`C��b �P�LL�@g!���@l�UBN�M�(U.�>bs� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��~�`C��b �P�LL�@g���@l�UBN�M�(U.�>Z3� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��~�`C��a �P�PL�@g���@l�UBN�M�(U.�>Z3� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��~�`C��a �P�PL�@h���@l�UBN�M�(U.�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��n�_C�|a �P�TL�@h���@l�UBN�M� (U.�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��n�_C�|a �P�TL�@h���@l�UBN�M� (U.�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��n�^C�|a �P�XL�@h���@l�UBN�M� (@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  .�/    � ��n�^C�|a �P�XL�@h���@l�UBN�M��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��n�]C�|` �P�\L �@h���@l�UBN�M��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��n�]Dx` �O�\L �<h���@l�VBN�M��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^�]Dx` �O�`L �<i���@l�VBN�L��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^�]Dt` �O�`L �<i���@l�VBN�L��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^�\Dt` �O�dL �<i���@l�VBN�L��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^�\Dp_ �O�dL �<i���@l�VBN�L��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^�\Dp_ �O�dM �<i���@l�VBN�K��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�\Dp_ �O�hM �<i���@l�VBN�K��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�[Dl^ �O�hM �<i���@l�VBN�K��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q ��/    � ��^�[Dl^ �O�lM �<i��#�@l�VBN�J��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����[Dl^ �O�lM<i��#�@l�VBN�J��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����[Lh] �O�lM<i��#�@l�VBN�J��(@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����ZLh] �O�pM<i��#�@l�VBN�J��)@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/   � ����ZLh] �O�pM8i��#�@l�VBN�I��)@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����ZLh] �N�pM8j��#�@l�VBN�I��)@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����ZLd] �N�pM�8j��#�@l�VBN�I��)@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����ZLd] �N�pM�4j��#�@l�VBN�I��)@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����ZL`] �N�pM�4j��#�@l�VBN�H��)@n�>Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����ZL`\ �N�pM�4j��#�@l�VBN�H��)@n�=Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����ZL\\ �N�pM�0j��#�@l�VBN�H��)@n�=Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����[L\\ �N�pM�0k��#�@l�VBN�H��)@n�=Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����[L\\ �N npM�,k��#�@l�VBN�G��)@n�=Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����[LX[ �N npM�(k��#�@l�VBN�G��)@n�=Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����[LX[ �N npM�(k��#�@l�VBN�G��)@n�=Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����[LX[ �N npM�$k��#�@l�VBN�G��)@n�<Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����\L.X[ �N npM� k��#�@l�WBN�F��)@n�<Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����\L.X[ �NNpM� k��#�@l�WBO F��)@n�<Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����\L.X[ �NNpM�j��#�@l�WBO F��)@n�<Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����\L.X[ �NNpM�j��#�@l�WBO F��)@n�<Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����]L.X[ �NNpM�j��#�@l�WBO F��)@n�<Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/   � ����]L.X[ �NNpM�j��#�@l�WBO E��)@n�;Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ����]L.X[ �N �pM�i��#�@l�WBOE��)@n�;Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/   � ����]L.X[ �N �pMi��#�@l�WBOE��)@n�;Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���^L.X\ �M �pMh��#�@l�WBOE��)@n�;Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/   � ���^L.X\ �M �pMh��#�@l�WBOE��)@n�;Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���^L.T\ �M �pMg��#�@l�WBOD��)@n�;Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���^L.T\ �M�pMg��#�@l�WBOD��)@n�;Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���^L.T\ �L�pM�f��#�@l�WBOD��)@n�:Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��ޜ_L.P\ �L�lM�f��#�@l�WBOD��)@n�:Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��ޘ_L.P\ �L�lM�e��#�@l�WBOD��)@n�:Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��ޔ_L.P] �L�lN�e��#�@l�WBOD��)@n�:Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��ޔ_L.L] �K�lN�d��#�@l�WBOC��)@n�:Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/   � ��ސ_L.H] �K�hN�d��#�@l�WBOC��)@n�:Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���_L.D] �K�hO�d��#�@l�WBOC��)@n�:Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���_L.@] �K�dO�d��#�@l�WBOC��)@n�:Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���_L.@] �K�dO�c��#�@l�WBOC��)@n�9Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���_L.@] �J�`O�c��#�@l�WBOC��)@n�9Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���_L.@] �J�`O� c��#�@l�WBOB��)@n�9Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��>�_L.@^ �J�`O� c��#�@l�WBOB��)@n�9Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��>�_L.@^ �J�\O� c��#�@l�WBOB��)@n�9Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��>�_L.@^ �J�\O��c��#�@l�WBOB��)@n�9Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��>�_L.@^ �I�XO��c��#�@l�WBOB��)@n�9Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��>�_L.<^ �I�XO��c��#�@l�WBOB��)@n�9Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^|_L.8^ �I�XO��c��#�@l�WBOA��)@n�9Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^|_L.8^ �I�TO��c��#�@l�WBOA��)@n�9Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^x_L.8^ �I�TO��c��#�@l�WBOA��)@n�8Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^x_L.8^ �I�TO��c��#�@l�WBOA��)@n�8Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^x_L.4_ �H�TO��c��#�@l�XBOA��)@n�8Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^x_L.0_ �H�TO��c��#�@l�XBOA��)@n�8Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��^t_L.0_ �H�TO��c��#�@l�XBOA��)@n�8Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���t_L.0_ �H�TO��b��#�@l�XBOA��)@n�8Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���t_L.0_��H�TO��b��#�@l�XBO@��)@n�8Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���t_L.,_��HTO��b��#�@l�XBO@��)@n�8Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���t_L.,_��HTO�b��#�@l�XBO@��)@n�8Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���p_L.,_��HPO�a��#�@l�XBO@��)@n�8Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��p_L.,_��HPO�a��#�@l�XBO@��)@n�7Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/   � ��p_L(_��HPO�a��#�@l�XBO@��)@n�7Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��p_L(_��H�PP�`��#�@l�XBO@��)@n�7Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��p_L(_��H�PP��`��#�@l�XBO@��)@n�7Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��l_L$_��H�PP��`��#�@l�XBO@��)@n�7Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��l_L$_��H�LP��`��#�@l�XBO?��)@n�7Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��h_L$_��H�LP��`��#�@l�XBO?��)@n�7Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��h_C�$_��G�LP��`��#�@l�XBO?��)@n�7Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��h_C�$_��G�HP��`��#�@l�XBO?��)@n�7Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��h_C�$^��G�HP��`��#�@l�XBO?��)@n�6Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��d`C�$^��G�DP��`��#�@l�XBO?��)@n�6Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��d`C�$^��G�DP��_��#�@l�XBO?��)@n�6Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��.d`C�$^��G�DP��_��#�@l�XBO?��)@n�6Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ��.d`C�$^��G�DP��_��#�@l�XBO?��)@n�6Z3� T0 k� ������	E1 4#Q&�1D"3Q  ��/    � ���PE˙	.��M+�s�|�=�E}��O��B��GZ3��T0 k� � �	E1 4#Q&�1D"3Q  ��U    � 
�d�XEә	.��M'�s�|�=�E}��O��B��GZ3��T0 k� ��	E1 4#Q&�1D"3Q  ��U    � 
�e�`Eט	.��M'��w�|�=�E}��O��B� GZ3��T0 k� ��	E1 4#Q&�1D"3Q  ��U    � 
�f�pE�	.��M��{�|�=�E~�O(��B�GZ3��T0 k� ��	E1 4#Q&�1D"3Q  ��U    � 
�g�xE�	��M��{�} M�E��O0��J@GZ3��T0 k� ��	E1 4#Q&�1D"3Q  ��U    � 
�h�� E�	��M���}M�E��O4 �#�J@ GZ3��T0 k� ��	E1 4#Q&�1D"3Q  ��U    � 
�i��"E���	��=���}M�E��O<!�'�J@(GZ3��T0 k� �� 	E1 4#Q&�1D"3Q  ��U    � 
�j��$E��	��=����}
M�E��OL#�3�J@4HZ3��T0 k� �$	�(		E1 4#Q&�1D"3Q  ��U    � 
�k��&E��	.��=����}
M�E��OT$�;�E0<HZ3��T0 k� �(
�,
	E1 4#Q&�1D"3Q  ��U   � 
�l��'E��	.��=����}M�E�#�OX%�C�E0DHZ3��T0 k� �,
�0
	E1 4#Q&�1D"3Q  ��U    � 
�m��(E�#�	/�<�����}M�E�'�O`&�G�E0HIZ3��T0 k� �,�0	E1 4#Q&�1D"3Q  ��U    � 
�n��*E�+�	/�<�����}M�F+�Oh'�O�E0PIZ3��T0 k� �0�4	E1 4#Q&�1D"3Q  �U    � 
�o��,E�;�	/�������}$=�F3�Ot(�_�E0`JZ3��T0 k� �8�<	E1 4#Q&�1D"3Q  ��U    � 
�p��-E�C�	�������}(=�F7�O|)�c�E0dKZ3��T0 k� �<�@	E1 4#Q&�1D"3Q  ��U    � 
�q��/E�K�	�������},=�F;�O�*�k�E0lKZ3��T0 k� �@�D	E1 4#Q&�1D"3Q  ��U    � 
�r��0E�S�	�������},=�F?�O�+�s�E0pLZ3��T0 k� �@�D	E1 4#Q&�1D"3Q  ��U    � 
�s��1E[�	�������}0=�FG�O�+�{�E0xMZ3��T0 k� �D�H	E1 4#Q&�1D"3Q  ��U    � 
�t��3Ek�	�������}8��FO�O�-���E@�NZ3��T0 k� �L�P	E1 4#Q&�1D"3Q  ��U    � 
�u��5Es�	/��������<��FS�O�.ϓ�E@�OZ3��T0 k� �L�P	E1 4#Q&�1D"3Q  ��U    � 
�v��6E{�	/��������<��F[�O�.ϛ�E@�PZ3��T0 k� �H�L	E1 4#Q&�1D"3Q  ��U    � 
�w� 7E��	/��������@��F_�O�/ϣ�E@�QZ3��T0 k� �L�P	E1 4#Q&�1D"3Q  ��U    � 
�x�8E��	/��������D��E�g�B��0ϫ�E@�RZ3��T0 k� �P�T	E1 4#Q&�1D"3Q  ��U    � 
�y�:E��	/��������L��E�o�B��1ϻ�E@�TZ3��T0 k� �X �\ 	E1 4#Q&�1D"3Q  ��U    � 
�z�;E��	��������P��E�w�B��2���E@�UZ3��T0 k� �\"�`"	E1 4#Q&�1D"3Q  ��U    � 
�|� <E��	��������T��E��B��3���E@�VZ3��T0 k� �`$�d$	E1 4#Q&�1D"3Q  ��U    � 
�}�$=E��	��������X��B���B��3���E@�WZ3��T0 k� �d%�h%	E1 4#Q&�1D"3Q  ��U    � 
��,>E��	��������\�B���B��4���E@�XZ3��T0 k� �h&�l&	E1 4#Q&�1D"3Q  �U    � 
���0?E��	��������`�B���@�5 ��E@�YZ3��T0 k� �l'�p'	E1 4#Q&�1D"3Q  ��U    � 
���4@E× o��������d�B���@�5 ��E@�ZZ3��T0 k� �p(�t(	E1 4#Q&�1D"3Q  ��U    � 
���<AE˘ o���� ��h�B���@�6 ��E@�[Z3��T0 k� �p)�t)	E1 4#Q&�1D"3Q  ��U    � 
���@BEә o���� ��l�@��@�7 ��E@�[Z3��T0 k� �t*�x*	E1 4#Q&�1D"3Q  ��U    � 
���DCEי o���� ��p�@��@�7 �E@�\Z3��T0 k� �x+�|+	E1 4#Q&�1D"3Q  ��U    � 
���LDA�ߚ o���� ��t#�@��@ 8 �J��]Z3��T0 k� �|,��,	E1 4#Q&�1D"3Q  ��U    � 
���PEA�� o���� ��|'�@��@9 �J��^Z3��T0 k� ��-��-	E1 4#Q&�1D"3Q  ��U    � 
���TFA�� o���� #�̀ '�@��@9 �J��_Z3��T0 k� ��.��.	E1 4#Q&�1D"3Q  ��U    � 
���XGA�� o���� '�̈́!+�@��@: '�J� `Z3��T0 k� ��/��/	E1 4#Q&�1D"3Q �U    � 
���`HA��� o���� /��"/�@��@: /�J�aZ3��T0 k� ��0��0	E1 4#Q&�1D"3Q ��    � 
���dHA��� o���� 3��#3�@��@ ; 7�J�bZ3��T0 k� ��2��2	E1 4#Q&�1D"3Q ��    � 
���hIA�� o���� 7��$3�@��@$; ;�J�bZ3��T0 k� ��3��3	E1 4#Q&�1D"3Q ��    � ���lJA�� o���� ?��%7�@��@(< C�J�cZ3��T0 k� ��5��5	E1 4#Q&�1D"3Q ��    � ���pKA�� o���� C��&;�@��@0< K�J�dZ3��T0 k� ��6��6	E1 4#Q&�1D"3Q ��    � ���xLA�� o���� G��&?�@��@4= S�J� eZ3��T0 k� ��8��8	E1 4#Q&�1D"3Q ��    � ���|MA�� o���� O��'-C�@��@<> W�J�(eZ3��T0 k� ��9��9	E1 4#Q&�1D"3Q ��    � ����MA�� o���� S�-�(-G�@��@@> _�J�,fZ3��T0 k� ��:��:	E1 4#Q&�1D"3Q ��    � ����NA�#� o���� W�-�)-K�@��@D? g�J�0gZ3��T0 k� ��<��<	E1 4#Q&�1D"3Q ��    � ����OA�+� o���� [�-�*-O�@��@L? k�J�8hZ3��T0 k� �=�=	E1 4#Q&�1D"3Q ��    � ����PA�/� o���� _�-�+-S�@��@P@ s�J�<hZ3��T0 k� �?�?	E1 4#Q&�1D"3Q ��    � ����PA�3� o���� g�-�+-W�@�@T@ w�J�@iZ3��T0 k� �@�@	E1 4#Q&�1D"3Q ��    � ����QA�;� o���� k�-�,-[�@�@XA �J�DjZ3��T0 k� �$B�(B	E1 4#Q&�1D"3Q	 ��    � ����RA�?� o���� o�-�--_�@�@`A ��J�HkZ3��T0 k� �0C�4C	E1 4#Q&�1D"3Q	 ��    � ����RA�C� o���� s�-�.-c�@�@dA ��J�PkZ3��T0 k� �<D�@D	E1 4#Q&�1D"3Q
 ��    � ����SA�G� o��� w�-�/-g�@ @hB ��J�TlZ3��T0 k� �HF�LF	E1 4#Q&�1D"3Q
 ��    � ����TA�K� o��� {��/�o�@@lB ��J�XmZ3��T0 k� �TG�XG	E1 4#Q&�1D"3Q
 ��    � ����UA�O� o��{� ��0�w�@@pC ��J�\mZ3��T0 k� �\I�`I	E1 4#Q&�1D"3Q ��   � ����UA�W� o��{� ���1� @ @tC ��J�`nZ3��T0 k� �hJ�lJ	E1 4#Q&�1D"3Q ��    � ����VA�[� o��w� ���1�@$@xD ��J�dnZ3��T0 k� �tL�xL	E1 4#Q&�1D"3Q ��    � ����VA�_� o��w� ���2�@(@�D ��J�hoZ3��T0 k� ��M��M	E1 4#Q&�1D"3Q ��    � ����WA�c� o��s� ���3�@,@�E ��J�lpZ3��T0 k� ��N��N	E1 4#Q&�1D"3Q ��    � ����XA�g� o��s� ���4�	@0@�E ��J�ppZ3��T0 k� ��P��P	E1 4#Q&�1D"3Q ��    � ����XA�k� o��o� ���4�@4@�E ��J�tqZ3��T0 k� ��Q��Q	E1 4#Q&�1D"3Q ��    �  ����YA�o� o��o� ���5�@8@�F ��J�xqZ3��T0 k� ��S��S	E1 4#Q&�1D"3Q ��    � !����YA�s� o��k� ���6�@<@�F ��J�|rZ3��T0 k� ��T��T	E1 4#Q&�1D"3Q ��    � "����ZA�w� o��k� ���6��@@@�F ��J��sZ3��T0 k� ��V��V	E1 4#Q&�1D"3Q ��    � #����[A�{� o��g� ���7��@D	@�G ��J��sZ3��T0 k� ��W��W	E1 4#Q&�1D"3Q ��    � $����[A�� o��g� ���7��@H
@�G ��J��tZ3��T0 k� ��X��X	E1 4#Q&�1D"3Q ��    � %����\A��� o��g� ���8��@L
@�H ��J��tZ3��T0 k� ��Z��Z	E1 4#Q&�1D"3Q ��    � &����\A��� o��c� ���9��@P@�H ��J��uZ3��T0 k� ��[��[	E1 4#Q&�1D"3Q ��    � ' ��]A��� o��c� ���9��@P@�H ��J��uZ3��T0 k� � ]�]	E1 4#Q&�1D"3Q ��    � ( ��]A��� o��_� ���:��@T@�I ��J��vZ3��T0 k� �^�^	E1 4#Q&�1D"3Q ��    � ) ��^A� o��_� ����:��!@X@�I ��J��vZ3��T0 k� �`�`	E1 4#Q&�1D"3Q ��    � * 
��^A� o��_� ����;��#@\@�I ��J��wZ3��T0 k� � a�$a	E1 4#Q&�1D"3Q ��   � + ��]A� o��[� é� ;� %@`@�J ��J��wZ3��T0 k� �,b�0b	E1 4#Q&�1D"3Q ��    � , ��]A� o��[� Ǩ� <�'@d@�J ��J��xZ3��T0 k� �8d�<d	E1 4#Q&�1D"3Q ��    � - ��]A� o��[� Ǩ�=�)@d@�J ��J��xZ3��T0 k� �De�He	E1 4#Q&�1D"3Q ��    � . ��]A� o��W� ˧�=�*@h@�K ��J��yZ3��T0 k� �Pg�Tg	E1 4#Q&�1D"3Q ��    � / ��\A� o��W� ϧ�>�,@l@�K �J��yZ3��T0 k� �Xh�\h	E1 4#Q&�1D"3Q
 ��    � 0 ��\A� o��S� Ӧ�>� .@p@�K �J��zZ3��T0 k� �dj�hj	E1 4#Q&�1D"3Q
 ��    � 1 ��\A� o��S� Ӧ�?�(0@t@�L �J��zZ3��T0 k� �pk�tk	E1 4#Q&�1D"3Q
 ��    � 2 "��\A� o��S� ץ�?�(0@t@�L �J��zZ3��T0 k� �|m��m	E1 4#Q&�1D"3Q	 ��    � 3 %��[A� o��O� ۥ�@�02@x@�L �J��{Z3��T0 k� ��n��n	E1 4#Q&�1D"3Q	 ��    � 4 (��[A� o��O� ۤ�A�43@|@�L �J��{Z3��T0 k� ��o��o	E1 4#Q&�1D"3Q ��    � 5 +��[A� o��O� ߤ�B�<5@|@�M �J��|Z3��T0 k� ��q��q	E1 4#Q&�1D"3Q ��    � 6 .� [A� o��O� ��B�D6@�@�M �J��|Z3��T0 k� ��r��r	E1 4#Q&�1D"3Q ��    � 7 1� [A� o��K� ��C�H7@�@�M #�J��|Z3��T0 k� ��t��t	E1 4#Q&�1D"3Q ��    � 8 4�ZA�ò o��K� ��D�P9@�@�M '�J��}Z3��T0 k� ��u��u	E1 4#Q&�1D"3Q ��    � 9 7�ZA�ò o��K� ��D�T:@�E��M +�J��}Z3��T0 k� ��w��w	E1 4#Q&�1D"3Q ��    � : :�ZA�ǳ o��G� ��E�\<@�E��M /�J��~bs��T0 k� ��x��x	E1 4#Q&�1D"3Q ��    � ; =�ZA�˳ o��G� ��F�d=@�E��M /�J��~bs��T0 k� ��y��y	E1 4#Q&�1D"3Q ��    � < @�ZA�˳ o��G� �� G�h>@�E��M 3�J��~bs��T0 k� ��{��{	E1 4#Q&�1D"3Q ��    � < C�ZA�ϴ o��C� �� G�p@@�E��M 7�J��bs��T0 k� ��|� |	E1 4#Q&�1D"3Q ��    � < F�ZA�Ӵ o��C� ��� H ntA@�E��N ;�J��bs��T0 k� �~�~	E1 4#Q&�1D"3Q ��    � < I�ZA�Ӵ o��C� ���$I nxB@�Ep�N ?�J�؀bs��T0 k� ��	E1 4#Q&�1D"3Q ��    � < L�ZA�״ o��C� ���$I n�D@�Ep�N ?�J��bs��T0 k� ��� �	E1 4#Q&�1D"3Q ��    � < O�ZA�۵ o��?� ���$J n�E@�Ep�N C�J��bs��T0 k� �(��,�	E1 4#Q&�1D"3Q ��    � < R� [A�۵ o��?� ���(K n�F@�Ep�N G�J��bs��T0 k� �4��8�	E1 4#Q&�1D"3Q  *�    � < U� [A�ߵ o��?� ��(K n�G@�Ep�N K�J��bs��T0 k�  @��D�	E1 4#Q&�1D"3Q  /�    � < X�$[A�ߵ o��?� ��(L n�H@�Ep�O K�J��~bs��T0 k�  H��L�	E1 4#Q&�1D"3Q  ��    � < [�([A�� o��;� ��,L n�J@�E`�O O�J��~Z3��T0 k�  T��X�	E1 4#Q&�1D"3Q  ��    � < ^�,[A�� o��;� ��,M n�K@�E`�P S�J��~Z3��T0 k�  `��d�	E1 4#Q&�1D"3Q  ��   � < a�,[A�� o��;� ��,N n�L@�E`�P S�J��~Z3��T0 k�  l��p�	E1 4#Q&�1D"3Q  ��    � < d�0[A�� o��;� ��,N n�M@�E`�Q W�J��}Z3��T0 k� �x��|�	E1 4#Q&�1D"3Q  ��    � < g�4[A�� o��7� ��0O n�N@�E`�R [�J��}Z3��T0 k� ������	E1 4#Q&�1D"3Q  ��    � < j�4\A�� o��7� ��0O n�O@�E��R [�J��}Z3��T0 k� ������	E1 4#Q&�1D"3Q  ��    � < m�8\A�� o��7� ��0P n�P@�E��S _�J��}Z3��T0 k� ����	E1 4#Q&�1D"3Q  ��    � < p�<\A�� o��7� ��4P n�Q@�E� T c�J��|Z3��T0 k� ����	E1 4#Q&�1D"3Q  ��    � < s�<\A�� o��7� ��4Q n�R@�E� U c�J��|Z3��T0 k� ����	E1 4#Q&�1D"3Q  ��    � < v�@\A��� o��3� ��4Q n�S@�E� U g�J��|Z3��T0 k� ���	E1 4#Q&�1D"3Q  ��    � < y�D\A��� o��3� ��4R n�T@�E� V k�J��|Z3��T0 k� ����	E1 4#Q&�1D"3Q  ��    � < |�D\A��� o��3� ��8R n�U@�E�W k�J� |b���T0 k� ��~��~	E1 4#Q&�1D"3Q  ��    � < �H\A��� o��3� ��8S n�V@�E�X o�J� {b���T0 k� ��~��~	E1 4#Q&�1D"3Q  ��    � < ��H]A��� o��3� ��8S n�W@�E�Y o�J� {b���T0 k� ��~��~	E1 4#Q&�1D"3Q  ��    � < ��L]A��� o��/� ��8T n�X@� E�[ s�J�{b���T0 k� ��}��}	E1 4#Q&�1D"3Q  ��    � < ��P]A�� o��/� #��<T n�Y@� E�\ w�J�{b���T0 k� ��}��}	E1 4#Q&�1D"3Q  ��    � < ��P]A�� o��/� #��<U n�Z@� E�] w�J�{b���T0 k� �}�}	E1 4#Q&�1D"3Q  ��    � < ��T]A�� o��/� '��<U n�[@�!E�^ {�J�{b���T0 k� �|�|	E1 4#Q&�1D"3Q  ��    � < ��T]A�� o��/� '��<V n�\@�!E�_ {�J�zb���T0 k� �|�|	E1 4#Q&�1D"3Q  ��    � < ��X]A�� o��+� +��@V n�]@�!E�a �J�zb���T0 k� �$|�(|	E1 4#Q&�1D"3Q  ��    � < ��X]A�� o��+� +��@W n�^@�!E�b �J�zb���T0 k� �,z�0z	E1 4#Q&�1D"3Q  ��    � < ��\]A�� o��+� +��@W n�^@�"H�c ��J�zb���T0 k� �z� z	E1 4#Q&�1D"3Q  ��    � < �1\]A�� o��+� /��@W n�_@�"H�e ��J�zZ3��T0 k� �y�y	E1 4#Q&�1D"3Q  ��    � < �1`]A�� o��+� /��DX o `@�"H�f ��J�zZ3��T0 k� �y�y	E1 4#Q&�1D"3Q  ��    � < �1`^A�� o��+� /��DX oa@�#H�g ��J�yZ3��T0 k� �z�z	E1 4#Q&�1D"3Q  ��    � < �1d^A�� o��'� 3��DY ob@�#H�i ��J�yZ3��T0 k� ��y��y	E1 4#Q&�1D"3Q �    � < �1d^A�� o��'� 3��DY oc@�#Hqj ��J�yZ3��T0 k� ��y��y	E1 4#Q&�1D"3Q ��    � < |1h^A�� o��'� 3��DZ oc@�#Hqk ��J�yZ3��T0 k� ��x��x	E1 4#Q&�1D"3Q ��    � < v1h^A�� o��'� 7��HZ od@�$Hql ��J�yZ3��T0 k� ��x��x	E1 4#Q&�1D"3Q ��    � < p1l^A�� o��'� 7��HZ oe@�$Hqn ��J�yZ3��T0 k� ��x��x	E1 4#Q&�1D"3Q ��    � < j1l^A�� o��'� ;��H[ of@�$Hqo ��J�yZ3��T0 k� ��w��w	E1 4#Q&�1D"3Q	 ��    � < e �p^A�� o��#� ;��H[ of@�$Hap ��J� xZ3��T0 k� ��w��w	E1 4#Q&�1D"3Q
 ��    � < ` �p^A�� o��#� ;��H[ o g@�%Haq ��J� xZ3��T0 k� �v��v	E1 4#Q&�1D"3Q ��    � < [ �p^A�� o��#� ?��L\ o h@�%Har ��J� xZ3��T0 k� �v��v	E1 4#Q&�1D"3Q ��    � < V �t^A�� o��#� ?��L\ o$h@�%Has ��J�$xZ3��T0 k� �u��u	E1 4#Q&�1D"3Q ��    � < Q �t^A�� o��#� ?��L\ o(i@�%Hat ��J�$xZ3��T0 k� �u��u	E1 4#Q&�1D"3Q ��    � < M �x_A�#� o��#� ?��L] o,j@�&Hau ��J�$xZ3��T0 k� �u��u	E1 4#Q&�1D"3Q ��    � < I �x_A�#� o��#� C��L] o0j@�&Hav ��J�(xZ3��T0 k� ��t��t	E1 4#Q&�1D"3Q ��    � < E �|_A�#� o�<#� C��P^ o0k@�&Hav ��J�(wZ3��T0 k� ��t��t	E1 4#Q&�1D"3Q ��    � < A �|_A�'� o�<� C��P^ o4l@�&Hav ��J�(wZ3��T0 k� �xs�|s	E1 4#Q&�1D"3Q ��    � < = �|_A�'� o�<� G��P^ o8l@�&Hav ��J�(wZ3��T0 k� �ps�ts	E1 4#Q&�1D"3Q ��    � < 9 ��_A�'� o�<� G��P^ o8m@�'Hau ��J�,wZ3��T0 k� �ds�hs	E1 4#Q&�1D"3Q ��    � < 5 ��_A�+� o�<� G��P_ o<m@�'Hau ��J�,wZ3��T0 k� �\r�`r	E1 4#Q&�1D"3Q ��    � < 1 ��_A�+� o�<� G��P_ o@n@�'Hau ��J�,wZ3��T0 k� �Tr�Xr	E1 4#Q&�1D"3Q ��    � < - ��_A�+� o�<� K��T_ o@o@�'Ha u ��J�0wZ3��T0 k� �Hq�Lq	E1 4#Q&�1D"3Q ��    � < ) ��_A�/� o�<� K��T` oDo@�'Ha t ��J�0wZ3��T0 k� �@q�Dq	E1 4#Q&�1D"3Q ��    � < & ��_A�/� o�<� K��T` oHp@�(Ha t ��J�0wZ3��T0 k� �8p�<p	E1 4#Q&�1D"3Q ��    � < # ��_A�/� o� �� O��T` oHp@�(Ha t ��J�0vZ3��T0 k� �0p�4p	E1 4#Q&�1D"3Q ��    � <   ��_A�/� o� �� O��Ta oLq@�(A� t ��J�4vZ3��T0 k� �$p�(p	E1 4#Q&�1D"3Q ��    � <  ��_A�3� o� �� O��Ta oPq@�(A� t ��J�4vZ3��T0 k� �o� o	E1 4#Q&�1D"3Q ��    � <  ��`A�3� o� �� O��Ta oPr@�(A� s ��J�4vZ3��T0 k� �o�o	E1 4#Q&�1D"3Q  ��    � <  ��`A�3� o� �� S��Xa oTs@�)A�$s ��J�8vZ3��T0 k� �n�n	E1 4#Q&�1D"3Q! ��    � <  ��`A�7� o� �� S��Xb oTs@�)A�$s ��J�8vZ3��T0 k� � n�n	E1 4#Q&�1D"3Q! ��    � <  ��`A�7� o� �� S��Xb oXt@�)A�$s ��J�8vZ3��T0 k� ��m��m	E1 4#Q&�1D"3Q" ��    � <  ��`A�7� o� �� S��Xb o\t@�)A�$s ��J�8vZ3��T0 k� ��m��m	E1 4#Q&�1D"3Q# ��    � <  ��`A�7� o� �� S��Xb o\u@�)A�$r ��J�8vZ3��T0 k� ��m��m	E1 4#Q&�1D"3Q$ ��    � <  ��`A�;� o� �� W��Xc o`u@�)A�$r ��J�<vZ3��T0 k� ��l��l	E1 4#Q&�1D"3Q% ��    � <  ��`A�;� o� �� W��Xc o`v@�*A�$r ��J�<uZ3��T0 k� ��l��l	E1 4#Q&�1D"3Q% ��    � <  ��`A�;� o� �� W��\c odv@�*A�(r ��J�<uZ3��T0 k� ��k��k	E1 4#Q&�1D"3Q& ��    � <�� ��`A�;� o� �� W��\c odw@�*A�(r ��J�<uZ3��T0 k� ��k��k	E1 4#Q&�1D"3Q' ��    � <�� ��`A�;� o� �� [��\d ohv@�*A�(q ��J�@uZ3��T0 k� ��j��j	E1 4#Q&�1D"3Q' ��    � <�� ��`A�?� o� �� [��\d ohv@�*A�(q ��J�@uZ3��T0 k� ��j��j	E1 4#Q&�1D"3Q( ��    � <�� ��`A�?� o� �� [��\d olv@�*A�(q ��J�@uZ3��T0 k� ��j��j	E1 4#Q&�1D"3Q( ��    � <�� ��`A�?� o� �� [��\d olv@ +A�(q ��J�@uZ3��T0 k� ��i��i	E1 4#Q&�1D"3Q) ��    � <�� ��`A�?� o� �� [��\e opu@ +A�(q ��J�@uZ3��T0 k� ��i��i	E1 4#Q&�1D"3Q* ��    � <�� ��`A�C� o� �� _��\e opu@ +A�(q ��J�DuZ3��T0 k� ��h��h	E1 4#Q&�1D"3Q* ��    � <�� ��`A�C� o� �� _��\e otu@ +A�,p ��J�DuZ3��T0 k� ��h��h	E1 4#Q&�1D"3Q+ ��    � <�� ��`A�C� o� �� _��`e otu@ +A�,p ��J�DuZ3��T0 k� �tg�xg	E1 4#Q&�1D"3Q+ ��    � <�� ��aA�C� o� �� _��`e oxt@+A�,p ��J�DuZ3��T0 k� �lg�pg	E1 4#Q&�1D"3Q+ ��    � <�� ��aA�C� o� �� _��`f oxt@+A�,p ��J�DtZ3��T0 k� �dg�hg	E1 4#Q&�1D"3Q, ��    � <�� ��aA�G� o� �� c��`f o|t@,A�,p ��J�HtZ3��T0 k� �Xf�\f	E1 4#Q&�1D"3Q, ��    � <�� ��aA�G� o� �� c��`f o|t@,A�,p ��J�HtZ3��T0 k� �Pf�Tf	E1 4#Q&�1D"3Q- ��    � <�� ��aA�G� o� �� c��`f o|s@,A�,o ��J�HtZ3��T0 k� �He�Le	E1 4#Q&�1D"3Q- ��    � <�� ��aA�G� o� �� c��`f o�s@,A�,o ��J�HtZ3��T0 k� �@e�De	E1 4#Q&�1D"3Q- ��    � <�� ��aA�G� o� �� c��`g o�s@,A�,o ��J�HtZ3��T0 k� �4d�8d	E1 4#Q&�1D"3Q- ��    � <�� ��aA�K� o� �� c��`g o�s@,A�0o ��J�LtZ3��T0 k� �,d�0d	E1 4#Q&�1D"3Q. ��    � <�� ��aA�K� o� �� g��dg o�s@,A�0o ��J�LtZ3��T0 k� �$d�(d	E1 4#Q&�1D"3Q. ��    � <�� ��aA�K� o� �� g��dg o�r@,A�0o ��J�LtZ3��T0 k� �c�c	E1 4#Q&�1D"3Q. ��   � <�� ��aA�K� o� �� g��dg o�r@-A�0o ��J�LtZ3��T0 k� �c�c	E1 4#Q&�1D"3Q. ��    � <�� ��aA�K� o� �� g��dh o�r@-A�0n ��J�LtZ3��T0 k� �b�b	E1 4#Q&�1D"3Q. ��    � <�� ��aA�K� o� �� g��dh o�r@-A�0n ��J�LtZ3��T0 k� ��b� b	E1 4#Q&�1D"3Q/ ��    � <�� ��aA�O� o� �� g��dh o�r@-A�0n ��J�PtZ3��T0 k� ��a��a	E1 4#Q&�1D"3Q/ ��    � <�� ��aA�O� o� �� k��dh o�r@-A�0n ��J�PtZ3��T0 k� ��a��a	E1 4#Q&�1D"3Q/ ��    � <�� ��aA�O� o� �� k��dh o�q@-A�0n ��J�PtZ3��T0 k� ��a��a	E1 4#Q&�1D"3Q/ ��    � <�� ��aA�O� o� �� k��dh o�q@-A�0n ��J�PsZ3��T0 k� ��`��`	E1 4#Q&�1D"3Q/ ��    � <�� ��aA�O� o� �� k��di o�q@-A�0n ��J�PsZ3��T0 k� ��`��`	E1 4#Q&�1D"3Q/ ��    � <�� ��aA�O� o� �� k��di o�q@.A�4n ��J�PsZ3��T0 k� ��_��_	E1 4#Q&�1D"3Q/ ��    � <�� ��aA�S� o� �� k��hi o�q@.A�4n ��J�TsZ3��T0 k� ��_��_	E1 4#Q&�1D"3Q/ ��    � <�� ��aA�S� o� �� k��hi o�q@.A�4m ��J�TsZ3��T0 k� ��^��^	E1 4#Q&�1D"3Q. ��    � <�� ��aA�S� o� �� o��hi o�p@.A�4m ��J�TsZ3��T0 k� ��^��^	E1 4#Q&�1D"3Q. ��    � <��                                                                                                                                                                            � � �  �  �  d A�  �K����   �      6 \��g\ ]�&&
 8 �) `t�   � �
	  �����     `Us��+�     ��              /	 Z��           ���  &  ���  (
	           ^�  > > 
	   ���<~     ^�4��c�     �             Y	 Z��          � �     ���   
	           GZb   � �
     ���     Gq����    �� �   
         8  Z��           ��  $  ���  8	 

          PCS   : :     ���     PB���@�      �!               	 Z��          ��    ���  0
3
          _&�   * *	     /�yA(     _rn�y?]    �� �                 Z��           +0�     ���   H


          �H  ��    C�}.     �H�}.                            ���I              ^  ���    		 5 	           ���p         W�H|H    �����H|H    ��             
 
            �     ��@   0
&


          X�R       k�;m<     X}��;m<     Q             
 
 �          !�     ��@   (
 
           ?(Q $ $     ��o�     ??���W    ��q                �         q�     ��@   0	
           )��        ��.W�     )�f�.sN     �a                  T         	        ��H   H	$
          6�         ���l�     6���`�    �� �                 ��         
 �     ��@   03 
            ����     � ��7      �� ��7                             ���4              ^  ��@   P		 5                   ��      �                                                                           �                               ��        ���          ��                                                                 �                         ���?  ��        ����!    �������Z    �	�W "                  x                j  �   �	   �                         ��    ��        ���      ��  ��           "                                                 �                         ���������y��H�;���.�� ������� 
   	             
  C   �p� h��A       �� �[� �� \� � ]  �$ ]  �D ]@ �d ]`���J ����X ����� � �� ]� �� ]����. ����< ����J ����X � �� u� � �r` �  s` 
�\ V� 
� W  
�\ W  �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0� ���� ����� � � �r` � s` � s� �� �o� �� p� � q  �$  q  �d q` �� q� �� �j� �� k� @� 0e� @� @f@ Ad f� A� @f� B  g` �d 0t� �� 0u@ �$ u� �D  u� ��  v  Ƥ �h` Ǥ i` ��  i� � �m` �  n` �d  }� �� }����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������� �� y  ������  
�fD
��L���"����D"� �  " `   J jF��     �j   
��
��
���    "�j��" " �
� �  �  
�  '    ��     ��R  �    G    ��     ���       )    ��     ��.          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �/$ $      ��D �  ���        �O �  ���        �        ��        �        ��        � 	 	 �     "������        ��                         T�) , ��� �                                     �                  ����           	 '�S 	���&��   �� 2 F�2       �     9 Pelle Eklund        1:54                                                                        4  3     �s � �r � �S CC �[CD �s CJ �[CK �2c�J c� �$	kk12
ks!cW �- c_ � �C/: � C72 � C82 �J�8 � J�0 �C. � C!. � C"> �B�9 � B�I � B�1 � B�4 � B�: � B�< �C  �C �C0 �k� �k� � � k � !k�* �""� � #"�/ �$"� �%*�(T&"� �T '"�D(� �D 
�
B*� �B 
�
/,� �/ 
�	, 
�	+ 
�	*0� �* 
�	*2� �* 
�	 �{ � 5"�9 �6"�# �7*�2,8"� �, 9"�:� � 
�X  *LU.  "Q v6 >"E vN  "S v                                                                                                                                                                                                                         �� R        �     @ 
             ^ P E g  ��        	            ������������������������������������� ���������	�
���������                                                                                          ��    �g�� ��������������������������������������������������������   �4, ?   6 � � � @(�@<@���A+��2�J�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             2    2    �� 
İJ          	                           ������������������������������������������������������                                                                   
                                                	                   ����  �  �                                           ���������������� �������� �������� ������������������������������������������� ���������������� ������������ � �������������  �������������� �������������������� ��������������  � ���������������������� �������� ������������������  �                    	      
        c    -     � ��J     �U                              ������������������������������������������������������                                                                                                                                        ����  ��                                             � ������������������������������ ������������������� ��������������������� ������� ������������������������ ����� ��� ����� ������� �������������������� ������������������������ ���������� ������  � �������������� ������ ��� �������                                                                                                                                                                                                                                           	          
                                                                      �              


             �  }�           �  0�             M     M                                                      ���      K  g�����  W  8�����������������������������������������������������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � ���� �[�                                                                                                                                                                                                                                                                                           )n)n1n  	n�              k      b      m      d      k      m                                                                                                                                                                                                                                                                                                                                                                                                                > �  
>�   J�   Q  (�  Cm�  ��8�� �N \�̞����&�[�̎���˶���̞�J��� �                      �: {        $   �   & QW  �   l                  �                                                                                                                                                                                                                                                                                                                                      0 K K   �                       !��                                                                                                                                                                                                                            Z��   �� �� �      �� M      ���������������� �������� �������� ������������������������������������������� ���������������� ������������ � �������������  �������������� �������������������� ��������������  � ���������������������� �������� ������������������  �� ������������������������������ ������������������� ��������������������� ������� ������������������������ ����� ��� ����� ������� �������������������� ������������������������ ���������� ������  � �������������� ������ ��� �������             $����������������UUUU�����UUU�U{�����������������UUUW����x�����w�����������������UUuU������wxwwww����������������WwwU�������wwwwx����������������UUUU����w�xw�w������������������Uuww���uUw��uU���Uz��uz��Wz��wzu�wYW�wxw�uxwwuW���������wx��UUwwX�xuy����u������wwww�wwwwwwwwwwwUUwWuUuu�UWW�wwwwy��x���x���ww�uwuuwwx��x�����Y����������w��www�wwwy��wyx�wyx��x�U���U���U���uy��u���u��uu��uU���wx��wxxwuW�WuuxU�uWW�UUU�uWu��W�y���wx�ww��wxx����wwwwwWwwwwwuW��ww��wx��w��xww��WwxUW�wWW�wy����w����������x�www��xwx�w��w�Ww����w��xwx�xwwwx�xwww��ww�wwwwwww�Wy�x�xuw��UwuwWwuwWwxwX�xwW�wuW�z�u�Y�u�X�u�U��yUU�Uuw�yUX��UX�uWwuWuwWwUwwUUUwUUWUUUUuUUWWUUWwwuW�WUW�XUuwx�UXx�Uxwwwxww�xww����ww��UwuwwW��ww��ww��ww��xw��xwwwwwwwwwwwwxwwwxuwwxwwwwUwwwWwwwwywX��yWx�Xxy�W��uXYwWuZ��u��w���ux���w���U���U���U���u���UZ��UWUUwWuUUU�Uu��Uw��UWx�UUW��UU��UUwwwxUwww��wx��������x���w���Ux�wx�wwwwww���w���U��ww��ww�wwwuwwwWwwxWwwywww�wwx�ww��xx��wx��w����WU��WY��uY��Wx��Wy�Uxz�Xw��Xw�W���W���U��������������������������UUW�uUUX�U�U�W�uWW��WU���u���WUUUWUUwuuwwwwx��wwx�wwwwwwwwuwwwWuwwWwwwuwwx�ww�wwwx�w�xxw��wx��xw�Uw��W���Xx�U��uW��UxwUWwwUwww�w�W�x�W�y�wx��wx�Wwx�Wyz�wz��x�q��    B      0   � ��                       M     �  �����J���J'    ��     ~         �      �   �      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ��  � ��     � ��  � ��  p �� �� �z  p���� �$ ^h  ��  p  ����     �           �� �     ��  H ��   �� �� �z  ���� �$ ��  n ��     �� �� �� ��  �� �� [� �� �� �z [� �� �$  �q  �� I      �  ��   �������2����  g���  �     f ^�         ��              ��g����2�������J��(2���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                         E  �\       U TUTQ�T\�jA���̪������ UTDDEUU�����j������������������DUP UUTD�����v����������������    U�UPUDDE��\����������������        U   TE ��@ x�@ �lE �|U  E� \� �Q� _ǪE�L��\��\�������������������E�lTP��E ��P �����������UDL�_UL�_L�UL�L�̪�������U������D���EU��E��E���E���������z��Q�j�T_�z �_�  T\  E��U ��T ����|��E |P �E  @  \��\��\��Ez� Oʪ UǪ \� Eʪ�P ��E �|�P���D��lϪ�����������L��L��L�UUL�QDL�_���Ua��̪��w���E��EU��E���E��DU�����wz��   �  �E �ETOQ���j����������UO  �T  ��P ��O ��� �����O���E  T\  E   T                   ����Ǫ��\ʪ�E\ʪUE\� UDU  UT    ����������������z������DUUUUTD�������������������|���UUTDDUU�����������̧|�T�TUUDP U       ��TQ�TE TE  E                   wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwtwwwCwwt1wwCwt1wC�t1��C1����������""""���������������!���""!����,���ww��7����������������wwwwwwwwwwwwwwwwwwww7wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwws��w1wt1�wC�t1��s��s��s������"$��Gw�!������������L���q��"r��������!�����!ww�r�w�ww!�wwrwwwwwwqwwwrwwww�7ww�ww�ww��7w��w���G��'!wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                 �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "" "  """     " ""   "" !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ "!    " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """     " ""   "" !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                             �   �   �   r�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  bp gp �'������ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     "  �           �   �   �                     .  ". "  ""                       "  .���"    �     �                                               ���                          ����                  �   �� �       �  �  "�  "   "                                             � 
��	�˽���w��rb��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            .  .     �   �           / �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��  .�"." "."   /�  �  �              � ��         �� �� �� g} &' vw     ���.�                     �"�!/"�  �                                                                                                                                                                                 ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   �"   ".   .                  �   �   �   �   �   �   �   �                .         �  �  �  �                                  � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                                       � �� �������ۛ˽���� �ͼ ��+ �""�B.�R#Z�C U�D �T Z� �; � �� ��� ��  ��� ˽� �wp �&  �vp �w� ��� ˙� ̻� �۰ �ِ ��� Ш� �� >�" 3��.30" ��  �   �                �"/ "" ""  ��  ��                       .  .  "   "       �          �  �" �"" �"   �                    .   .   �            �  "�  "  "  �   �         �        �   �     �       �       "       .      �                    �"  �""� "�                        ����                               ���                          ����                  �   �� �       �  �  "�  "   "                                                                  
   �   �  ��  �� ������-�� "��  �  
�  �C 
UU US �UD TE0 �� 
�� ʐ �  ̻  "�  "   " �� ����   �  �˰ ̻� �ݰ �w� ��� ����������˹�̹���ڙ��ٻ��ݰ̻� ˘  ��  3D  TD� 340 340 3D0 30 
��  ��  "/  "/  �� ���� �    ��                  "      �              "   "   "�  �            ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �                    �"  �""� "����                                                                                                                                                                                                             �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �         �� �� �� �� �݉���̙�  ���                              �������  �                     �  .   .     �   �  ��  �                                                                                                                                                                                                   �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���                            "  ""�����"    /   �  �   ��                         �    �                    .   .                    �EU �E  
�   �               �"�!/"�  �                       � ".��".��/����  �                                                                                                                                                              	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           "� /���  �       �   �   �                                                   ��  ����   �       �                                   �    ��"  �"                    ".  ".  ���                        "  "  "      � ".��".��/����  �                                                                                                                                             �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   �   " � ��      �    �      �                         ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �                            � ��       "   "   "�  �                            �   ���                            �   "                                                                                                   �� ��� ��� ww� &'� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                               " "/ �/� ��             �   "   "  "                 �   �   "   "�  �                    �� ��� ��� ����                            �                               � ��       "   "   "�  �                            �   ���                            �   "                                                                                                                         	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           "� /���  �       �   �   �                         �   �     �   �        �   �"/� ����                                     �"  �"  �                  �  ".��".� ��                        ���                                                                                                                                                                                                   �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ���������""��""��""�����        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                   2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��   �  �   
�  �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                             "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�GwDGwqwDDwtwwww3333DDDD �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�""""����������A��I��I = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=""""�����A�DA�I��I�    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"��������I���I���I���I��� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(XxMAMAMMMM�M�M����3333DDDD w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xwwD�����MD��M����3333DDDD  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���4���4���4���4���4���43334DDDD �  + � � � � � � � � � � ��	� � � ��� � � � � � � � � � � ��	� � � ��� �� ����(+((�""""wwwwqqqqwGwGGG ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""wwwwwwqqDAwG M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M������������������333DDD � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�M��M��D��M����������3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DD��D�M��D����3333DDDD 5 6  X � �F � � � � � ����� � ����������� � ����� � � � � ��	F ��(X((6(5""""������DH�H� x �  l � �G � � � � � � � � � � ������������� � � � � � � � � � ��	G ��l((�x""""�������H�H��D!�!�!�5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�vw��(W(�""""��������H��H��H��H�� !�!�AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���&2�(a(�DD������L��DL����3333DDDD;'(!�AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(�L�A�AAD��DL�����3333DDDD<34!�AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� SA��l(=���4���4���4L��4L��4���43334DDDD  � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� SA��(( """"���������M�MMM X � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� SA��(Xx""""�������A��AA w � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� )��:	9ww��������������333DDD � � �!�AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(I��I����������������3333DDDD  � �!�AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((���A���I��I���I�����3333DDDD m � �!�A�A� � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""������������������������  � �!�AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M""""������D�D��� 
 � �!�AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�""""������������������������ - � �!�!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�wqwwqwwwwwqwwwDwwww3333DDDD 69�:���  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5qqwwwDDwtGwwww3333DDDD x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xwww4www4www4www4www4www43334DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwqwwwqwqwq + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""wwwwwwwDwGwA � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(��A�L�L�L��L���333DDDLDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDDs � �r � �S CC �[CD �s CJ �[CK �2c�J c� �$	kk12
ks!cW �- c_ � �C/: � C72 � C82 �J�8 � J�0 �C. � C!. � C"> �B�9 � B�I � B�1 � B�4 � B�: � B�< �C  �C �C0 �k� �k� � � k � !k�* �""� � #"�/ �$"� �%*�(T&"� �T '"�D(� �D 
�
B*� �B 
�
/,� �/ 
�	, 
�	+ 
�	*0� �* 
�	*2� �* 
�	 �{ � 5"�9 �6"�# �7*�2,8"� �, 9"�:� � 
�X  *LU.  "Q v6 >"E vN  "S v3333DDDDAqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD��������������������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ��������������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ��������������������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE��������������������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD��������������������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD��������������������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD��������������������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� ����7�\�J��<�V�I�P�[�H�P�S�S�L�������8�>�7���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� ����>�L�L�T�\��=�L�S�H�U�U�L��������>��<���""""������A�D��I��""""�������D����� ��%��:�L�S�S�L��0�R�S�\�U�K���������8�>�7���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �>��<��� ���A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �8�>�7���!��""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,�����������DDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II�""""������D""""������IADD���I""""��������D��""""�������I��I�I�I�""""�������A�D�II�I""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            