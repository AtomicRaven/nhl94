GST@�                                                            \     �                                               ���      �  ��  K         ���2�������ʱ�����������������        i     #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    "�j��,  " ��
  D                                                                               ����������������������������������       ��    =b= 0Q0 44 111  4            	 
                    ��� �� � � ��                 nn 	)
         8�����������������������������������������������������������������������������������������������������������������������������  bb    41  c  c  c                   	  
        G  �  (  (                  n�  1)          8= �����������������������������������������������������������������������������                                �          �   @  &   �   �                                                                                 '    	n)n
  1n)�    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    AP7�ARS�PHq ��&+�|/�n�OLN�bLaP *�k"��T0 k� ����U2d  U8D"!  ��?    � ��AP7�ARS�PHq ��&+�|/�n�OLN�cLbP *�k"��T0 k� ����U2d  U8D"!  ��?    � ��AP3�ARS�PHq ��&+�|/�n�OLN�cLcP *��k"��T0 k� ����U2d  U8D"!  ��?    � ��AP3�ARS�PHq ��&+�|/�n�OLN�dLdP *��k"��T0 k� ����U2d  U8D"!  ��?    � ��AP3�ARS�PHq ��&+�|/�n�OLN�dLeP *��k"��T0 k� ����U2d  U8D"!  ��?    � ��AP3�ARS�PHq ��&+�|/�n�OLN�eLfP *��k"��T0 k� ����U2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&+�|/� ��OLN�eLgP *��k"��T0 k� ����U2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&+�|/� ��OLN�fLiP *��k"��T0 k� �߬��U2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&+�|/� ��OL>�fL jP *��k"��T0 k� �߫��U2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� ��OL>�gL kP *��k"��T0 k� �۫�߫U2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� ��OL>�gL�lP *��k"��T0 k� �۪�ߪU2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� ��OL>�gL�mP +�k��T0 k� �ש�۩U2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� n�OL>�hL.�n_�+�k��T0 k� �ө�שU2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� n�OL>�hL.�o_�+�k��T0 k� �Ө�רU2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� n�OL>�iL.�p_�+�k��T0 k� �Ϩ�ӨU2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� n�OL>�iL.�q_�+�k��T0 k� �ϧ�ӧU2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� n�OL>�iL.�r_�+�k��T0 k� �˦�ϦU2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� n�OL>�jL.�s_�+�k��T0 k� �˦�ϦU2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� n�OL>�jL.�s_�+�k��T0 k� �ǥ�˥U2d  U8D"!  ��?    � ��AP3�ARO�PHq ��&'�|/� n�OL>�jL.�t_�+�k��T0 k� �å�ǥU2d  U8D"!  ��?   � ��AP3�ARO�PHq ��&'�|/� n�OL>�jL.�u_�+�k��T0 k� �ä�ǤU2d  U8D"!  ��?    � ��AP/�ARO�PHq ��&'�|/� n�OL>�jL.�v_�+��k��T0 k� ����ãU2d  U8D"!  ��?    � ��AP/�ARO�PHq ��&'�|/� n�OL>�jL.�w_�+��k��T0 k� ����ãU2d  U8D"!  ��?    � ��AP/�ARO�PHq ��&'�|/� n�OL>�jL.�x_�+��k��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARO�PDq ��&'�|/� �OL>�jL.�y�+��k��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARO�PDr ��&'�|/� �OL>�jL.�z�+ |j��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARO�P@r ��&'�|/� �OL>�jL.�z�+ xj��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARO�P<r ��&'�|/� �OA��jL.�{�+ tj��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARO�P<r ��&#�|/� �OA��jL.�|�+ tj��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARO�P8s ��&#�|/� �OA��jL.�}�+ pi��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARO�P8s ��&#�|/� �OA��jL.�}�+ li��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�P4s ��&#�|/� �OA��jL.�~�+ hi��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�P0s ��&#�|/� �OA��jL.��+ di��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�P0t ��&#�|/� �OBN�jL.܀�+ `i��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�P,t ��&#�|/� �OBN�jL.��+ \h��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�P,t ��&#�|/� �OBN�jL.��+ \h��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�P(t ��&#�|/�N�OBN�jL.��+Xh��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�P$u ��&#�|/�N�OBN�jL.��+Th��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�P$u ��&#�|/�N�O@�jL.�~/�+Ph��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�P u ��&#�|/�N�O@�jL.�~/�+Lg��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�P v ��&#�|/�N�O@�jL.�~/�+Dg��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�Pv ��&#�|/�N�O@�jL.�~/�+@g��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�Pv ��&#�|/�~�O@�jL.�~/�+8g��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�Pv ��&#�|/�~�O@n�jL.�}/�+4g��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�Pw ��&#�|/�~�O@n�jL.�}/�+0f��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�Pw ��&#�|/�~�O@n�jL.�}/�+(f��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�Pw ��&#�|/�~�O@n�jL.�}/�+$f��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�Pw ��&#�|/�~�O@n�jL.�|/�+�f��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�Pw ��&#�|/�~�OB��jL.�|/�+�f��T0 k� ������U2d  U8D"!  ��?    � ��AP/�ARK�Px ��&#�|/�~�OB��iL.�|/�+�f��T0 k� ������U2d  U8D"!  ��?    � ��AP+�ARK�Px ��&#�|/�~�OB��iL.�|/�+�e��T0 k� ������U2d  U8D"!  ��?    � ��AP+�ARK�Px ��&#�|/�~�OB��iL.�|/�+� e��T0 k� �����U2d  U8D"!  ��?    � ��AP+�ARK�Px ��&#�|/�~�OB��hL.�{/�+��e��T0 k� �����U2d  U8D"!  ��?    � ��AP+�ARK�Py ��&#�|/�~�OB��hL�{/�+��e��T0 k� �{���U2d  U8D"!  ��?    � ��AP+�ARK�Py ��&#�|/�~�OB��hL�{/�+��e��T0 k� �{���U2d  U8D"!  ��?    � ��AP+�ARK�P y ��&#�|/�~�OB��gL�{/�+��e��T0 k� �w��{�U2d  U8D"!  ��?    � ��AP+�ARK�P y ��&#�|/���OC�gL�{/�+��e��T0 k� �w��{�U2d  U8D"!  ��?    � ��E,EB��w��.��|/�r��IlgI�����o����T0 k� ����U2d  U8D"!  ��    ��� E�4DB��{��,��|/�r��IpgI�����s����T0 k� ����U2d  U8D"!  ��    ��� E�<DBì���+��|/�r��ItgI�����w����T0 k� ��ÿU2d  U8D"!  ��    ��� E�PDB˰���)��|/����I"xgI!��C��{����T0 k� ������U2d  U8D"!  ��    ��� E�XDB˱	2��� (�#�|/����I"|gI!��C������T0 k� ������U2d  U8D"!  ��    ��� E�`DBϳ	2���('�+�|/����I"�gI!��C#�	�����T0 k� ������U2d  U8D"!  ��    ��� E�hDBӵ	2���,%�/�|/����I"�gI!��C'�	�����T0 k� ������U2d  U8D"!  ��    ��� E�pDB׶	2���4$�3�|/����I"�gI!��C+�	�����T0 k� ������U2d  U8D"!  ��    ��� E�|DB۸	2���8#�7�|/��I�gE��C+�	�����T0 k� ������U2d  U8D"!  ��    ��� E��DEc߼	2���D!�C�|/��I�gE��C3�
�����T0 k� ������U2d  U8D"!  ��    ��� E��DEc�	B���L �G�|/��I�gE��C7�
�����T0 k� ������U2d  U8D"!  ��    ��� E��DEc�	B���TK�|/�#�I�gE�S;�
�����T0 k� ������U2d  U8D"!  ��    ��� Es�EEc��	B���XO�|/�+�I"�gE�S?�
�����T0 k� �����U2d  U8D"!  ��    ��� Es�EEc��	B���`S�|/�/�I"�gE�S?�
�����T0 k� �����U2d  U8D"!  �    ��� Es�EE���	B���l_�|/��?�I"�gE�SG������T0 k� #�����U2d  U8D"!  ��    ��� Es�FE������tc�|/��G�I"�gE'�SK������T0 k� #�����U2d  U8D"!  ��    ��� Es�FE���� �xg�|/��K�I�gE�+�SK������T0 k� #�����U2d  U8D"!  ��    ��� Es�GE���� ��k�|/��S�I�gE�3�SO������T0 k� #�����U2d  U8D"!  ��    ��� D��GE������s�|/��[�I�gE�;�SS������T0 k� #�����U2d  U8D"!  ��    ��� D��HE������{�|/��k�I�gE�G�#W������T0 k� #�����U2d  U8D"!  ��    ��� D��IE���������|/��s�I"�gE�O�#[������T0 k� �����U2d  U8D"!  ��    ��� D� JD���������|/���I"�gE�W�#_������T0 k� �����U2d  U8D"!  ��    ��� EtKD���������|/���I"�gE�[�#c������T0 k� �����U2d  U8D"!  ��    ��� EtKD���������|/�Ç�I"�gE�c�#g�	�����T0 k� �����U2d  U8D"!  ��    ��� EtMD��������|/�Ó�@�gE�s�#o�	�����T0 k� �����U2d  U8D"!  �    ��� Et$NR��������|/�Û�@�gE�{�#s�	�����T0 k� �����U2d  U8D"!  ��    ��� Et(OR��������|/�ã�@�gE��#w�	�����T0 k� �����U2d  U8D"!   �    ��� Et0PR���������|/�ç�@�gEr��#{�	�����T0 k� �����U2d  U8D"!  �� 
   ��� Et<RR����$�����|/�÷�@�gEr��#��
�����T0 k� �����U2d  U8D"!  �� 
   ��� EtDSR����(�����|/�û�@�gEr��#��
�����T0 k� �����U2d  U8D"!  �� 
   ��� EtLUR����0���ǝ|/���@b�gEr��#��
�����T0 k� �����U2d  U8D"!  �� 
   ��� EdXWR����<���Ӛ|/���@b�gEr��#��
�����T0 k� �����U2d  U8D"!  �� 
   ��� Ed\XR����D���ۘ|/���@b�gEr��#��������T0 k� �����U2d  U8D"!  �� 
   ��� EddYR���L���ߗ|/���@b�gEr��#��������T0 k� �����U2d  U8D"!  �� 
   ��� Edp\R���X���|/���@b�gEr��#��������T0 k� �����U2d  U8D"!  �� 
   ��� Edt]R���\����|/���@��gEr��#��������T0 k� �����U2d  U8D"!  �� 
   ��� Edx^R���d����|/���@��gEr�� s��������T0 k� �����U2d  U8D"!  �� 
   ��� Ed�`R��sl���|/���@��gEr�� s��������T0 k� �����U2d  U8D"!  �� 
   ��� Ed|`R��st���|/���@��gEr�� s������T0 k� �����U2d  U8D"!  �� 
   ��� Edx`R��s�� ��|/���@��gEb�� s������T0 k� ������U2d  U8D"!  �� 
   ��� EdtaR��s�� ��|/���@��gEb���������T0 k� ������U2d  U8D"!  �� 
   ��� EdpaR��s��$ �'�|/���A�gEb���������T0 k� ������U2d  U8D"!  �� 
   ��� ETlbR��s��,!�3�|/���A�gEc����/����T0 k� ������U2d  U8D"!  �� 
   ��� EThbR��s��,"�;�|/���A�gEc����7����T0 k� ������U2d  U8D"!  �� 
   ��� ETdbR��s��0#�C�|/���A�gEc����?����T0 k� ������U2d  U8D"!  �� 
   ��� ET`bR��s��0#�K�|/���A�gEc����G����T0 k� ������U2d  U8D"!  �� 
   ��� C�XcR��s� �4$�W�|/���AR�gEc�����W����T0 k� ������U2d  U8D"!  �� 	   ��� C�TcR��c���4%�_�|/���AR�gEc�����_����T0 k� ������U2d  U8D"!  �� 	   ��� C�LcR��c���4&�c�|/��AR�gEc�����g����T0 k� ������U2d  U8D"!  �� 	   ��� C�DdR�#�c���8'�o�|/��AR�gES'�����w����T0 k� ������U2d  U8D"!  �� 	   ��� �C�@dR�#�c���8'�w�|/��C�gES+���������T0 k� ������U2d  U8D"!  �� 	   ��� �C�<dR�#�c���8'�{�|/���C�gES+����������T0 k� ������U2d  U8D"!  �� 	   ��� �C�0eR�'�c���8(���|/���C�gES/����������T0 k� ������U2d  U8D"!  �� 	   ��� �I�,eR�+�c���8(�|/���C�gES3���������T0 k� ������U2d  U8D"!  ��) 	   ��� �I�$eR�+�c���8(�|/���C�gES3���������T0 k� ������U2d  U8D"!  ��) 	   ��� �I�eR�/�c���4)�|/���C�gES7����t{����T0 k� ������U2d  U8D"!  ��) 	   ��� �I�fR�/�c��24)£�|/��#�C�gC�7����t{����T0 k� ������U2d  U8D"!  ��) 	   ��� �I�fR�/�3��24)§�|/��'�C�|gC�7����tw����T0 k� ������U2d  U8D"!  ��) 	   ��� �I�fR�/�3��24)«�|/��+�C�|gC�7����tw����T0 k� ������U2d  U8D"!  ��) 	   ��� �I�fR�3�3��20)¯�|/��/�C�xgC�4 ���ts����T0 k� ������U2d  U8D"!  ��) 	   ��� �I�fR�3�3��20)·�|/��7�C�pgC�4���ts����T0 k� ������U2d  U8D"!  ��) 	   ��� �I� fR�3�3��2,)»�|/��;�C�lgC�4���do����T0 k� ������U2d  U8D"!  ��) 	   ��� �I��fR�7�3��2,(¿�|/��C�C�dgC�4���do����T0 k� ������U2d  U8D"!  ��) 	   ��� �I��fR�7�3��2((�Ë|/��C�C�`gC�4���dk����T0 k� ������U2d  U8D"!  ��)    ��� �I��fR�7�3��2$(�ǌ|/��G�C�XgC�0���dk����T0 k� ������U2d  U8D"!  ��)    ��� �I��fR�;�#��2$'�ˍ|/��K�DPgC�0���dk����T0 k� ������U2d  U8D"!  ��)    ��� �I��fR�;�#��B '�ˍ|/��O�DLgES0	���dk����T0 k� ������U2d  U8D"!  ��)    ��� �I��fR�;�#��B '�ˎ|/��S�DHgES,
���dg����T0 k� ������U2d  U8D"!  ��)    ��� �I��fR�;�#��B&�ώ|/��W�D@gES,���Tg����T0 k� ������U2d  U8D"! $�)    ��� �I��fR�;�#��B&�Ϗ|/��W�D<gES(���Tc����T0 k� ������U2d  U8D"! ��/    ��� �I��fR�?�#��B&�Ϗ|/��[�D4gES(���Tc����T0 k� ������U2d  U8D"! ��/    ��� �I��fR�?�#��R%�Ϗ|/�t_�D0gES$���T_����T0 k� ������U2d  U8D"! ��/    ��� �I��fR�?�#��R%�Ӑ|/�tg�D$gES ����[�c��T0 k� #�����U2d  U8D"! ��/    ��� �I��fR�?�#��R$�ӑ|/�tk�DgEC����[�c��T0 k� #�����U2d  U8D"! ��/    ��� �I��fR�C�#��R$�ӑ|/�to�DgEC����W�c��T0 k� #�����U2d  U8D"!  ��/    ��� �I��fR�C�#��R #�Ӓ|/�ts�DgEC����S�c��T0 k� #�����U2d  U8D"!  ��/    ��� �I��fR�C�#�Q�#�ϒ|/�ts�DgEC����O�c��T0 k� #�����U2d  U8D"!  ��/    ��� �I��fR�C�#{���#�ϒ|/�tw�D gEC���TK�c��T0 k� ������U2d  U8D"!  ��/    ��� �I��fR�C�#w���#�ϓ|/�t{�D�gC����TG�c��T0 k� ������U2d  U8D"!  /�+    ��� �I��fR�C�#s���"�˓|/�d�D�gC����TC�s��T0 k� ������U2d  U8D"!  ��+    ��� �I��fR�G�#o���"�˔|/�d�EA�gC����TC�s��T0 k� ������U2d  U8D"!  ��+    ��� �I��fR�G�#g���"�˔|/�d��EA�gC����T;�s��T0 k� ������U2d  U8D"!  ��+    ��� �I��fR�G�#c���!�ǔ|/�d��EA�fC� ���T7�s��T0 k� ������U2d  U8D"!  ��+    ��� �I��fR�G�#_���!�Ǖ|/�d��EA�fC�����T3�s��T0 k� ������U2d  U8D"!  ��+    ��� �I��fR�G�#[���!�Õ!�/�d��EA�fC�����T/�s��T0 k� ������U2d  U8D"!  ��+    ��� �A�fR�G�#W��� �!�/�d��EA�fC�����T+�s��T0 k� ������U2d  U8D"!  ��+    ��� �A�fR�K�#S��� �!�/�d��EA�eC�����D'�s��T0 k� ������U2d  U8D"!  ��+    ��� �A�fR�K�#O��� �!�/�d��EA�eC�����D#�s��T0 k� ������U2d  U8D"!  ��+    ��� �A�fR�K�#K�� �!�/�T��EA�eC�����D�s��T0 k� ������U2d  U8D"!  ��+    ��� �A�fR�K�#G���!�/�T��C��dC�����D�s��T0 k� ������U2d  U8D"!  ��+    ��� �A�fR�K�c?���!�/�T��C��cC�������s��T0 k� ������U2d  U8D"!  ��+    ��� �A�fR�O�c;����!�/�T��C��cC����������T0 k� ������U2d  U8D"!  ��+    ��� �A�fR�O�c7����!�/�䓴C��bC����������T0 k� ������U2d  U8D"!  ��+    ��� �A�fR�O�c/����!�/�䓳Iq|bC�����������T0 k� ������U2d  U8D"!  ��+    ��� �A�fR�O�c+����|/�䓲IqtbC�����������T0 k� ������U2d  U8D"!  ��+    ��� �@��fR�O�S'����|/�䓱IqpbC����������T0 k� ������U2d  U8D"!  ��+    ��� �@��fR�O�S#����|/�䓰IqhaC����������T0 k� ������U2d  U8D"!  ��+    ��� �@��fR�O�S��|��|/�䏯IqdaC����������T0 k� ������U2d  U8D"!  ��+    ��� �@��fR�S�S��l��|/�䋭I�XaC������۠���T0 k� ������U2d  U8D"!  ��+    ��� �@��fR�S�S�d�|/�䇬I�PaC�� c���Ӡ���T0 k� ������U2d  U8D"!  ��+    ��� �@��fR�S�S�`{�|/�䇫I�LaC�� c���Ϡ���T0 k� ������U2d  U8D"!  ��+    ��� �@��fR�S�R��Xs�|/��I�HaC�� c���Ǡ���T0 k� ������U2d  U8D"!  ��+    ��� �@��fR�S�R��Po�|/���I�@aC�� c���à���T0 k� ������U2d  U8D"!  ��+    ��� �@��fR�S�B�Hg�|/��{�EA<`C�� c��C�����T0 k� ������U2d  U8D"!  ��+    ��� �@��fR�S�B�@c�!�/��w�EA4`C�� ��C�����T0 k� �����U2d  U8D"!  ��+    ��� �@��fR�W�B߱4W�!�/��s�EA(`C�� ��C��ӳ�T0 k� �{���U2d  U8D"!  ��+    ��� �A�fR�W�B۰,O�!�/��o�EA$_C ��C��ӫ�T0 k� �����U2d  U8D"!  ��+    ��� �A�fR�W�Bӯ$G�!�/��k�EA_C�| ��C��ӧ�T0 k� �����U2d  U8D"!  ��+    ��� �A�fR�W�B˯C�!�/��g�EA_C�xC��C��ӣ�T0 k� �����U2d  U8D"!  ��+    ��� �A�fR�W�BǮ;�!�/��c�EA^C�pC��3��ӟ�T0 k� �����U2d  U8D"!  ��+    ��� �A�fR�W�B��3�!�/��[�EA^C�lC��3�����T0 k� �s��w�U2d  U8D"!  ��+    ��� �AS�fR�W�B�� �'�!�/�S�E1 ]C�`C��3{����T0 k� �_��c�U2d  U8D"!  ��+    ��� �AS�fR�[�B�����!�/�O�E0�\C�X
C��3s����T0 k� �W��[�U2d  U8D"!  ��+    ��� �AS�fR�[�2�����|/�G�E0�[C�T
C��3o����T0 k� �K��O�U2d  U8D"!  ��+    ��� �AS�fR�[�2�����|/�C�E0�[C�L
C��3g�c�T0 k� �G��K�U2d  U8D"!  ��+    ��� �AS�fR�[�2�����|/�?�E0�ZC�D
C��3c�c{�T0 k� �C��G�U2d  U8D"!  ��+    ��� �C��fR�[�2������|/�7�E0�YC�@
C��3[�cw�T0 k� �;��?�U2d  U8D"!  ��+    ��� �C��fR�[�2������|/�3�E0�XC�8
s��CW�co�T0 k� �7��;�U2d  U8D"!  ��+    ��� �C��fR�[�B{����|/�'�E0�VC�,	
s��CK�cc�T0 k� �+��/�U2d  U8D"!  ��+    ��� �C��fR�[�Bs���ߠ|/��E0�UC�$
s��CC�c_�T0 k� �'��+�U2d  U8D"!  ��+    ��� �C��fR�_�Bo���Ӡ|/��E0�TC� 
s��C?�#[�T0 k� �+��/�U2d  U8D"!  ��+    ��� �C��fR�_�Bg���ˡ|/��E0�SC���C7�#S�T0 k� �/��3�U2d  U8D"!  ��+    ��� �C��fR�_�Bc���á|/��E �RC���C3�#O�T0 k� �/��3�U2d  U8D"!  ��+    ��� �C��fR�_�2W����|/���E �OC���C'�#C�T0 k� �+��/�U2d  U8D"!  ��+    ��� �C��fR�_�2O����|/���E �NC����C#��?�T0 k� �'��+�U2d  U8D"!  ��+    ��� �C��fR�_�2K����|/��E �MC����C��;�T0 k� �'��+�U2d  U8D"!  ��+    ��� �C��fR�_�2C����|/��E �LC�� ��C��3�T0 k� 3���U2d  U8D"!  �+    ��� �C�fR�_�2?��x�|/��E �JC���S��S��/�T0 k� 3���U2d  U8D"! ��/ 	   ��� �C�fR�_�27�	�p�|/�ۖE �IC���S��S��+�T0 k� 3���U2d  U8D"! ��/ 	   ��� C�fR�_�23�	�l�{�|/�ӖE �HC���S��S�S#�T0 k� 2����U2d  U8D"! ��/ 	   ��� {C�fR�c�2'�	�\�k�|/��ǕE �EC���S��S�S�T0 k� ������U2d  U8D"! ��/ 	   ��� wC�fR�c�2#�	�Xc�|/�㿔E �CC���S��R��S�T0 k� ������U2d  U8D"! ��/ 	   ��� sD�fUtc�2�	�P[�|/�㷔E�BC������R��S�T0 k� ������U2d  U8D"! ��/ 	   ��� oD�fUtc�2�	�LO�|/�㯓E�AC������R�c�T0 k� ������U2d  U8D"! ��/ 	   ��� kD�fUtc�2�	�HG�|/�㧓E�?C������R�c�T0 k� ������U2d  U8D"! ��/ 	   ��� gD�fUtc�2�	�@?�|/�㟒E�>C������R��c�T0 k� � �� U2d  U8D"! ��/ 	   ��� dD�fUtc�2�	�<7�|/�㗒E�<C������R��b��T0 k� ���U2d  U8D"!	 ��/ 	   ��� aEC�fUtc�2�	�8/�|/�㏑B��;C���3��b��b��T0 k� ���U2d  U8D"!
 ��/ 	   ��� ^EC�eUtc�1��	�4#�|/�㇑B��:C���3��b��b��T0 k� ���U2d  U8D"!
 ��/ 	   ��� [EC|eUtc�1��	�,�|/���B��9C���3��b��b��T0 k� ���U2d  U8D"! ��/ 	   ��� XECxeUtc�1��	�(�|/��w�B��7C���3��b��b��T0 k� B���U2d  U8D"! ��/ 	   ��� UECteA�c�1��	�$�|/��o�B��6C���3��b��b��T0 k� Bt�xU2d  U8D"! ��/ 	   ��� RECleA�c�1��	� �|/��g�B��5C���S��2��R��T0 k� Bl�pU2d  U8D"! ��/ 	   ��� OECheA�g�1��	� ��|/��_�B��4C�{�S��2��R��T0 k� B`�dU2d  U8D"! ��/ 	   ��� LEC`dA�g�1��	��|/��W�B��2C�w�S��2��R��T0 k� BT�XU2d  U8D"! ��/ 	   ��� IEC\dA�g�1��	��|/��O�B��1EAo�S��2��R��T0 k� "L�PU2d  U8D"! ��/ 	   ��� FECXdATg�1��	�ߥ|/��G�B��0EAg�S��2��R��T0 k� "@	�D	U2d  U8D"! ��/ 	   ��� CECPcATg�1��	�ӥ|/��?�B��/EAc�C��2��R��T0 k� "8
�<
U2d  U8D"! ��/ 
   ��� @E3LcATg�A��	�˦|/��7�B��.EA[�C��2��R��T0 k� ",�0U2d  U8D"! ��/ 
   ��� =E3DbATg�A��	�æ|/��/�B��-EAS�C��2��R��T0 k� " �$U2d  U8D"! ��/ 
   ��� :E3@bATg�A��	���|/��'�B��,EAO�C��2��R��T0 k� 2�U2d  U8D"! ��/ 
   ��� 7E38aAg�A��	���|/���B��+EAG�C��"��R��T0 k� 2�U2d  U8D"! ��/ 
   ��� 4E�,`Ag�1��	���|/���B��)EA;����"��R��T0 k� 1���U2d  U8D"! ��/ 
   ��� 1E�$`Ag�1��	����|/��B��(EA7����"��R��T0 k� 1���U2d  U8D"! ��/ 
   ��� .E� _Ag�1��	����|/���B��'EA/����"��R��T0 k� ����U2d  U8D"! ��/ 
   ��� +E�^C�g�1��	� ���|/���B��&E1'������R��T0 k� ����U2d  U8D"! ��/ 
   ��� (E�]C�g�1��	� �{�|/��B��%E1#������R��T0 k� ����U2d  U8D"! ��/ 
   ��� %E�]C�c�1��	� �s�|/��B��$E1������R��T0 k� ����U2d  U8D"! ��/ 
   ��� "C�\C�c�1��	� �k�|/�ۉB��#E1������R��T0 k� ����U2d  U8D"! ��/ 
   ��� C� [C�c�1��	� �c�|/�ӈB��"E1��������T0 k� ���U2d  U8D"! ��/    ��� C��ZC�c�1��	���[�|/�ˈB��!E1��������T0 k� ���U2d  U8D"! ��/    ��� C��ZC�_�1��	���O�|/�ÈB�� E1��������T0 k� ���U2d  U8D"! ��/    ��� C��YC�_�1��	���G�|/���B��E0���������T0 k� ���U2d  U8D"! ��/    ��� C��XC�[�1��	��@?�|/���B��E0���������T0 k� ���U2d  U8D"! ��/    ��� C��WC�[�1��	��@7�|/���B��E0��������� T0 k� A|��U2d  U8D"! ��/    ��� C��VC�[�1��	��@/�|/���B��E0��������T0 k� At�xU2d  U8D"! ��/    ��� 
C��UC�W�1��	��@#�|/���B��E ���{�����T0 k� Ah�lU2d  U8D"! ��/    ��� C��TC�S�1�	��@�|/���E�E ���w�����T0 k� A\�`U2d  U8D"! ��/    ��� C��SC�S�1���@�|/���E�E ���s�����T0 k� AT�XU2d  U8D"! ��/    ��� C��RC�O�1���@�|/���E�E ���k��� 2�
T0 k� !H�LU2d  U8D"! ��/    �����C��PC�K�1���O��|/�s�E�E ���c��� 2�T0 k� !4�8U2d  U8D"! ��/    �����C��OC�G�1���O�|/�k�E�E ���_��� 2�T0 k� !, �0 U2d  U8D"! ��/    �����C��NC�G�1|O���|/�c�E�E ���W��� 2�T0 k� !  �$ U2d  U8D"! ��/    �����C��LC�C�1xO��߫|/�[�E E ���S��� B�T0 k� �!�!U2d  U8D"! ��/    �����C��KC�?�1tO��׬|/��S�EE ���O��  B�T0 k� �"�"U2d  U8D"! ��/    �����C��JC�;�1tO��ˬ|/��K�EE ÿ�G�� B�T0 k� � #�#U2d  U8D"! ��/    �����C��IC�7�1pO��í|/��C�EE���C�� B�T0 k� ��$��$U2d  U8D"! ��/    �����C�xHC�3�1p ����|/��;�E�E��C?�� B�T0 k� ��$��$U2d  U8D"! ��/    �����C�pFC�/�1l ����|/��3�E�$E��C7�� B�T0 k� ��%��%U2d  U8D"! ��/    �����C�hEE�+��h ����|/��+�E�(E��C3��	 B�T0 k� ��&��&U2d  U8D"! ��/    �����C�dDE�'��h! ����|/��#�E�0E��C+��
 B�T0 k�  �'��'U2d  U8D"! ��/    �����C�\CE�#��d# ����|/���E�8E��C'�� B�T0 k�  �(��(U2d  U8D"!
 ��/    �����C�TAE���`%�����|/���E�@E��C#�� R�T0 k�  �)��)U2d  U8D"!
 ��/    �����C�L@E���`'�����|/���E�HE��C�� R�T0 k�  �)��)U2d  U8D"!	 ��/    �����C�D?E���\)� ��|/���E�LE��3�� S T0 k�  �*��*U2d  U8D"! ��/    �����E�<>C���\+� �w�|/����E�TE��3�"� ST0 k� �+��+U2d  U8D"! ��/    �  ��E�8<C���X-� �o�|/���E�\E��3�"� ST0 k� �,��,U2d  U8D"! ��/    � ��E�0;C���T/� �g�|/���E�dE���3�"� ST0 k� ��-��-U2d  U8D"! ��/    � ��E�(:C���P1� �_�|/���EqlE���2��"� ST0 k� �|.��.U2d  U8D"! ��/    � ��E� 9C����P3��W�|/��ۀEqtE���	R��"� ST0 k� �p.�t.U2d  U8D"! ��/    � ��E�7C����L5��O�|/��ӁEq|E���	R��"� $T0 k� �h/�l/U2d  U8D"! ��/    � ��E�6C���H7��C�|/��ˁEq�E���	R��"� (T0 k� �\0�`0U2d  U8D"! ��/    � ��E�5C���D9��;�|/��ÁEq�E���	R��"� 0T0 k�  P1�T1U2d  U8D"! ��/    � ��E�4C���@;��3�|/��Eq�E���	R��"�! 4T0 k�  H2�L2U2d  U8D"! ��/    � ��E��2C�߸�@= �+�|/��Eq�E���	b��"�# <T0 k�  <2�@2U2d  U8D"!  ��/    � ��E��1C�׷�<? �#�|/��Eq�E���	b��"�% #@T0 k�  0/�4/U2d  U8D"!  ,�3    � ��E��0C�ӷ�8@ ��|/��Eq�Ep��	b��"�' #HT0 k�  ,-�0-U2d  U8D"!  �3    � ��E��/AS˶�4B ��|/�Q��Eq�Ep��	b����) #LT0 k� �,+�0+U2d  U8D"!  �3    � ��E��-ASǶ�0D ��|/�Q��Ea�Ep��	b����+ #TT0 k� �,+�0+U2d  U8D"! ��3    � ��E��,AS��Q,F���|/�Q��Ea�Ep�������, #XT0 k� �0+�4+U2d  U8D"! ��3    � ��E��+AS��Q(H���|/�Q�Ea�Ep�������.�\T0 k� �0+�4+U2d  U8D"! ��3    � ��E��*AS��Q$I��|/�Qw�Ea�Ep�������0�dT0 k� �4+�8+U2d  U8D"! ��3    � ��E��)AS��Q K��|/�Qo�Ea�E`�������2�hT0 k� �4+�8+U2d  U8D"! ��3    � ��AQ�(AS��QM���|/�Qg�Ea�E`�������4�lT0 k� �4,�8,U2d  U8D"! ��3    � ��AQ�'AS��QN���|/�Q_�Ea�E`��¿���6�pT0 k�  4,�8,U2d  U8D"! ��3    � ��AQ�&AS��QP���|/�QW�Ea�E`��»���7�xT0 k�  8,�<,U2d  U8D"! ��3    � ��AQ�%AS��QQ���|/�AO�Ea�E`��ҷ���9�|T0 k�  8,�<,U2d  U8D"! ��3    � ��AQ�$AS��QS���|/�AG�Ea�D0��Ұ ��;��T0 k�  8,�<,U2d  U8D"! ��3   � ��AQ�#AS��QT `��|/�A?�Ea�D0��Ҩ��=��T0 k�  8-�<-U2d  U8D"! ��3    � ��AQ�"AS��QV `��|/�A7�EQ�D0��Ҥ��?��T0 k� �8-�<-U2d  U8D"! ��3    � ��AQ�!AS��QW ` ��|/�A/�EQ�D0��Ҡ��A��T0 k� �8-�<-U2d  U8D"! ��3    � ��AQ� AS�Q Y ` ��|/��'�EQ�D0�����C��T0 k� �<-�@-U2d  U8D"! ��3    � ��AQ�ASw�Q Z ` ��|/���EQ�D0�����D��T0 k� �<.�@.U2d  U8D"! ��3    � ��AQ�ASs�P�\  ��|/���EQ�D0�����F��T0 k� �0/�4/U2d  U8D"! ��3    � ��AQ|ASo�P�]   ��|/���EQ�D0�����H��T0 k� �(0�,0U2d  U8D"! ��3    � ��AQtASk�P�^   ��|/���EQ�D@�����J��T0 k� �$0�(0U2d  U8D"! ��3    � ��AQpASg�P�` $ ��|/����C��D@�����L��T0 k�   1�$1U2d  U8D"! ��3    � ��AQlAS_�P�a $!��|/����C��D@���x��N��T0 k�  ,0�00U2d  U8D"! �3    � ��AQdAS[�P�b�$!��|/���C��D@���t��P��T0 k�  4/�8/U2d  U8D"! ��?    � ��AQ`ASW�P�d�$!�|/���C�� D@���l	��R��T0 k�  @/�D/U2d  U8D"! ��?    � ��AQ\ASS�P�e�$!w�|/��ߊC�� D@���d
��T��T0 k�  H.�L.U2d  U8D"!
 ��?    � ��AQTASO�P�f�$"s�|/��׋C��!D@���`��V��T0 k� �T-�X-U2d  U8D"! ��?    � ��AQPASK�P�g�("k�|/��ϋC��"D@���X��W��T0 k� �\,�`,U2d  U8D"! ��?    � ��AQLASG�P�i�("g�|/��ǌC��"D@���T� Y��T0 k� �h,�l,U2d  U8D"! ��?    � ��AQHASC�P�j�("c�|/�@��C��#D@���L� [��T0 k� �p+�t+U2d  U8D"! ��?    � ��AQDAS?�P�k�("[�|/�@��C��#D@���D� ]��T0 k� �|*��*U2d  U8D"! ��?    � ��AQ@AS;�P�l�(#W�|/�@��C��$DP���<� _��T0 k� ��*��*U2d  U8D"! ��?    � ��AQ8AS7�P�m�(#S�|/�@��C��%DP���4�a��T0 k� ��)��)U2d  U8D"! ��?    � ��AQ4AS3�P�n�(#O�|/�@��C��%DP���0�c��T0 k�  �(��(U2d  U8D"! ��?    � ��AQ0AS/�P�p�,#G�|/�@��C��&DP���(�e��
T0 k�  �(��(U2d  U8D"! ��?    � ��AQ,AS+�P�q�,$C�|/�@��C��&DP�� �g��
T0 k�  �'��'U2d  U8D"! ��?    � ��AQ(AS'�P�r�,$?�|/�0��C��'DP���i��
T0 k�  �&��&U2d  U8D"! ��?    � ��AQ$AS#�P�s�,$;�|/�0��C��(DP���k��	T0 k�  �%��%U2d  U8D"! ��?    � ��AQ AS�P�t�,$7�|/�0{�EQ�(DP���l��	T0 k� ��%��%U2d  U8D"! ��?    � ��AQAS�P�u�,$3�|/�0s�EQ�)DP�� � n��	T0 k� ��$��$U2d  U8D"! ��?    � ��AQAS�P�v�,%+�|/�0k�EQ�)DP���� p��T0 k� ��#��#U2d  U8D"! ��?    � ��AQAS�P�w�,%'�|/�0c�EQ�*DP��� r��T0 k� ��#��#U2d  U8D"! ��?    � ��AQAS�P�x�0%#�|/�0_�EQ�*D`{��� s��T0 k� ��"��"U2d  U8D"! ��?    � ��AQAS�P�y�0%�|/�0W�E��*D`w����u��T0 k� ��!� !U2d  U8D"!  ��?    � ��AQAS�P�z �0%�|/�0O�E��+D`s����w��T0 k� �!�!U2d  U8D"!! ��?    � ��AQ
AS�P�{ �0&�|/�0K�E��+D`s����x��T0 k� ! � U2d  U8D"!" ��?    � ��AQ 	AS�P�{ �0&�|/�@C�E��,D`o����z� T0 k� !� U2d  U8D"!# ��?    � ��AP�	AS�P�| �0&�|/�@;�E��,D`k����{� T0 k� !$�(U2d  U8D"!$ ��?    � ��AP�AR��P�} �0&�|/�@7�E��-D`g����}�T0 k� !0�4U2d  U8D"!$ ��?    � ��AP�AR��P�~ �0&�|/�@/�E��-D`c���~�T0 k� !8�<U2d  U8D"!% ��?    � ��AP�AR��P� �0&�|/�@+�EѼ-L0[����T0 k� �D�HU2d  U8D"!& ��?    � ��AP�AR��P�� �4'��|/�@#�C�.L0W����T0 k� �L�PU2d  U8D"!' ��?    � ��AP�AR�P�� �4'��|/�@�C�.L0S����T0 k� �X�\U2d  U8D"!( ��?    � ��AP�AR�P� �4'��|/�@�C�/L0S����T0 k� �`�dU2d  U8D"!( ��?    � ��AP�AR�P� �4'��|/�@�C�/L0O���~�T0 k� �l�pU2d  U8D"!) ��?    � ��AP�AR�P� �4'��|/�@�C�/L0K�x�~�T0 k� �t�xU2d  U8D"!* ��?    � ��AP�AR�P� �4'��|/�@�C�0L0G�Qp�~�T0 k� ����U2d  U8D"!+ ��?    � ��AP�AR�P�~ �4'��|/�@�C�0L0C�Qh�}� T0 k� !���U2d  U8D"!+ ��?    � ��AP�AR�P�~ �4(��|/�_��C�1L0?�Q`�}� T0 k� !���U2d  U8D"!, ��?    � ��AP�ARߠP�~ �4(��|/�_��C�1L0;�QX�}� T0 k� !���U2d  U8D"!, ��?   � ��AP�ARߠP�~ �4(��|/�_�C�1L07�QP�|� T0 k� !���U2d  U8D"!- ��?    � ��AP�AR۟P�} �8(��|/�_�C�|2L03�QH�|� T0 k� !���U2d  U8D"!- ��?    � ��AP�AR۟P�} �8(��|/�_�C�t2L0/�Q@�|� T0 k� ���U2d  U8D"!. ��?    � ��AP�ARןP�} �8(��|/�_�C�p2L0/�Q8"�{� T0 k� ����U2d  U8D"!. ��?    � ��AP� ARӟP�} �8(��|/�_ߵC�h3L@+�Q0"�{��T0 k� ����U2d  U8D"!/ ��?    � ��AP� ARӟP�} �8)��|/�_׷C�`3L@'�Q("�{��	T0 k� ����U2d  U8D"!/ ��?    � ��AP��ARϞP�| �8)��|/�_ӸC�X3L@#�Q "�{��	T0 k� ����U2d  U8D"!0 ��?    � ��AP��ARϞP�| �8)��|/�_ϺC�T4L@�Q"�z��	T0 k� ����U2d  U8D"!0 ��?    � ��AP��AR˞P�| �8)��|/�_˼C�L4L@�Q"�z��	T0 k� ����U2d  U8D"!0 ��?    � ��AP��AR˞P�| �8)��|/�oǽC�D4L@�Q "�z��	T0 k� " �U2d  U8D"!1 ��?    � ��AP��ARǝP�| �8)��|/�oÿC�<5L@�Q "�z��	T0 k� "�U2d  U8D"!1 ��?    � ��AP��ARǝP�{ �8)��|/�o��C�45L@�P� "�y��
T0 k� "�U2d  U8D"!1 ��?    � ��AP��ARÝP�{ �8*��|/�o��C�,5L@�P�!"�y��
T0 k� "� U2d  U8D"!2 ��?    � ��AP��ARÝP�{ �<*��|/�o��C�$5L@��!"�y��
T0 k� "(�,U2d  U8D"!2 ��?   � ��AP��AR��P�{ �<*��|/�o��D6L@��!"�x��
T0 k� �0�4U2d  U8D"!2 ��?    � ��AP��AR��P�{ �<*��|/�o��D6L@��""�x��
T0 k� �<�@U2d  U8D"!2 ��?    � ��AP��AR��P�z �<*��|/�o��D6L@��""�x��
T0 k� �D
�H
U2d  U8D"!2 ��?    � ��AP��AR��P�z �<*��|/�o��D7L@��""�x��
T0 k� �P	�T	U2d  U8D"!2 ��?    � ��AP��AR��P�z �<*��|/�o��D �7L@��#"�x��T0 k� �X	�\	U2d  U8D"!3 ��?    � ��AP��AR��P�z �<*��|/�o��D �7LO���#"�w��T0 k� �d�hU2d  U8D"!3 ��?    � ��AP��AR��P�z �<*��|/���D �7LO���#"�w��T0 k� �l�pU2d  U8D"!3 ��?    � ��AP��AR��P�z �<+��|/���D �8LO���$"�w��T0 k� "x�|U2d  U8D"!3 ��?    � ��AP��AR��P�y �<+��|/���D �8LO���$"�w��T0 k� "���U2d  U8D"!3 ��?    � ��AP��AR��P�y �<+��|/���D �8LO���$"�v��T0 k� "���U2d  U8D"!3 ��?    � ��AP��AR��P�y �<+��|/���D �8LO���$"�v��T0 k� "���U2d  U8D"!2 ��?    � ��AP��AR��P�y �<+��|/�߇�D�9LO���%"�v��T0 k� "���U2d  U8D"!2 ��?    � ��AP��AR��P�y �<+��|/�߃�D�9LO���%"�v��T0 k� ���U2d  U8D"!2 ��?    � ��AP��AR��P|y �@+��|/���D�9LO�� �%"�v��T0 k� ���U2d  U8D"!2 ��?    � ��AP��AR��P|y �@+��|/��{�D�9LO�� �%"�u��T0 k� ���U2d  U8D"!2 ��?    � ��AP��AR��P|x �@+��|/��{�D�9LO�� �&"�u��T0 k� ����U2d  U8D"!2 ��?    � ��AP��AR��P|x �@+��|/��w�D�:LO�� �&"�u��T0 k� �� �� U2d  U8D"!1 ��?    � ��AP��AR��Pxx �@,��|/��s�D�:LO�� �&"�u��T0 k� �� �� U2d  U8D"!1 ��?    � ��AP��AR��Pxx �@,��|/��o�D|:LO�� �'"�u��T0 k� ������U2d  U8D"!1 ��?    � ��AP��AR��Pxx �@,��|/��k�Dp:LO�� �'"�t��T0 k� "�����U2d  U8D"!1 ��?    � ��AP��AR��Pxx �@,��!�/��k�Dh;LO�� �'"�t��T0 k� "�����U2d  U8D"!0 ��?    � ��AP��AR��Pxx �<,��!�/��g�D`;LO�� |'"�t��T0 k� #���U2d  U8D"!0 ��?    � ��AP��AR��Ptw �<,��!�/��c�C�T;LO�� |'"�t��T0 k� #���U2d  U8D"!0 ��?    � ��AP��AR��Ptw �<,��!�/��_�C�L<LO�� x'"�t��T0 k� #���U2d  U8D"!/ ��?    � ��AP��AR��Ptw �<,��!�/��_�C�D<LO�� x'"�t��T0 k� �#��'�U2d  U8D"!/ ��?    � ��AP��AR��Ptw �8+��!�/��[�C�<=LO�� t'"�s��T0 k� �/��3�U2d  U8D"!. ��?    � ��AP��AR��Ptw �4+��!�/��W�C�4=LO�� p'"�s��T0 k� �7��;�U2d  U8D"!. ��?    � ��AP�AR��Ppw �0+�!�/��W�E�,>LO�� p'"�s��T0 k� �C��G�U2d  U8D"!- ��?    � ��AP�AR��Ppw �0+�!�/��S�E� >LO�� l'"�s��T0 k� �K��O�U2d  U8D"!- ��?    � ��AP�AR��Ppw �,+�!�/��O�E�?LO�� l'"�s��T0 k� �W��[�U2d  U8D"!, ��?    � ��AP{�AR��Ppw �(+{�!�/��O�E�?LO�� h'�s��T0 k� �_��c�U2d  U8D"!+ ��?    � ��AP{�AR��Ppv �(+{�|/��K�E�@L?�� h(�r��T0 k� #k��o�U2d  U8D"!+ ��?    � ��AP{�AR��Plv �$+w�|/��G�E��@L?�� d(�r��T0 k� #s��w�U2d  U8D"!* ��?    � ��APw�AR��Plv � +w�|/��G�E��AL?�� d(�r��T0 k� #����U2d  U8D"!* ��?    � ��APw�AR��Plv � +w�|/��C�E��AL?�� `(�r��T0 k� #�����U2d  U8D"!) ��?    � ��APw�AR��Plv �*s�|/��C�E��BL?�� `(�r��T0 k� #�����U2d  U8D"!( ��?    � ��APs�AR��Plv �*s�|/��?�E��CL?�� \(�r��T0 k� �����U2d  U8D"!' ��?    � ��APs�AR��Phv �*o�|/��;�E��CE��� \(�r��T0 k� �����U2d  U8D"!' ��?    � ��APs�AR��Phv �*o�|/��8 E��DE��� X(�q��T0 k� �����U2d  U8D"!& ��?    � ��APo�AR��Phv �*o�|/��4E��EE��� X(�q��T0 k� �����U2d  U8D"!% ��?    � ��APo�AR��Phv �*k�|/��4E�EE��� X(�q��T0 k� ������U2d  U8D"!$ ��?    � ��APo�AR��Phu �*k�|/��0E�FE��� T(�q��T0 k� ������U2d  U8D"!# ��?    � ��APo�AR��Phu �*k�!�/��0E�GE��� T(�q��T0 k� ������U2d  U8D"!" ��?    � ��APk�AR��Phu �*g�!�/��,D?�GE��� P(�q��T0 k� #�����U2d  U8D"!! ��?    � ��APk�AR�Pdu �*g�!�/��,D?�HE��� P(�|q��T0 k� #�����U2d  U8D"!  ��?    � ��APk�AR�Pdu �*g�!�/��(D?�IE��� L(�|q��T0 k� #�����U2d  U8D"! ��?    � ��APg�AR�Pdu �*g�!�/��(	D?�JE��� L(�xp��T0 k� #����U2d  U8D"! ��?    � ��APg�AR�Pdu � )c�!�/��$
D?xJD��� L(�tp��T0 k� $���U2d  U8D"! ��?    � ��APg�AR{�Pdu � )c�!�/��$I�pKD��� H(�pp��T0 k� ����U2d  U8D"! ��?    � ��APg�AR{�Pdu ��)c�!�/�� I�hLD��� H(�lp��T0 k� ����U2d  U8D"! ��?    � ��APc�AR{�Pdu ��)_�!�/�� I�`LD��� H(�hp��T0 k� �'��+�U2d  U8D"! ��?    � ��APc�AR{�P`u ��)_�!�/��I�XMD��� D(�dp��T0 k� �/��3�U2d  U8D"! ��?    � ��APc�ARw�P`u ��)_�!�/��I�TMD��� D(�`p��T0 k� �;��?�U2d  U8D"! ��?    � ��APc�ARw�P`t ��)[�|/��I�LND��� @(�\p��T0 k� �C��G�U2d  U8D"! ��?   � ��AP_�ARw�P`t ��)[�|/��I�DND���@(�Xp��T0 k� �O��S�U2d  U8D"! ��?    � ��AP_�ARw�P`t ��)[�|/��I�@OD���@)�Tp��T0 k� $W��[�U2d  U8D"! ��?    � ��AP_�ARw�P`t ��)[�|/��I�8OD���<)�Po��T0 k� $c��g�U2d  U8D"! ��?    � ��AP_�ARs�P`t ��)W�|/��I�4OD���<)�Lo��T0 k� $k��o�U2d  U8D"! ��?    � ��AP[�ARs�P`t ��)W�|/��I�,OD���<)�Do��T0 k� $w��{�U2d  U8D"! ��?    � ��AP[�ARs�P\t ��)W�|/��I�(PD���8)@o��T0 k� $����U2d  U8D"! ��?    � ��AP[�ARs�P\t ��)W�|/��I�$PD���P8)<o��T0 k� �����U2d  U8D"! ��?    � ��AP[�ARs�P\t ��)S�|/��I� PD���P8)4o��T0 k� ������U2d  U8D"! ��?    � ��AP[�ARo�P\t ��)S�|/��I�PD���P8)0o��T0 k� ������U2d  U8D"!
 )�?    � ��APW�ARo�P\t ��(S�|/��I�PD���P4),o��T0 k� ������U2d  U8D"!
 ��?    � ��APW�ARo�P\t ��(S�|/��I�PD���P4)$o��T0 k� ������U2d  U8D"!	 ��?    � ��APW�ARo�P\t ��(O�|/��I�PD���P4) o��T0 k� �����U2d  U8D"!	 ��?    � ��APW�ARo�P\t ��(O�|/��I�PD���P0)o��T0 k� �����U2d  U8D"! ��?    � ��APW�ARo�P\t ��(O�|/��I�PD���P0)n��T0 k� �����U2d  U8D"! ��?    � ��APS�ARk�PXt ��(O�|/�� I�PD���P0)n��T0 k� �����U2d  U8D"! ��?    � ��APS�ARk�PXs ��(O�|/�� I� PD���P,)n��T0 k� �����U2d  U8D"! ��?    � ��APS�ARk�PXs ��(K�|/�O I��PD���P,) n��T0 k� ԋ����U2d  U8D"! ��?    � ��APS�ARk�PXs ��(K�|/�N�I��PD���P,)�n��T0 k� ԇ����U2d  U8D"! ��?    � ��APS�ARk�PXs ��(K�|/�N�I��PD���P,)�n��T0 k� ԇ����U2d  U8D"! ��?    � ��APO�ARg�PXs ��(K�|/�N� I��PD���P()�n��T0 k� �����U2d  U8D"! ��?    � ��APO�ARg�PXs ��(G�|/�N�!I��PD���P()�n��T0 k� ����U2d  U8D"! ��?    � ��APO�ARg�PXs ��(G�|/�N�"I��PD���P()�n��T0 k� {���U2d  U8D"!  ��?   � ��APO�ARg�PXs ��(G�|/�N�#I��PD���P$)�n��T0 k� w��{�U2d  U8D"!  ,�?    � ��APO�ARg�PXs ��(G�|/�N�$I��PD���P$)�n��T0 k� w��{�U2d  U8D"!  ��?    � ��APK�ARg�PTs ��(G�|/�N�%I��PD��P$)�n��T0 k� s��w�U2d  U8D"!  ��?    � ��APK�ARg�PTs ��(C�|/�N�&I��PD��P$)�m��T0 k� �s��w�U2d  U8D"! ��?    � ��APK�ARc�PTs ��(C�|/�N�(I��PD��P )�m��T0 k� �o��s�U2d  U8D"! ��?    � ��APK�ARc�PTs ��(C�|/�^�)I��PD��P )�m��T0 k� �k��o�U2d  U8D"! ��?    � ��APK�ARc�PTs ��(C�|/�^�*I��PD��P )�m��T0 k� �k��o�U2d  U8D"! ��?    � ��APK�ARc�PTs ��(C�|/�^�+I��PD��
P )�m��T0 k� �g��k�U2d  U8D"! ��?    � ��APG�ARc�PTs ��'C�|/�^�-I��PD��P )�m��T0 k� �g��k�U2d  U8D"! ��?    � ��APG�ARc�PTs ��'?�|/�^�.I��PEo�P)�m��T0 k� �c��g�U2d  U8D"! ��?    � ��APG�ARc�PTs ��'?�|/�^�0I��PEo�P)�m��T0 k� �_��c�U2d  U8D"! ��?    � ��APG�ARc�PTs ��'?�|/�^�1I��PEo�P)!�m��T0 k� �_��c�U2d  U8D"! ��?    � ��APG�AR_�PTs ��'?�|/�^�2L>�PEo�P*!�m��T0 k� �[��_�U2d  U8D"! ��?    � ��APG�AR_�PTs ��'?�|/�^�4L>�PEo�P*!�m��T0 k� �W��[�U2d  U8D"! ��?    � ��APG�AR_�PTr ��'?�|/�^�5L>�PEo�P*!�m��T0 k� �W��[�U2d  U8D"! ��?   � ��APC�AR_�PPr ��';�|/�^�7L>�PEo�P*!|m��T0 k� �S��W�U2d  U8D"! ��?    � ��APC�AR_�PPr ��';�|/�n�9L>�PEo|P*!xm��T0 k� �S��W�U2d  U8D"! ��?    � ��APC�AR_�PPr ��';�|/�n�:L>�PEo|P*!pm��T0 k� �O��S�U2d  U8D"! ��?    � ��APC�AR_�PPr ��';�|/�n�<L>�PD?x P*!lm��T0 k� �K��O�U2d  U8D"! ��?    � ��APC�AR_�PPr ��';�|/�n�>L>�PD?x!P*!hm��T0 k� �K��O�U2d  U8D"! ��?    � ��APC�AR_�PPr ��';�|/�n�?L>�PD?x#P*!dm��T0 k� �G��K�U2d  U8D"! ��?    � ��APC�AR[�PPr ��';�|/�	^�?L>�QD?t%P*!`l��T0 k� �C��G�U2d  U8D"! ��?   � ��APC�AR[�PPr ��';�|/�	^�?L>�QD?p'P*!Xl��T0 k� �C��G�U2d  U8D"! ��?    � ��AP?�AR[�PPr ��'7�|/�	^�@LN�RD?p)P*!Tl��T0 k� �?��C�U2d  U8D"! ��?    � ��AP?�AR[�PPr ��'7�|/�	^�@LN�RD?l+P*!Pl��T0 k� �?��C�U2d  U8D"! ��?    � ��AP?�AR[�PPr ��'7�|/�	^�ALN�SD?l-P*!Ll��T0 k� �;��?�U2d  U8D"! ��?    � ��AP?�AR[�PPr ��'7�|/�	n�ALN�TD?h/P*!Hl��T0 k� �7��;�U2d  U8D"! ��?   � ��AP?�AR[�PPr ��'7�|/�	n�BLN�TD?h1P*!Dl��T0 k� �7��;�U2d  U8D"! ��?    � ��AP?�AR[�PPr ��'7�|/�	n�BLN�UD?d3P*!@l��T0 k� 3��7�U2d  U8D"! ��?    � ��AP?�AR[�PPr ��'7�|/�	n�BLN�UD?`4P*!<l��T0 k� 3��7�U2d  U8D"! ��?    � ��AP?�AR[�PPr ��'7�|/�	n�CLN�VDO`6P*!8l��T0 k� /��3�U2d  U8D"! ��?   � ��AP?�AR[�PPr ��'3�|/�	^�CLN�VDO\8P*!4l��T0 k� +��/�U2d  U8D"!  ��?    � ��AP?�ARW�PLr ��'3�|/�	^�CLN�WDOX:P*!0l��T0 k� +��/�U2d  U8D"!  ��?    � ��AP;�ARW�PLr ��'3�|/�	^�CLN�WDOX<P*!,l��T0 k� �'��+�U2d  U8D"!  ��?    � ��AP;�ARW�PLr ��'3�|/�	^�DLN�XDOT>P*!(l"��T0 k� �#��'�U2d  U8D"!  .�?    � ��AP;�ARW�PLr ��'3�|/�	^�DLN�XEoP@P*!$l"��T0 k� �#��'�U2d  U8D"!  ��?    � ��AP;�ARW�PLr ��'3�|/�N�ELN�YEoLAP*! l"��T0 k� ���#�U2d  U8D"!  ��?    � ��AP;�ARW�PLr ��'3�|/�N�ELN�YEoLCP*!l"��T0 k� ���#�U2d  U8D"!  ��?    � ��AP;�ARW�PLr ��'3�|/�N�FLN�ZEoHEP*!l"��T0 k� ���U2d  U8D"!  ��?    � ��AP;�ARW�PLr ��'3�|/�N�FLN�ZEoDGP*!l"��T0 k� ���U2d  U8D"!  ��?    � ��AP;�ARW�PLr ��'/�|/�N�GLN�[Eo@IP*!l"��T0 k� ���U2d  U8D"!  ��?    � ��AP;�ARW�PLr ��'/�|/�N�HLN�[Eo@KP*!l"��T0 k� ���U2d  U8D"!  ��?    � ��AP;�ARW�PLr ��'/�|/�N�ILN�\E_<LP*!l"��T0 k� ���U2d  U8D"!  ��?    � ��AP;�ARW�PLr ��'/�|/�N�ILN�\E_8NP*!l"��T0 k� ����U2d  U8D"!  ��?   � ��AP7�ARW�PLr ��'/�|/�^�JLN�]E_4PP*!l"��T0 k� ����U2d  U8D"!  ��?    � ��AP7�ARS�PLr ��'/�|/�^�KLN�]E_0RP*!l��T0 k� ����U2d  U8D"!  ��?    � ��AP7�ARS�PLr ��&/�|/�^�KLN�]E_,SP*! l��T0 k� ����U2d  U8D"!  ��?    � ��AP7�ARS�PLr ��&/�|/�^�LLN�^E_(UP* �k��T0 k� ����U2d  U8D"!  ��?    � ��AP7�ARS�PLr ��&/�|/�^�LLN�^E_$VP* �k��T0 k� ����U2d  U8D"!  ��?    � ��AP7�ARS�PLr ��&/�|/�^�MLN�_E_ XP* �k��T0 k� �����U2d  U8D"!  ��?    � ��AP7�ARS�PLq ��&/�|/�^�MLN�_E_ZP* �k��T0 k� �����U2d  U8D"!  ��?    � ��AP7�ARS�PLq ��&+�|/�^�NLN�_E_ZP* �k��T0 k� ������U2d  U8D"!  ��?    � ��AP7�ARS�PLq ��&+�|/�^�NLN�`E_\P*�k��T0 k� ������U2d  U8D"!  ��?    � ��AP7�ARS�PLq ��&+�|/�^�NLN�aE_]P*�k��T0 k� ������U2d  U8D"!  ��?    � ��AP7�ARS�PLq ��&+�|/�^�OLN�aL^P*�k��T0 k� �����U2d  U8D"!  ��?    � ��AP7�ARS�PLq ��&+�|/�n�OLN�bL_P*�k��T0 k� �����U2d  U8D"!  ��?    � ��                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��p ]�'�'� � ����2d       � 
��    ��5� 
��    ����               
   �          ��     ���   8	          ���w  ,      � �c�    ���� �h)    ����              A��          ��     ���   0	%           y��            "s     yv�  ��    �e   
         
  ; 7         �  �  ���   0
 	          &z�          ��>�     &z���K�      �?              	 ��$          \�  �  ���   8         ���         .�Hl    ���H2     X��                �$          �0     ���   P	         ��r2  ��     B�6i    ��r2�6i                           
  ���s              g  ���    P              O�k  � �
	   V��6�     O�k��6�                    	 Z��         �`�  '  ��`  (

          g4 0 0  
  j��j     g������    ��H           ( Z��          ���  	  ��@  8�           {<� � � 
	   ~���8     {j���X    �R��           O Z��         � �    ��` 	@


           +:1  � �
	   ����\     +:1���u      �w              . Z��         	 ��    ��h   H	$
          e  > >  	   ����     e'?����    ���               Z��         
 @�     ��@   H

!          `E ��     � �@�     ]& �@�     /                       ��V             �  ��@    0                ��      �                                                                           �                               ��        ���          ��                                                                 �                         ���  ��        � ��    ���o ݗ!    �m�: "                 x                j  �   �   �                         ��    ��       � �      ��   �           "                                                  �                          
 �  ���H����������� ��� � � 
  	              
   �  
,� ��A        �m@ �$ �j� �$ k� �D k� �d l  Є l  Ф l@ �d q@ �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À���� � � }`���� � .� s@ .�  s` � �h@ � 0i@ �d  i� פ i� �� �j� ¤ 0k� � l  �$ l@ � �^@ � _@ ބ �c@ �$ �m@ �$ n@ �D n` �d n� Є n� Ф n� �� t� �� �t� �� u� ބ �[�  � �e� � f� ބ �o����� � 
�< U� 
� V  
�\ V  
�\ V� 
�� V� 
�| W                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �������� �� D  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    "�j�� , " �
� �  �  
�  !��  ��     � 	  �    &��  ��     ���       +    ��     ���          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �?$      ��5 �  ���        � �  ���        �        ��        �        ��        �    ��    ���� ��        ��                         �w� $ �� ����                                     �                ����              	���%��   ����                15 Kevin Todd rson y   4:32                                                                        4  4     �LC. �dC6 � �kjS �k~g � k�o �cV= � c^E � c_5 � 	c`5 � 
ca@ � cb; �C � C"+ � c�e �c� � c�* � c� � c� � c� y c� �Ci � Cq �J� � � J� � �"� � "�  �"� �*� �"� � "�) �� � 
�" �!"� � ""�) �#� � 
�" � 
�" � 
�! ~'
� q ("J �I  "J q �*!� y/  "  y � ,"�1 �-� �.
�& �  "P � �  "P � �1
�% p2"8 � �  "P � �  "P � �  "P �  6"J �8 !� |@ !� |@ !� |(  "P �(  "P �X <*CT` =*G\`  *K<,  *F�                                                                                                                                                                                                                         �� R @       �     @ 
        �     a P E c  ���� Z   	           	 �������������������������������������� ���������	�
��������                                                                                          ��    �MJ�� ��������������������������������������������������������   �4, ?  * =�� t� @��@���	��ς	������                                                                                                                                                                                                                                                                                                                                �                                                                                                                                                                                                                                             
      \    (    ��  D�J    	  B                             ������������������������������������������������������                                                                       	                                                                    �      �      �        �        � �          	  
 	 
 	 	 ��������������������� ��������� ������������������� ���� �����������������������������������  � ����������  ����������������������� � ������������ �  ����� � ��� ���������� ������ ������������ ����������� �� �����������                     
     	           $     ��  H�J      ��  	                           ������������������������������������������������������                                                                    
                                                              
       �        �      �        �    ��              
 	  
	 
 	 	 ������������������������� � ������������ ����������������� � � ���������������������� � ��� �������� ����������� � �� ��   � ���� ����������������������������������� ������ ����� �������������������������� ������������ �����������            x                                                                                                                                                                                                                                                                                                           �             


           �   }�         ��������������������������������    ����������������  R������������������������  N���������������������                              Rw                        'u                        �ww�ww333wwwwwwww�ww�ww�ww�ww333wwww I @ 5 
              	                  � 1��� �\                                                                                                                                                                                                                                                                                         	n)n
  1n)�              a      l            b      a      m                                                                                                                                                                                                                                                                                                                                                                                                                  O  � ��  � @��  � ��  � #��  � ��  ��8�������������������9�����y�����������]�����y          :   4 
  ��� 	       	 	 �   & AG� �  �   
           � �                                                                                                                                                                                                                                                                                                                                     p B C   �     p                !��                                                                                                                                                                                                                            Y   	�� �� Ѱ��      �� B 	     ��������������������� ��������� ������������������� ���� �����������������������������������  � ����������  ����������������������� � ������������ �  ����� � ��� ���������� ������ ������������ ����������� �� ������������������������������������ � ������������ ����������������� � � ���������������������� � ��� �������� ����������� � �� ��   � ���� ����������������������������������� ������ ����� �������������������������� ������������ �����������   �� �     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    3      1   � ��                       B     �   ����������      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��     �� p���� ��    ���  �  �(����     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@     H 
o� ��  H 
o� �$ ^$   8 � ��� �� � ��� � �� �  ��  �      �  ��   K�������2����   g��� 	 �     f ^�         ��&       K      ������2�������J��\���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ""   "! " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               ""   "! " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """     " ""   "" !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��   "  " "  ��  �           ���  +"  "" ���������                   �                        ���� ��� ����               �  �  �  �                            �  �˰ ��� �wp ���    �   ��  ���  � �    �                                                                                                                                                   � ""�""�"" ���      � ""+ "" "   ���4 �4ED@�DUT�4DU��3E�4EU�EU\�EU���"+��2"ʀ""��//���/�� �   �   �ɪ��˙�ݹ��ݪ��]����ˊ ̻? ˴?�C��?� ������� �� �  �                �   �     �   �       � "� "  "+���� ��  ݚ                          ��������                          ��  ��  ��  }�  ��  vw� wz� ��� �����        "  ""  ""/ �"� ��          �   �  � �� ��  �                        �   ��  �   ��  ��  �  �  �   �                        �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                        �          �   � � �  ��� ��  �                    �                        ���� ��� ����        �   �   ��� ������ �   �      �       �                        �   ��  ���  � �    �                               �   �                                                                                                                 �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                            ��  ��  ��                          �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������             ��  �   ��  �                                                                                                                                                                                                                               �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �            �  ��  �  �  ��  �                       ����               �   �   �                   �  �  ��  �   �   �        ��  �  �  �   �                                                                                                                                                                                              �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �                              �           �  � � �� ��     �  � � �    �                    ��      �                       �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                     �� ̽ ̽��۽ }�  wz  � ��������ɜ���̚��̸ ��  ��  �  �  T�  T�  H� �E �E �D�[ ˻  ˸  ��  
� ,"�"" �"  �"              "   *�  ��� ��� �ة��ڋ�̽� ��  ��  ̻� ̻� ��� ��@ ��@ DD0 T30 B3� ��  ��  ��  
� +� �"" �"� �" ��� ����  ��          ���    �                       
 "� ""� ""� "                       �                             ���                         �  ��                    �����                       �       �                        �   ��  ���  � �    �                                                                                                                                               �   �  �  �  	�  �  EH  ET DU CE DD4 DD3 DC0 �3 ɰ �  ,�  +�  "/  ������ � ̹�p�˚��̹���ː�̼�̻���ۜ��۩�ݍ���=��J�ܰT�� EJ�0 EJ� I�  ��  �"  ""  "/  "�� ���                    ̰ ̻ ̻	���̚�w��  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                    "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                  ���� �                                                                                                                                                                                          �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw  ��  �   ��  �                                   � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                              �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��               �  �� ��  �    � ���                                                                                                                                                                                              � 
��	�˽���w��{k��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            �  �  �  ��  �            ��  ��                                �  �� �  �  �   �     ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw �   �  ���� �   �             �   ��  ��  ��  �  �   ��  ��                                                                                                                                                                   �  �  �� ̹ ��� ��� ����U���U � U� �� ۻ�������۹�ɧ������٪��̙͉��؝���˳��̽� ˈ� �ɍ �ɀ �ɏ �Ɏ��̎�����      ��  ��  ��� ؙ� ��  ��  �                   �    �������       ���                                    �� ̽ �����ȭ���� (���+�����"/  ��        �  ��  ��� ���� �   ����   �                    ��� ��� ����    �   �   �   ��  �                                            �   �           �   ̰  �˰                                                                                                                                                                                                              �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    DD@DD@                        �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqLC. �dC6 � �kjS � kpS �k~g � k�o �cV> �c^6 � 	ca. �
cb& �C � C"+ �c�U � c�e �c� � c�* � c� � c� � c� y c� �Ci � Cq �J� � � J� � �"� � "�  �"� �*� �"� � "�) �� � 
�" �!"� � ""�) �#� � 
�" � 
�" � 
�! ~'
� q ("J �I  "J q �*!� y/  "  y � ,"�1 �-� �.
�& �  "P � �  "P � �1
�% p2"8 � �  "P � �  "P � �  "P �  6"J �8 !� |@ !� |@ !� |(  "P �(  "P �X <*CT` =*G\`  *K<,  *F�3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.����������������������������������������#� ��9�K�Z�X��5�R�O�S�G� � � � � � � � � � �/�.�7����������������������������������������� ��5�K�\�O�T��=�U�J�J� � � � � � � � � � �/�.�7�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������/�.�7� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $������������������������     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %������������������������ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�A�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                