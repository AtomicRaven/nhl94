GST@�                                                           @r�                                                      ���   ��             
      ����e j�	 ʱ����������`���z���        �h     #    z���                                d8<n    �  ?     ����  �
fD�
�L���"����D"� j   " B   J  jF�"   "�j  ����
��
�"    
 �j� �  
  ��
  Z                                                                               ����������������������������������      ��    bb= QQ0 4 111 44              		 

                     ��� �   � �                 nn ))
         88�����������������������������������������������������������������������������������������������������������������������������  bb    41  c  c  c                    	  
        G  �  (  (                  n�  1)          8= �����������������������������������������������������������������������������                                         �   @  &   }   �                                                                                 '       )n)n
  1n)�    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    A��{	�(:��KD�'�|(	GnToXR�7��4B3�C�TT0 k� �\.�`.!2�$ !A&0   ��    � <�eA��{N��	�$9��KD�#�|(	Gn SoTP�;��0B3�C�PT0 k� �d+�h+!2�$ !A&0   ��    � <�hA��{N��	� 8��KD�#�|(	G]�RoPO�?��(B3�C�LT0 k� �l(�p(!2�$ !A&0   ��    � <�kA��|N��	� 7��KD��|(	G]�RoLN�C�$B3�C�DT0 k� �x%�|%!2�$ !A&0   ��    � <�nA��|N�	�6�KD��|(	G]�QoHL�G� B3�C�@T0 k� ��"��"!2�$ !A&0   ��    � <�qA��|Nw�	�5�KI��|(G]�P_@K�K�B3�D<T0 k� ����!2�$ !A&0   ��    � <�tA��|No��4�KI� |(G]�P_<I�K�B3�D8T0 k� ����!2�$ !A&0   ��    � <�wA��}Ng��3 �KI�|(GM�O_8H�O�B3�D4T0 k� ����!2�$ !A&0   ��    � <�zA��}N_��2 �KI�|(GM�N_4G�S�B3�D,T0 k� ����!2�$ !A&0   ��    � <�}A��}NW��1 �KI�|(GM�M_,E�W�B3�D(T0 k� ����!2�$ !A&0   ��    � ;��A��}NK��0 �KI�|,GM�M�(D�[� B3�D$T0 k� ����!2�$ !A&0   ��    � :��A��~NC��/ �KI�|,GM�L� C�_��B3�DT0 k� ����!2�$ !A&0   ��    � 9��A��~>;��- xKI�|,GM�K�B�c��B3�DT0 k� ��
��
!2�$ !A&0   ��    � 8��A��~>3�� , lKI�|,GM�K�@�g��B3�DT0 k� ����!2�$ !A&0   ��    � 7��A��~>+���+ dKI�|,GM�J�?�g��B3�DT0 k� ����!2�$ !A&0   ��    � 6��A��~>#���) \KE}	|,GM�J�>�k��B3�DT0 k� �� �� !2�$ !A&0   ��    � 5��A��>���( TKE}
|,GM�I�=�o��B3�D T0 k� ������!2�$ !A&0   ��    � 4��A��~>���& LKE}|,GM�H��<�s��B3�D�T0 k� ������!2�$ !A&0   ��    � 2��A��~>���%@KE}|,GM�H��:�w��B3�D�T0 k� ����!2�$ !A&0   ��    � 0��A��~>���#8KE}|,GM�G��9�{��B3�D�T0 k� ����!2�$ !A&0    ��    � .��A��~=����"0KEm|,GM�G��8���B3�D�T0 k� ����!2�$ !A&0    ��    � ,��A��}=��� (KEm|,GM�F��6���B3�D�T0 k� �#��'�!2�$ !A&0    ��    � *��A��}=��� KEm|,GM|F��5����B3�D�T0 k� �+��/�!2�$ !A&0    /�    � (��A��}-���KEm|,GMxE��4���ҨB3�D�T0 k� �3��7�!2�$ !A&0    �    � (��A��}-ߦ��PKEm|,GMtDn�2O��ҤB3�D�T0 k� �;��?�!2�$ !A&0    �    � (��A��|-ק��PKEm|,GMlDn�1O��ҜB3�D�T0 k� �G��K�!2�$ !A&0    ��    � (��A��|-Ө��_�KEm|,E�hCn�/O��ҔB3�D�T0 k� �O��S�!2�$ !A&0    ��    � (��A��|-˩��_�KEm|,E�dCn�.O��ҌB3�C�T0 k� �W��[�!2�$ !A&0    ��    � (��A��|-Ǫ��_�KEm|,E�`Bn�-O��҄B3�C�T0 k� �c��g�!2�$ !A&0    ��    � (��A��|-����_�KEm|,E�XBn�+O���|B3�C�T0 k� �k��o�!2�$ !A&0    ��    � (��A��{-����_�KEm|,E�TAn�*O���tB3�C�T0 k� �s��w�!2�$ !A&0    ��    � (��A��{ m����_�KEm|,E�PAn�(O���lB3�C�T0 k� �{���!2�$ !A&0    ��    � (��A��{ m����_�KEm|,E�L@^�'O���dB3�C�T0 k� ������!2�$ !A&0    ��    � (��A��{ m����_�KA�|,E�H@^�&O���\B3�C�T0 k� ������!2�$ !A&0    ��   � (��A��{ m����_�KA�|,EMD?^�$ ����PB3�C�|T0 k� ������!2�$ !A&0    ��    � (��A��z m����	_�KA�|,EM<?^�# ����HB3�C�tT0 k� ������!2�$ !A&0    ��    � (��A��z m����_�KA� |,EM8>^|" ����@B3�C�lT0 k� ������!2�$ !A&0    ��    � (��A��z m����_�KA�!|,EM4=^x  ����8B3�C�`T0 k� ������!2�$ !A&0    ��    � (��A��z m����_�KA�"|,EM0=^p ����0B3�C�XT0 k� ������!2�$ !A&0    ��    � (��A��z m����_�KA�"|,EM(<^h ����(B3�C�PT0 k� ������!2�$ !A&0    ��    � (��A��y m���_�KA�#|,E=$;^` ���� B3�C�HT0 k� ������!2�$ !A&0    ��    � (��A��y m{���_�KA�$|,E= :^X �û�B3�C�@T0 k� ������!2�$ !A&0    ��    � (��A��y ms��� _�KA�%|,E=9NP �ý�B3�C�4T0 k� ������!2�$ !A&0    ��    � (��A��y mo����_�KA�&|,E=8NL �Ǿ�B3�C�,T0 k� ������!2�$ !A&0    ��    � (��A��y mk����_xKA�'|,E=7ND �˿� B3�C�$T0 k� ������!2�$ !A&0    ��    � (��A��y mg����_tKA�'|,E=7N< �����B3�C�T0 k� ������!2�$ !A&0    ��    � (��A��x mc����_lKA�'|,E=7N4 �����B3�C�T0 k� ������!2�$ !A&0    ��    � (��A��x m[����_hKA�&|,E=7N, �����B3�C�T0 k� ������!2�$ !A&0    ��    � (��A��x mW����_`KA�&|,E= 7N$ �����B3�C� T0 k� ������!2�$ !A&0    ��    � (��A��x mS����_\KA�&|, E,�7N �����B3�C��T0 k� ������!2�$ !A&0    ��    � (��A��x mO����_TKA�&|, E,�6N �����B3�D�T0 k� ������!2�$ !A&0    ��   � (��A��x mK����_PKA�&|, E,�6N �����B3�D�T0 k� ������!2�$ !A&0    ��    � (��A��x mG����_LKA�&|, E,�6N ����B3�D�T0 k� ������!2�$ !A&0    ��    � (��A��w mC����_DKA�&|, E,�6=� ����B3�D�T0 k� ������!2�$ !A&0    ��    � (��A��w m;����_@KA�&|, K��6=� ����B3�D�T0 k� ������!2�$ !A&0    ��    � (��A��w m7����_<KA� &|, K��6=� ����B3�D�T0 k� ������!2�$ !A&0    ��    � (��A��w m3����_4KA� %|, K��5=� ����B3�D�T0 k� ������!2�$ !A&0    ��    � (��A��w m/����_0KA� %|, K��5=� ����B3�D�T0 k� ������!2�$ !A&0    ��    � (��A��w m+����_,KA� %|, K��5=� ����B3�D�T0 k� ������!2�$ !A&0    ��    � (��A��w m'����_$KA��%|, K��5=� ����B3�D�T0 k� ������!2�$ !A&0    ��    � (��A��w m#����_ KA��%|, K��4=� ���xB3�EјT0 k� ������!2�$ !A&0    ��    � (��A��v m����_KA��%|/�K��4=� ���pB3�EьT0 k� ������!2�$ !A&0    ��    � (��A��v m����_KA��%|/�K��4=� ���hB3�EфT0 k� ������!2�$ !A&0    ��    � (��A��v m����_KA��%|/�K��4=� ���`B3�E�|T0 k� ������!2�$ !A&0    ��    � (��A��v m����_KA��$!�/�K��3-� ���XB"s�E�tT0 k� ������!2�$ !A&0    ��    � (��A��v m����_KA��$!�/�K��3-� ���PB"s�E�hT0 k� ������!2�$ !A&0    ��    � (��A��v m����_KA��$!�/�K��3-� ���HB"s�E�`T0 k� ������!2�$ !A&0    ��    � (��A��v m����_ KA��$!�/�K��3-� ���@B"s�E�XT0 k� ������!2�$ !A&0    ��   � (��A��v m����^�KA��$!�/�K��2-� ��8B"s�E�PT0 k� ������!2�$ !A&0    ��    � (��A��u m����^�KA��$!�/�K��2-� ��0B"s�E�HT0 k� ������!2�$ !A&0    ��    � (��A��u m����^�KA��$!�/�K��2-� ��(B"s�D1<T0 k� ������!2�$ !A&0    ��    � (��A��u l�����^�KA��$!�/�K̼2-� �� B"s�D14T0 k� ������!2�$ !A&0    ��    � (��A��u l�����^�KA��$!�/�K̼1-� ��B"s�D1,T0 k� ������!2�$ !A&0    ��    � (��A��u l�����^�KA��$!�/�K̸1-� ��B"s�D1$T0 k� ������!2�$ !A&0    ��    � (��A��u l�����^�KA��#!�/�K̴1�| ��B"s�D1T0 k� ������!2�$ !A&0    ��    � (��A��u l�����^�KA��#|/�K̴1�x ���B3�D1T0 k� ������!2�$ !A&0    ��    � (��A��u l�����^�KA��#|/�K̰1�x ���B3�D1T0 k� ������!2�$ !A&0    ��    � (��A��u l�����^�KA��#|/�K̰0�t ���B3�D1 	T0 k� ������!2�$ !A&0    ��    � (��A��u l�����^�KA��#|/�K̬0�p ����B3�D0�	T0 k� �����!2�$ !A&0    ��    � (��A��t l�����^�KA��#|/�K̬0�l ����B3�D0�
T0 k� �����!2�$ !A&0    ��    � (��A��t l�����^�KA��#|/�K̨0�l ����B3�D0�
T0 k� ����!2�$ !A&0    ��    � (��A��t l�����^�KA��#|/�K̨0�h ����B3�D0�T0 k� ����!2�$ !A&0    ��    � (��A��t l�����^�KA��#|/�K̤/�h ����B3�D@�T0 k� ����!2�$ !A&0    ��    � (��A��t l�����^�KA��#|/�K̤/�d ���B3�D@�T0 k� ����!2�$ !A&0    ��    � (��A��t l�����^�KA��#|/�K̠/�d ���B3�D@�T0 k� ����!2�$ !A&0    ��    � (��A��t l�����^�KA��#|/�K̠/�` ���B3�D@�T0 k� ����!2�$ !A&0    ��    � (��A��t l�����^�KA��#!�/�K̜/` ���B"��D@�T0 k� ����!2�$ !A&0    ��    � (��A��t l�����^�KA��"!�/�K̜/\ ����B"��D@�T0 k� ����!2�$ !A&0    ��    � (��A��t l�����^�KA��"!�/�K̘.\ �#���B"��D@�T0 k� ����!2�$ !A&0    ��    � (��A��t l�����^�KA��"!�/�K̘.\ �#���B"��D@�T0 k� ����!2�$ !A&0    ��    � (��A��t l�����^�KA��"!�/�K̔.\ �'���B"��D@�T0 k� ����!2�$ !A&0    ��   � (��A��t l�����^�KA��"!�/�K̔.\  �'��xB"��D@�T0 k� ����!2�$ !A&0    ��    � (��A��s l�����^�KA��"!�/�K̔.\! �'��pB"��D@�T0 k� ����!2�$ !A&0    ��    � (��A��s l�����^�KA��"!�/�K̐.X"�+��hB"��DPxT0 k� ����!2�$ !A&0    ��    � (��A��s l�����^�KA��"!�/�K̐-X#�+��`B"��DPpT0 k� ���#�!2�$ !A&0    ��    � (��A��s l�����^�KA��"!�/�Ǩ-X$�+��XB"��DPhT0 k� ���#�!2�$ !A&0    ��    � (��A��s l�����^�KA��"!�/�Ǩ--\%�+��PB"��DP`T0 k� ���#�!2�$ !A&0    ��    � (��A��s l�����^�KA��"|/�Ǩ--\&�/��HB3�DPXT0 k� �#��'�!2�$ !A&0    ��    � (��A��s l�����^�KA��"|/�K̈--\'�/��<B3�DPPT0 k� �#��'�!2�$ !A&0    ��    � (��A��s l����^�KA��"|/�K̈--\)�/��4B3�DPHT0 k� �#��'�!2�$ !A&0    ��    � (��A��s l����^�KA��"|/�K̄--\*�3��,B3�DP@T0 k� �'��+�!2�$ !A&0    ��    � (��A��s l����^�KA��"|/�K̄,-\+�3� $B3�DP8T0 k� �'��+�!2�$ !A&0    ��    � (��A��s l����^�KA��!|/�K̄,-`,�3� B3�DP0T0 k� �'��+�!2�$ !A&0    ��    � (��A��s l����^�KA��!|/�K̀,-`.�7� B3�DP(T0 k� �+��/�!2�$ !A&0    ��    � (��A��s l����^�KA��!|/�K̀,`/�7� B3�D` T0 k� �/��3�!2�$ !A&0    ��    � (��A��s l���{�^�KA��!|/�K̀,d0�7� B3�D`T0 k� �/��3�!2�$ !A&0    ��    � (��A��s l���{�^�KA��!|/�K�|,d1�7��B3�D`T0 k� �/��3�!2�$ !A&0    ��    � (��A��r l���{�^�KA��!|/�K�|,h2�;��B3�D`T0 k� �/��3�!2�$ !A&0    ��    � (��A��r l���{�^|KA��!|/�K�|+h4�;��B3�D`  T0 k� �3��7�!2�$ !A&0    ��    � (��A��r l���{�^|KA��!|/�K�x+�l5�;��B3�L?�!T0 k� �3��7�!2�$ !A&0    ��    � (��A��r l���{�^xKA��!|/�K�x+�p6�;��B3�L?�"T0 k� �3��7�!2�$ !A&0    ��    � (��A��r l���{�^xKA��!|/�K�x+�t7�?��B3�L?�#T0 k� �3��7�!2�$ !A&0    ��    � (��A��r l���w�^tKA��!|/�K�t+�t8�?��B3�L?�$T0 k� �7��;�!2�$ !A&0    ��    � (��A��r l���w�^tKA��!|/�E,t+�x9�?��B3�L?�$T0 k� �7��;�!2�$ !A&0    ��    � (��A��r l���w�^pKA��!|/�E,t+�|:�?��B3�L?�%T0 k� �7��;�!2�$ !A&0    ��    � (��A��r l���w�^pKA��!|/�E,t*��;�C��B3�L?�&T0 k� �7��;�!2�$ !A&0    ��    � (��A��r l���w�^lKA��!|/�E,t*��<�C��B3�L?�'T0 k� �;��?�!2�$ !A&0    ��    � (��A��r l���w�^lKA��!|/�E,t*��=�C��B3�L?�(T0 k� �;��?�!2�$ !A&0    ��    � (��A��r l���w�^hKA��!|/�@t*��>�C��B3�L?�(T0 k� �;��?�!2�$ !A&0    ��    � (��A��r l���s�^hKA��!|/�@t)��?�C��B3�L?�)T0 k� �;��?�!2�$ !A&0    ��    � (��A��r l���s�^dKA��!|/�@t)��@�G�_�B3�L?�*T0 k� �?��C�!2�$ !A&0    ��    � (��A��r l���s�^dKA��!|/�@t)��A�G�_�B3�LO�+T0 k� �?��C�!2�$ !A&0    ��    � (��A��r l���s�^`KA��!|/�@x)��B�G�_xB3�LO�+T0 k� �?��C�!2�$ !A&0    ��    � (��A��r l���s�^`KA��!|/�@x)��C�G�_pB3�LO�,T0 k� �?��C�!2�$ !A&0    ��    � (��A��r l���s�^\KA�� |/�B�x(��D�G�_dB3�LO�-T0 k� �?��C�!2�$ !A&0    ��    � (��A��r l���s�^\KA�� |/�B�|(��E�K�\B3�LO�.T0 k� �C��G�!2�$ !A&0    ��    � (��A��r l���s�^\KA�� |/�B�|(��F�K�TB3�LO�.T0 k� �C��G�!2�$ !A&0    ��    � (��A��r l���s�^XKA�� |/�B��(��F�K�LB3�LO�/T0 k� �C��G�!2�$ !A&0    ��    � (��A��r l���o�^XKA�� |/�B��(��G�K�HB3�LOx0T0 k� �C��G�!2�$ !A&0    ��    � (��A��q l���o�^TKA�� |/�B��'��H�K�@B3�LOt0T0 k� �C��G�!2�$ !A&0    ��    � (��A��q l���o�^TKA�� |/�B��'��I�O�8B3�LOp1T0 k� �G��K�!2�$ !A&0    ��    � (��A��q l��o�^TKA�� |/�B��'��J�O�0B3�LOh2T0 k� �G��K�!2�$ !A&0    ��    � (��A��q l��o�^PKA�� |/�B��'��K�O�(B3�LOd2T0 k� �G��K�!2�$ !A&0    ��    � (��A��q l��o�^PKA�� |/�B��'��K�O� B3�LO`3T0 k� �G��K�!2�$ !A&0    ��    � (��A��q l��o�^LKA�� |/�B��'��L�O�B3�LOX3T0 k� �G��K�!2�$ !A&0    ��    � (��A��q l{��o�^LKA�� |/�B��'��M�S�B3�LOT4T0 k� �K��O�!2�$ !A&0    ��    � (��A��q l{��o�^LKA�� |/�B��(��N�S�B3�LOP5T0 k� �K��O�!2�$ !A&0    ��    � (��A��q l{��o�^HKA�� |/�B��(��N�S�B3�LOL5T0 k� �K��O�!2�$ !A&0    ��    � (��A��q lw��k�^HKA��|/�B��(��O�S�/ B3�LOD6T0 k� �K��O�!2�$ !A&0    ��    � (��A��q lw��k�^HKA��|/�B��(�P�S�.�B3�LO@6T0 k� �K��O�!2�$ !A&0    ��    � (��A��q lw��k�^DKA��|/�B��(�P�S�.�B3�LO<7T0 k� �K��O�!2�$ !A&0    ��    � (��A��q lw��k�^HKA��|/�B��(�P�W�.�B3�LO87T0 k� �K��O�!2�$ !A&0    ��    � (��A��q ls��k�^HKA��|/�B��(�Q�W�.�B3�LO48T0 k� �O��S�!2�$ !A&0    ��    � (��A��q ls��k�^HKA��|/�B��(�R�W�.�B3�LO09T0 k� �O��S�!2�$ !A&0    ��    � (��A��q ls��k�^LJA��|/�B��(�S�W�.�B3�LO,9T0 k� �O��S�!2�$ !A&0    ��    � (��A��q ls��k�^LJA��|/�B��(�T�W�.�B3�LO$:T0 k� �O��S�!2�$ !A&0    ��    � (��A��q lo��k�^LJA��|/�B��)�U�W�.�B3�LO :T0 k� �O��S�!2�$ !A&0    ��    � (��A��q lo��k�^LJA��|/�B̴)�U�W�.�B3�LO;T0 k� �O��S�!2�$ !A&0    ��    � (��A��q lo��k�^PIA��|/�B̸)�V�[�.�B3�LO;T0 k� �S��W�!2�$ !A&0    ��    � (��A��q lo��k�^PIA��|/�B̸)� W�[�.�B3�LO<T0 k� �S��W�!2�$ !A&0    ��    � (��A��q lk��g�^PIA��|/�B̼)� X�[�.�B3�LO<T0 k� �S��W�!2�$ !A&0    ��    � (��A��q lk��g�^TIA��|/�B��)�$Y�[�.�B3�LO=T0 k� �S��W�!2�$ !A&0    ��    � (��A��q lk��g�^THA��|/�B��*�(Y�[�.�B3�LO=T0 k� �S��W�!2�$ !A&0    ��    � (��A��q lk��g�^THA��|/�B��*�,Z�[�.�B3�LO=T0 k� �S��W�!2�$ !A&0    ��    � (��A��q lk��g�^THA��|/�B��*�,[ �[�.�B3�LO >T0 k� �L�P!2�$ !A&0    ��    � (��A��q lg��g�^XHA��|/�B��*�0[ �[�.�B3�LN�>T0 k� �L�P!2�$ !A&0    ��    � (��A��q lg��g�^XGA��|/�B��*�4\ �_�.�B3�LN�?T0 k� �P�T!2�$ !A&0    ��    � (��A��q lg��g�^XGA��|/�B��+�4] �_�.�B3�LN�?T0 k� �P	�T	!2�$ !A&0    ��    � (��A��q lg��g�^XGA��|/�B��+�8^ �_�.�B3�LN�@T0 k� �P�T!2�$ !A&0    ��    � (��A��q lg��g�^TGA��|/�B��+�8^ �_�.�B3�LN�@T0 k� �P�T!2�$ !A&0    ��    � (��A��q lc��g�^TGA��|/�B��+�<_ �_�.�A3�LN�@T0 k� �P�T!2�$ !A&0    ��    � (��A��q lc��g�^PGA��|/�B��+�@` �_�.�A3�LN�AT0 k� �P�T!2�$ !A&0    ��   � (��A��q lc��g�^PGA��|/�B��+�@` �_�.�A3�L>�AT0 k� �P�T!2�$ !A&0    ��    � (��A��q lc��g�^PGA��|/�B� ,�Da �\ .�A3�L>�BT0 k� �P�T!2�$ !A&0    ��    � (��A��q lc��g�^LGA��|/�B�,�Da �` .�A3�L>�BT0 k� �T�X!2�$ !A&0    ��    � (��A��q l_��c�^LGA��|/�B�,�Hb �` .�A3�L>�BT0 k� �T�X!2�$ !A&0    ��    � (��A��q l_��c�^HGA��|/�B�,�Lc �` .�@3�L>�CT0 k� �T�X!2�$ !A&0    ��    � (��A��q l_��c�^HGA��|/�E,�Lc �` .�@3�L>�CT0 k� �T�X!2�$ !A&0    ��    � (��A��q l_��c�^HGA� |/�E ,�Pd �`.�@3�D>�DT0 k� �T�X!2�$ !A&0    ��    � (��A��p l_��c�^DGA� |/�E0-�Te �`.�@3�D>�DT0 k� �T�X!2�$ !A&0    ��    � (��A�|p l[��c�^@GA� |/�E4-�Tf �`.�?3�D>�ET0 k� �T�X!2�$ !A&0    ��    � (��A�|p l[��c�^@GA�|/�K�<-�Xf �`.�?3�D>�ET0 k� �T�X!2�$ !A&0    ��    � (��A�|p l[��c�^@GA�|/�K�D-�Xg �`.|?3�E��FT0 k� �T�X!2�$ !A&0    ��   � (��A�|p l[��c�^<GA�|/�K�H-�\g �d.|?3�E�GT0 k� �T�X!2�$ !A&0    ��    � (��A�|p l[��c�^<HA�|/�K�P.�\h �d.|?3�E�GT0 k� �T�X!2�$ !A&0    ��    � (��A�|p l[��c�^<HA�|/�K�T.�`h �d.x?3�E�HT0 k� �T�X!2�$ !A&0    ��    � (��A�|p lW��c�^8HA�|/�K�\.�`i �d.x>3�E�IT0 k� �T�X!2�$ !A&0    ��    � (��A�|p lW��c�^8HA�|/�K�`.�di �d.t>3�E��IT0 k� �T�X!2�$ !A&0    ��    � (��A�|p lW��c�^8HA�|/�K�h.�dj �dt>3�E��JT0 k� �T�X!2�$ !A&0    ��    � (��A�|p lW��c�^4HA�|/�K�l.�hj �dt>3�E��KT0 k� �T�X!2�$ !A&0    ��    � (��A�|p lW��c�^4HA�|/�K�t.�hk �dp>3�E��LT0 k� �T�X!2�$ !A&0    ��    � (��A�|p lW��c�^4HA�|/�K�x.�lk �dp>3�E��MT0 k� �T�X!2�$ !A&0    ��    � (��A�|p lW��c�^0HA�|/�K��/�ll �dp>3�D��MT0 k� �T�X!2�$ !A&0    ��    � (��A�|p lS��c�^0HA�|/�K��/�ll �dl=3�D��NT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lS��c�^0HA�|/�K��/�pm �h^l=3�D��OT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lS��_�^0HA�|/�K��/�pm �h^h=3�D��OT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lS��_�^,HA�|/�K��/�tn �h^h=3�D��PT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lS��_�^,HA�|/�K��/�tn �h^d=3�D��PT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lS��_�^,HA�|/�K��/�tn �h^d=3�D��PT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lS��_�^(HA�|/�K��/�xo �hN`=3�D��QT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lS��_�^(HA�|/�K��0�xo �hN\=3�D��QT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lO��_�^(HA�|/�K��0�|p �hN\=3�L^�QT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lO��_�^(HA�|/�K��0�|p �hNX=3�L^�RT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lO��_�^$HA�|/�K��0�|p �hNT=3�L^�RT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lO��_�^$HA�|/�K��0��q �hNT=3�L^�RT0 k� �X�\!2�$ !A&0    ��    � (��A�|p lO��_�^$HA�|/�K��0��q �hNT=3�L^�ST0 k� �X�\!2�$ !A&0    ��    � (��A�|p lO��_�^ HA�|/�K��0��r �lNP=3�L^�ST0 k� �\�`!2�$ !A&0    ��    � (��A�|p lO��_�^ HA�|/�K��0��r �l>P=3�L^|ST0 k� �\�`!2�$ !A&0    ��    � (��A�|p lO��_�^ HA�|/�K��0��r �l>P=3�L^|TT0 k� �\�`!2�$ !A&0    ��    � (��A�|p lO��_�^IA�|/�K��1��s �l>P=3�L^|TT0 k� �\�`!2�$ !A&0    ��    � (��A�|p lO��_�^IA�|/�K��1��s �l>L=3�L^xTT0 k� �\�`!2�$ !A&0    ��    � (��A�|p lK��_�^IA� |/�K��1��s �l>L>3�L^xTT0 k� �\�`!2�$ !A&0    ��    � (��A�|p lK��_�^IA� |/�K��1��t �l>H>3�L^xUT0 k� �\�`!2�$ !A&0    ��    � (��A�|p lK��_�^IA� |/�K��1��t �l.H?3�L^tUT0 k� �\�`!2�$ !A&0    ��    � (��A�|p lK��_�^JA� |/�K��1�t �l.D?3�L^tUT0 k� �\�`!2�$ !A&0    ��    � (��E��\��`H�8WEb8&|( C�$dSFcPS�I�C��T0 k� �A�A!2�$ !A&0    ��3    � $ �E��Z��XH�4WEb8'|( C� c� F3P
�I�C��T0 k� �A�A!2�$ !A&0    ��3    � % �E��Y��LG�0WEb8(|( C�b� F3P	�H�C��T0 k� �A�A!2�$ !A&0    ��3    � & �E��V��8G�0WER8*|( E3_��E3L�G�C��T0 k� �A� A!2�$ !A&0    ��3    � ' �E��U�
�,F�,WER8+|( E3^��E3L�F�C��T0 k� � @�$@!2�$ !A&0    ��3    � ( �E��S�	�$F�(WER8,|( E3\��E3L	��F�C��T0 k� �$@�(@!2�$ !A&0    ��3    � ) �EB�S��E$WER8-|( E3\��E3L	��E�A�T0 k� � @�$@!2�$ !A&0    ��3    � * �EB�Q��DVER8/|( E3Y��C3H	��D�A�T0 k� �@�@!2�$ !A&0    ��3    � + �EB�P��DVER40|( E3 W��C3D	��D�A�T0 k� �?�?!2�$ !A&0    ��3    � , �EB�O��CVER41|( E2�U2�B3D	��D�A�T0 k� �?�?!2�$ !A&0    ��3    � - �EB�N ��CUER42|( E2�T2�A3G�	��C�A�T0 k� �>�>!2�$ !A&0    ��3    � - �EB�K  ��B�TER04|( E2�T2�?CC�	��C�A�T0 k� ��>��>!2�$ !A&0    ��3    � - �EB�J���B� TEB,5|( CB�S2�=CC�	��C�C��T0 k� ��?��?!2�$ !A&0    ��3    � - �EB�I����A��SEB,6|( CB�RR�<C?�	�|B�C��T0 k� ��?��?!2�$ !A&0    ��3    � - �EB�H����A��SEB(7|( CB�PR�;C?�	�xB�C��T0 k� ��?��?!2�$ !A&0    ��3    � - �EB�E��Ѱ@��REB$8|( CB�NR�8C?�	�tB�	C��T0 k� ��>��>!2�$ !A&0    ��3    � - �E2�D��Ѩ?��QEB$9|( CB�LR�7C?�	�tB�	C��T0 k� ��=��=!2�$ !A&0    ��3    � - �E2�B���?��QEB :|( CB�KR�6C?�	�pB�	C��T0 k� ��=��=!2�$ !A&0    ��3    � - �E2�A���?��PEB:|( CB�IR�5C;�	�pB�	C��T0 k� ��<��<!2�$ !A&0    ��3    � - �E2t>���>��PE2;|( CB�FR�2C;�	�lB3�	C��T0 k� ��:��:!2�$ !A&0   �3    � - �E2l<����|=��OE2<|( E��DR�1S;�	�lB3�	C��
T0 k� ��9��9!2�$ !A&0   ��?    � - �E2h;����t=��OE2<|( E��C�0S;�	�hB3�	C��
T0 k� ��8��8!2�$ !A&0   ��?    � - �E2d9����l=��NE2<|( E��A�/S;�	�hB3�
C��	T0 k� �7�7!2�$ !A&0   ��?    � - �E2X6����\<��NE2=|( E��=�-S?�	�hB3�
C��	T0 k� �5� 5!2�$ !A&0   ��?    � - �E2T4���T<��MCB=|( E��<�,SC�	�dB3�
C��T0 k� �,4�04!2�$ !A&0   ��?    � - �E2L2���L;��MCB=|( E��:�+SC�	�dB3�
C��T0 k� �83�<3!2�$ !A&0   ��?    � - �E"H0��D;��LCB=|( E¼8�*SG�	�dB3�EӀT0 k� �D2�H2!2�$ !A&0   ��?    � - �E"D/��8:��LCB=|( E¸6�)SG�	�dB3�EӀT0 k� �P1�T1!2�$ !A&0   ��?    � - �E"@-��0:��LCB =|( E´4�)SG�	�dB3�E�|T0 k� �\0�`0!2�$ !A&0   ��?    � - �E"4)�� 9��KCA�=|( E´4�t&SK�	�dB3�E�xT0 k� �t.�x.!2�$ !A&0   $�?    � - �E",(��9��KCA�<|( E°2�l%cK�	�dB3�E�tT0 k� 2p.�t.!2�$ !A&0   ��?    � - �E"(&��8��JCA�<|( EҨ1Rh$cO�	�dB3�E�pT0 k� 2l/�p/!2�$ !A&0   ��?    � - �E"$$��8��JCA�<|( EҤ/Rh$cO�	�dB3�E�pT0 k� 2h/�l/!2�$ !A&0   ��?    � - �E" "�� 8��JCA�;|( EҠ-Rd"cO�	�dB3�E�lT0 k� 2d/�h/!2�$ !A&0   ��?    � - �E" ���7��ICA�;|( EҜ,R`!cO�SdB3�E�hT0 k� 2d/�h/!2�$ !A&0   ��?    � - �E"���7��ICQ�;|( EҜ,R\ cO�SdB3�E�dT0 k� �`/�d/!2�$ !A&0   ��?    � - �E"���6��HCQ�:|( EҔ*RPcO�SdB3�E�`T0 k� �X/�\/!2�$ !A&0   ��?    � - �E���5��HCQ�9|( EҌ(RLcO�SdB3�E�\T0 k� �T/�X/!2�$ !A&0   ��?    � - �E#���4��HCQ�8|( E҈'RDcO�SdB3�E�XT0 k� �P/�T/!2�$ !A&0   ��?    � - �E '���4��GCQ�8|( E҄&R@cK�SdB3�E�TT0 k� "L0�P0!2�$ !A&0   ��?    � - �E�'���3��GCQ�7|( E�|$R<3K�SdB3�E�PT0 k� "H0�L0!2�$ !A&0   ��?    � - �E�+��2��GCQ�6|( E�x#	�83K�SdB3�E�LT0 k� "D0�H0!2�$ !A&0   ��?    � - �E�/��1��FCQ�5|( E�x#	�83G�SdB3�E�DT0 k� "<0�@0!2�$ !A&0   ��?    � - �E�/��0�FCQ�4|( E�t"	�43G�SdB3�E�@T0 k� B@2�D2!2�$ !A&0   ��6    � - �E�3��/�ECa�3|( E�p!	�0cG�SdB3�E�@T0 k� B@2�D2!2�$ !A&0   ��6    � - �E�
3��.�|ECa�2|( E�h 	�,cC�SdB3�E�<T0 k� B<2�@2!2�$ !A&0   ��6    � - �E�7���,�xCCa�0|( E�h �$c?�SdB3�
E�4T0 k� B82�<2!2�$ !A&0   ��6    � - �E�;��|+�tCCa�/|( E�` � c?�SdB3�
F0T0 k� �42�82!2�$ !A&0   ��6    � - �E��;��t*tBE��.|( E�\�c;�SdB3�
F0T0 k� �42�82!2�$ !A&0   ��6    � - �E��?��l(pAE��,|( E�T�c;�SdB3�
F,T0 k� �02�42!2�$ !A&0   ��6    � - �E���C� `&l@E��*|( E�L�c7�SdB3�
F(	T0 k� �(1�,1!2�$ !A&0    -�6    � - �E���G� X%l?E��)|( E�D�c3�SdB3�	F$
T0 k� �$0�(0!2�$ !A&0    ��6    � - �E����G� T$l>E��(|( E�<�
S3�SdB3�	F$T0 k� �0� 0!2�$ !A&0    ��6    � - �E����K� L"h=E��'|( E�8�
S/�SdB3�	E�$T0 k� �$0�(0!2�$ !A&0    ��6    � - �E����S�p@ h;E��$|( E�,��S+�SdB3�	E� T0 k� � /�$/!2�$ !A&0   ��6    � - �E����W�p<h:E��#|( E�(a�S'�SdB3�	E� T0 k� 2 /�$/!2�$ !A&0   ��6    � - �E����[�p4�h9E��"|( E� a�S#�SdB3�	E� T0 k� 2 /�$/!2�$ !A&0   ��6    � - �E����[�p0�h8E�� |( E�a�S�SdB3�	E� T0 k� 2/� /!2�$ !A&0   ��6    � - �E����c�p$�h6E��|( E�a�S�SdB3�	E�T0 k� 20�0!2�$ !A&0   ��6    � - �E����g�p�h5E��|( E�a� ��SdB3�	E� T0 k� "0�0!2�$ !A&0   ��6    � - �E���sk���h4E��|( E�a����SdB3�	E� T0 k� "0�0!2�$ !A&0   ��6    � - �Eq��so���l3E��|( E� a����SdB3�	E� T0 k� "1�1!2�$ !A&0   ��6    � - �Eq��sw���l1EѤ|( E��a�����SdB3�	E� T0 k� "2�2!2�$ !A&0   ��6    � - �Eq��s{���t0EѤ|( E��Q�����SdB3�	E�$T0 k� � 2�2!2�$ !A&0   ��6    � - �Eq��s����|0EѠ|( F� Q�����SdB3�	E�$T0 k� � 1�1!2�$ !A&0   ��6    � - D���s������/Eќ|( F� Q����SdB3�	E�$T0 k� �1�1!2�$ !A&0   ��6    � - |D���s���
��.Eј|( F�!Q����SdB3�	E�(T0 k� �0�0!2�$ !A&0   ��6    � - yD���s�����,Eѐ|( F�#Q���߀SdB3�	E�,T0 k� � 1�1!2�$ !A&0    ��6    � - vD���s�����,Eш|( Eq�#Q���ہSdB3�	B�,T0 k� ��4��4!2�$ !A&0    �6    � - vD���s����,C�|( Eq�#Q���ӁSdB3�	B�0T0 k� !�5��5!2�$ !A&0    ��6    � - uD���s����,C�|( Eq�#Q���ˁSdB3�	B�0T0 k� !�6��6!2�$ !A&0    /�6    � - tD���c�����-C�|
|( Eq�#Q���ǂSdB3�	B�4T0 k� !�7��7!2�$ !A&0    ��6    � - sD���c�����-C�x	|( Eq�#Q���SdB3�	B�4T0 k� !�8��8!2�$ !A&0    ��6    � - rD���c�����-C�p|( Eq�$A{��SdB3�	B�8T0 k� !�9��9!2�$ !A&0    ��6    � - qD���c�����-C�l|( Eq�$Aw��SdB3�	E�<T0 k� ��9��9!2�$ !A&0    ��6    � - pD���c�����-C�`|( Eq�%Ag��SdB3�	E�@T0 k� ��:��:!2�$ !A&0    ��6    � - oD���c������-C�\|( Eq�&A_��SdB3�	E�DT0 k� ��;��;!2�$ !A&0    ��6    � - nD���c������-C�T|( Ea�&AW��SdB3�	E�HT0 k� ��:��:!2�$ !A&0    ��6    � - mD���c������-C�P|( Ea�'AO��SdB3�	E�LT0 k� ��9��9!2�$ !A&0    ��6    � - lD���c������-C�H |( Ea�(AG���SdB3�	E�PT0 k� ��9��9!2�$ !A&0    ��6    � - jD���c������-C�G�|( Ea�)A?�{�SdB3�	E�PT0 k� ��9��9!2�$ !A&0    ��6    � - iD���c������-C�?�|( Ea�)A;�s�SdB3�	E�TT0 k� ��9��9!2�$ !A&0    ��6    � - hD���S������.C�;�|( Ea�*A3�k�SdB3�	E�XT0 k� ��9��9!2�$ !A&0    ��6    � - fD���S������.C�3�|( Ea�+A+�c�SdB3�	E�\T0 k� ��:��:!2�$ !A&0    ��6    � - dD���S������.C�+�|( EQ�,1#�[�SdB3�	CC`T0 k� ��5��5!2�$ !A&0    ��6    � - bD���S������.C�'�|( EQ�,1�S�SdB3�	CC`T0 k� ��1��1!2�$ !A&0    ��6    � - `D���S������.C��|( EQ�,1�C�SdB3�	CChT0 k� ��.��.!2�$ !A&0    ��6    � - ^D���S������.C��|( EQ�-1�7�SdB3�	CChT0 k� ��,��,!2�$ !A&0    ��6    � - \D���S������/C��|( Aa�.0��/�SdB3�	CClT0 k� ��-��-!2�$ !A&0    ��6    � - ZD���S������/C��|( Aa�.0��R'�SdB3�	CClT0 k� ��-��-!2�$ !A&0    ��6    � - XD���S������/D ��|( Aa�.@��R�SdB3�	CCpT0 k� ��-��-!2�$ !A&0    ��6    � - WD���㯋����/D ��|( Aa�.@��R�SdB3�	CCpT0 k� ��-��-!2�$ !A&0    ��6    � - VD���㫉����/D ��|( Aa�.@��R�SdB3�	CCtT0 k� ��-��-!2�$ !A&0    ��6    � - UD���㫈�����/D ��|( Aa�/@��R�SdB3�	CCtT0 k� ��-��-!2�$ !A&0    ��6    � - TEq��㧆�����/D ��|( Aa�/@��Q��SdB3�	CStT0 k� ��.��.!2�$ !A&0    ��6    � - SEq��㧅�����/D ��|( Aa�0@��Q�SdB3�	CSxT0 k� ��/��/!2�$ !A&0    $�6    � - REq��㣃�����0D ��|( Aa�1@��Q�SdB3�	CSxT0 k� 1�/��/!2�$ !A&0    ��6    � - QEq��㟀�����0D ��|( Aa�2@��Q׋SdB3�	CSxT0 k� 1�0��0!2�$ !A&0    ��6    � - PEq��㛁�����0D ��|( Aq�2@��QϋSdB3�	CSxT0 k� 1�/��/!2�$ !A&0    ��6    � - OEq��㗁�����0D ��|( Aq�2@��AǋSdB3�	CSxT0 k� 1�/��/!2�$ !A&0    ��6    � - NEq��㓁�����0D��|( Aq�3@��A��SdB3�	CSxT0 k� ��/��/!2�$ !A&0    ��6    � - MEq��㏂�����0D��|( Aq�3P��A��SdB3�	CSxT0 k� ��/��/!2�$ !A&0    ��6    � - LEa�������0D��|( Aq�4P��A��SdB3�	CSxT0 k� ��0��0!2�$ !A&0    ��6    � - KEa�������0D��|( E��5P��A��SdB3�	@�xT0 k� ��7��7!2�$ !A&0    �6    � - KEa�������0D��|( E��6P��ћ�SdB3�	@�xT0 k� ��<��<!2�$ !A&0    ��6    � - KEa��������0D��!�( E��7P��ѓ�SdB"��	@�xT0 k� ��A��A!2�$ !A&0    ��6    � - KEa��{������0D��!�( E��8P��ч�SdB"��	@�xT0 k� ��E��E!2�$ !A&0    ��6    � - KEa��w�O����0D��!�( E��9P���SdB"��	@�xT0 k� ��H��H!2�$ !A&0    ��6    � - KE��
�s�@��0D��!�( E��:P��w�SdB"��	CCxT0 k� ��K��K!2�$ !A&0    ��6    � - KE���k�@��0D��!�( E��;0{��o�SdB"��	CCxT0 k� ��M��M!2�$ !A&0    ��6    � - KE���g�@��0D{�!�( E��<0s��g�SdB"��	CCxT0 k� ��O��O!2�$ !A&0    ��6    � - KE���[�@��0C�k�!�( A��>0k��S�SdB"��	CCxT0 k� ��O��O!2�$ !A&0    ��6    � - KE��W�@��0C�c�!�( A��?0c��K�SdB"��	CCxT0 k� ��O��O!2�$ !A&0    ��6    � - KE��S�@��0C�W�!�( A��A0_��C�SdB"��	CCxT0 k� ��P��P!2�$ !A&0    ��6    � - KE��K�@��0C�O�!�( A��B0[�A;�SdB"��	CCx
T0 k� ��P��P!2�$ !A&0    ��6    � - JE��G�@��0C�G�|( A��C0W�A/�SdB3�	CCx
T0 k� ��P��P!2�$ !A&0    ��6    � - IE��?�@��0C�?�|( A��E0O�A'�SdB3�	CCx	T0 k� ��R��R!2�$ !A&0    ��6    � - HEa�7�@��0C�7�|( A��F0O�A�SdB3�	CCxT0 k� ��S��S!2�$ !A&0    ��6    � - GEa�3�P��0C�/�|( A��G0K�A�SdB3�	CSxT0 k� ��T��T!2�$ !A&0    ��6    � - FEa�+�P��0C�#�|( A��I G�A�SdB3�	CSxT0 k� ��V��V!2�$ !A&0    ��6    � - EEa� #�P��0C��|( A��J C�A�SdB�	CSxT0 k� ��W��W!2�$ !A&0    ��6    � - DEa� �P��1C��|( A��L ?�@��SdB�	CSxT0 k� ��Y��Y!2�$ !A&0    ��6    � - CEa�!�P��2C��|( A��M ;�@�SdB�	CSxT0 k� ��Z��Z!2�$ !A&0    ��6    � - BEa�"�P��3C��|( A��O 7���SdB�
CSxT0 k� ��\��\!2�$ !A&0    ��6    � - AEa�#�P��3C���|( A��P 3���SdB�
CSxT0 k� ��]��]!2�$ !A&0    ��6    � - @Ea�#�P��4C���|( A��R 3��ەSdB�
CSxT0 k� ��_��_!2�$ !A&0    ��6    � - ?EQ�#��P��5C���!�( A��S /��ӕSdB"C�
CSxT0 k� ��a��a!2�$ !A&0    ��6    � - >EQ�$�P��6C���!�( A��U /��˖SdB"C�
CSxT0 k� ��b��b!2�$ !A&0    ��6    � - =EQ�%�P#��7Eo��!�( A��W�+����SdB"C�
CSxT0 k� ��d��d!2�$ !A&0    ��6    � . <EQ�&ۊ`#���8Eo��!�( Ea�Z�'����SdB"C�CcxT0 k� ��g��g!2�$ !A&0    ��6    � / ;C��'ӊ`#���9Eo��!�( Ea�\�'����SdB"C�CcxT0 k� ��i��i!2�$ !A&0    ��6    � 0 9C��(ˊ`#���:Eo��!�( Ea�]�'����SdB"C�CcxT0 k� ��k��k!2�$ !A&0    ��6    � 1 7C��)Ê`#���;Eo��!�( Ea�_�#����SdB"C�CcxT0 k� ��l��l!2�$ !A&0    ��6    � 2 5C��)⻊`'���<Eo��!�( Ea�`�#�Џ�SdB"C�CcxT0 k� ��n��n!2�$ !A&0    ��6    � 3 3C��*ⳋ`'���<Eo��!�( EQ�b�#�Ї�SdB"C�@�xT0 k� ��i��i!2�$ !A&0    ��6    � 4 1E��+⧋`'���=E��!�( EQ�c�#���SdB"C�@�xT0 k� ��f��f!2�$ !A&0    ��6 	   � 5 /E��,⟋`'���>E��|( EQ�e�#��s�SdB�@�xT0 k� ��d��d!2�$ !A&0    ��6 	   � 6 -E��,○`'���>E��|( EQ�f�#��k�SdB�@�xT0 k� �|c��c!2�$ !A&0    ��6 	   � 7 +E��-⏋`'���?E��|( EQ�h�#��c�SdB�@�xT0 k� �xb�|b!2�$ !A&0    ��6 	   � 8 )E��.⇋p'���@E��|( EQ�i #��[�SdB�@�xT0 k� �tc�xc!2�$ !A&0    ��6 	   � 9 'E�/�{�p+���AE��|( EQ�j   �S�SdB�@�xT0 k� �pc�tc!2�$ !A&0    ��6 	   � : %E�0�s�p+���AE�|( EQ�l  �K�SdB�AxT0 k� �lc�pc!2�$ !A&0    ��6 	   � ; #E�1�k�p+���BE{�|( EQ�m  �C�SdB�AxT0 k� �dd�hd!2�$ !A&0    ��6 	   � < !E�2�c�p+���CEs�|( EQ�o  �7�SdB�AxT0 k� �\e�`e!2�$ !A&0    ��6 
   � < E�3�[�p+���CEo�|( EAxp  �/�SdB�AxT0 k� �Xd�\d!2�$ !A&0    ��6 
   � < E�4�S�p+�� DEk�|( EApq $�'�SdB�AxT0 k� �Pd�Td!2�$ !A&0    ��6 
   � < E�5�G�p+� DE�c�|( EAlr $	��SdB�AxT0 k� �Lc�Pc!2�$ !A&0    ��6 
   � < E�6�?�p/� EE�_�|( EAds $��SdB�AxT0 k� �Dc�Hc!2�$ !A&0    ��6 
   � < E�7�7�p/� FE�[�|( EA`t (��SdB�AxT0 k� �<c�@c!2�$ !A&0    ��6 
   � < Ea�8�/��/� FE�S�|( AXu (��SdB�AxT0 k� �0d�4d!2�$ !A&0    ��6 
   � < Ea�9�'��/� GE�O�|( APv ,���SdB�AxT0 k� �$e�(e!2�$ !A&0    ��6 
   � < Ea�;���/� GE�K�|( AHw ,��SdB�AxT0 k� �e�e!2�$ !A&0    ��6 
   � < Ea�<���/�  HE�C�|( ADw0��SdB�AxT0 k� �f�f!2�$ !A&0    ��6 
   � < Ea�=���, $IE�?�|( A<x0��SdB�ASxT0 k� �g�g!2�$ !A&0    �� 
   � < Ea�>���, $IE�7�|( A4y4�ۧSdB�ASxT0 k� ��h� h!2�$ !A&0    �� 
   � < 	A��?����, (IE�3�|( A,y4�ӧSdB�ASxT0 k� ��h��h!2�$ !A&0    �� 
   � < A�|A��0 ,JE�+�|( A(z8�ǨSdB�ASxT0 k� ��i��i!2�$ !A&0    �� 
   � < A�xB��0	 0JE'�|( A z�<￨SdB�ASxT0 k� ��i��i!2�$ !A&0    ��    � < A�tCߎ�0 0KE�|( A{�<﷨SdB�ASxT0 k� ��j��j!2�$ !A&0    ��    � < A�pD׏�0 4KE�|( A{�@ﯩSdB�ASxT0 k� ��j��j!2�$ !A&0    ��    � <��A�lEϏ�0 8KE�|( A{�@!里SdB�ASxT0 k� ��j��j!2�$ !A&0    ��    � <��A�hFǏ�0 8KE�|( A! |�D#SdB�ASxT0 k� ��j��j!2�$ !A&0    ��    � <��A�dG���0 <KE�|( A �|�D%SdB�ASxT0 k� ��k��k!2�$ !A&0    ��    � <��A�`H���0 <KE�|( A �|�H'SdB�ASxT0 k� ��k��k!2�$ !A&0    ��    � <��A�\I���0 @KE��|( A �|�H)SdB�ASxT0 k� ��k��k!2�$ !A&0    ��    � <��A�XJ���, @KJ��|( A �|�L+�w�SdB�A�xT0 k� ��k��k!2�$ !A&0    ��    � <��A�XK���, @KJ��|( A �|�P-�o�SdB�A�xT0 k� ��k��k!2�$ !A&0    ��    � <��A�TL���, @KJ��|( A �|�P/�g�SdB�A�xT0 k� ��k��k!2�$ !A&0    ��    � <��A�PM���,  DKJ��|( A �|�P1�_�SdB�A�xT0 k� ��k��k!2�$ !A&0    ��    � <��A�LN��(" DKJ��|( A �|�T3�W�SdB�A�xT0 k� ��k��k!2�$ !A&0    ��    � <��A�HOw��($ DKJ��|( A �|�T5�O�SdB�A�xT0 k� ��k��k!2�$ !A&0    ��    � <��A�DPo��$& DKJ��|( A �|�T7�G�SdB�A�xT0 k� �|j��j!2�$ !A&0    ��    � <��A�@Qg��$( DKJ��|( A0�{�T9�?�SdB�A�xT0 k� �ti�xi!2�$ !A&0    ��    � <��A�@R_�� * DKJ��|( A0�{�X;�7�SdB�A�xT0 k� �lh�ph!2�$ !A&0    ��    � <��A�<SS�� , DKJ��|( A0�{�X>�/�SdB�A�xT0 k� �dg�hg!2�$ !A&0    ��    � <��A�8TK��. bDKE��|( A0�z�X@�'�SdB3�A�xT0 k� �\g�`g!2�$ !A&0    ��    � <��A�4UC��0 bDKE��|( A0�z�XB��SdB3�A�xT0 k� �Tg�Xg!2�$ !A&0    ��    � <��A�4U;��2 bDKE��|( E�|z�XD��SdB3�A�xT0 k� �Lk�Pk!2�$ !A&0    ��    � <��A�0V�3��4 bDKE��|( E�ty�XF��SdB3�A�xT0 k� �Ho�Lo!2�$ !A&0    ��    � <��A�,W�'��5 bDKE��|( E�ly�TH��SdB3�A�xT0 k� �Dr�Hr!2�$ !A&0    ��    � <��A�(X���7 �DKE��|( E�dy�TJ�SdB3�A�xT0 k� �<s�@s!2�$ !A&0    ��    � <��A�(Y���9 �DKE{�|( E�Xx�TL��SdB3�A�xT0 k� �4t�8t!2�$ !A&0    ��    � <��A�$Y���; �DKEs�|( E�Px�TN�SdB3�A�xT0 k� �,u�0u!2�$ !A&0    ��    � <��A� ZQ���< �DKEk�|( E�Hx�PP�SdB3�A�xT0 k� � u�$u!2�$ !A&0    ��    � <��A� [P����> �DKE.c�|( E�<w�PQ�SdB3�A�xT0 k� �v�v!2�$ !A&0    ��    � <��A�\P���@ �DKE.[�|( A`4w�PS�SdB3�A�xT0 k� �v�v!2�$ !A&0    ��    � <��A�\P���ADKE.S�|( A`,w�LUߟSdB3�A�xT0 k� ��u��u!2�$ !A&0    ��    � <��A�]P���CDKE.K�|( A`$v�HWמSdB3�A�xT0 k� ��u��u!2�$ !A&0    ��    � <��A�^Pے��DDKE.?�|( A`v�HXӝSdB3�A�xT0 k� ��u��u!2�$ !A&0    ��    � <��A�_PӒ��FDKJN7�|( A`v�DZϜSdB3�A�xT0 k� ��t��t!2�$ !A&0    ��    � <��A�_Pǒ��GDKJN/�|( E@u�D\˛SdB3�
A�xT0 k� ��o��o!2�$ !A&0    ��    � <��A�`@����IRDKJN'�|( E@ u�@]ǚSdB3�
A�xT0 k� ��l��l!2�$ !A&0    ��    � <��A�a@����JRDKJN�|( EO�u�<_�ÙSdB3�
A�xT0 k� ��i��i!2�$ !A&0    ��    � <��A�a@����LRDKJN�|( EO�t�8`���SdB3�
A�xT0 k� ��g��g!2�$ !A&0    ��    � <��A�b@����MRDKJN�|(EO�t�8a���SdB3�	A�xT0 k� ��e��e!2�$ !A&0    ��    � <��A�c@����NRDKJN�|(EO�s�4c���SdB3�	A�xT0 k� ��d��d!2�$ !A&0    ��    � <��A� cГ���P�@KJM��|(EO�s00d���SdB3�A�xT0 k� ��b��b!2�$ !A&0    ��    � <��A� dЋ���Q�@KJ]��|(EO�r0,e���SdB3�A�xT0 k� ��a��a!2�$ !A&0    ��    � <��A��dЃ���S�@KJ]��|(A�r0(f���SdB3�A�xT0 k� ��`��`!2�$ !A&0    ��    � <��A��e�{���T�<KJ]��|(A�q0$g���SdB3�A�xT0 k� ��`��`!2�$ !A&0    ��    � <��A��f�s���U�<KJ]��|(A�p0 h���SdB3�A�xT0 k� �|_��_!2�$ !A&0    ��    � <��A��f�k���V�8KJ]��|(A�p0 i���SdB3�A�xT0 k� �p^�t^!2�$ !A&0    ��    � <��A��g�_�ߌX�4KE��|(A�o0j���SdB3�A�xT0 k� �d^�h^!2�$ !A&0    ��    � <��A��g�W�߄Y�4KE��|(EO�n�j���SdB3�A�xT0 k� �d\�h\!2�$ !A&0    ��    � <��A��h�O��|Z�0KE��|(EO�n�k���SdB3�A�xT0 k� �`[�d[!2�$ !A&0    ��    � <��A��h�G��t[�,KE��|(EO�m�l���SdB3�A�xT0 k� �\[�`[!2�$ !A&0    ��    � <��A��i�?��p\�(KE��|(EOxl�m���SdB3�A�xT0 k� �TZ�XZ!2�$ !A&0    ��    � <��A��j�7��p\�$KE��|(EOxl�m���SdB3�A�xT0 k� �LY�PY!2�$ !A&0    �    � <��A��j�+��h\� KE��|(EOpl� n���SdB3�A�xT0 k� �HY�LY!2�$ !A&0    ��    � <��A��k�#��`\�KE���|(EOhl��n���SdB3�A�xT0 k� �DY�HY!2�$ !A&0    ��    � <��A��k���X\�KE���|(EO`l��o���SdB3�A�xT0 k� �<Y�@Y!2�$ !A&0    ��    � <��A��l���P\�KE���|(AXl��o���SdB3�A�xT0 k� �,Y�0Y!2�$ !A&0    ��    � <��A��l���D\�KE���|(APl��o���SdB3�A�xT0 k� � Y�$Y!2�$ !A&0    ��    � <��A��m����<\�KE���|(AHl��p���SdB3�A�xT0 k� �Y�Y!2�$ !A&0    ��    � <��A��m����4\�KE���|(A@l��p���SdB3�A�xT0 k� �X�X!2�$ !A&0    ��    � <��A��n���,\KE���|(A@l��p���SdB3�A�xT0 k� � X�X!2�$ !A&0    ��    � <�A��n���$[�KE���|(A8l��p���SdB3�A�xT0 k� ��X��X!2�$ !A&0    ��    � <�}A��n�ߖ�[�KE����(A0l��p���SdB3�A�xT0 k� ��X��X!2�$ !A&0    ��    � <�{A��o�ח�[�KE}��(A(l��p���SdB3�A�xT0 k� ��X��X!2�$ !A&0    ��    � <�yA��o�˗�[�KE}{��(A k��p���SdB3�A�xT0 k� ��X��X!2�$ !A&0    ��    � <�wA��p�×� Z�KE}w��(Ak��p���SdB3�A�xT0 k� ��X��X!2�$ !A&0    ��    � <�uA��p�����Z�KE}w��(Aj��o�ÃSdB3�A�xT0 k� ��W��W!2�$ !A&0    ��    � <�sA��q�����Z�KE}s��(Aj��o�ǃSdB3�A�xT0 k� ��W��W!2�$ !A&0    ��    � <�qA��q�����Y�KD�o��(A.�i��o�ǂSdB3�A�xT0 k� ��V��V!2�$ !A&0    ��    � <�oA��q�����Y�KD�k��(	A.�i��n�˂SdB3�A�xT0 k� ��V��V!2�$ !A&0    ��    � <�mA��r�����Y�KD�k��(	A.�i��n�ςSdB3�A�xT0 k� ��U��U!2�$ !A&0    ��    � <�kA��r�����X�KD�g��(	A.�i��m�ӂSdB3�A�xT0 k� ��U��U!2�$ !A&0    ��    � <�iA��s����W�KD�c��(	A.�h��m�ӂSdB3�A�xT0 k� ��U��U!2�$ !A&0    ��    � <�gA��s���W�KD�_��(	A.�h��lׂSdB3�A�xT0 k� ��T��T!2�$ !A&0    ��    � <�eA��sw���V�KD�_��(	A.�g��lۂSdB3�A�xT0 k� ��T��T!2�$ !A&0    ��    � <�cA��tk���U�KD�[��(	A.�f��k߂SdB3�A�xT0 k� ��S��S!2�$ !A&0    ��    � <�aA��tc���T�KD�W��(	A.�f��j�SdB3�A�xT0 k� ��R��R!2�$ !A&0    ��    � <�_A��t[���S�KD�W��(	A.�e��i�SdB3�A�xT0 k� ��R��R!2�$ !A&0    ��    � <�]A��uS���R�KD�S��(	A.�d��i���dB3�A�xT0 k� �xQ�|Q!2�$ !A&0    ��    � <�[A��uK���Q�KD�O��(	A>�d��h���dB3�ASxT0 k� �pP�tP!2�$ !A&0    ��    � <�YA��v?���P|KD�O��(	A>�c��g���dB3�ASxT0 k� �hO�lO!2�$ !A&0    ��    � <�WA��v7���OtKD�K��(	A>�b��f����`B3�ASxT0 k� �`O�dO!2�$ !A&0    ��    � <�UA��v/���N�lKD�G��(	A>�a��e����`B3�ASxT0 k� �TN�XN!2�$ !A&0    ��    � <�SA��w'��xM�dKD�G��(	A>�`��d����`B3�ASxT0 k� �LM�PM!2�$ !A&0    ��    � <�QA��w��tK�\KD�C��(	A>x`��c���\B3�C�xT0 k� �DL�HL!2�$ !A&0    ��    � <�OA��w��lJ�TKD�C��(	A>p_��b���\B3�C�tT0 k� �<K�@K!2�$ !A&0    ��    � <�MA��w��hH�LKD�?��(	A>h^o�a���XB3�C�tT0 k� �4K�8K!2�$ !A&0    ��    � <�KA��x��`G�DKD�;��(	A>`]o�_���XB3�C�tT0 k� �,J�0J!2�$ !A&0    ��    � <�IA��x���\F�8KD�;��(	A>X\o�^���TB3�C�pT0 k� � I�$I!2�$ !A&0    ��    � <�GA��x��TD�0KD�7��(	A>P[o|]���TB3�C�lT0 k� �H�H!2�$ !A&0    ��    � <�FA��y��PC�(KD�7��(	AND[ox\���PB3�C�lT0 k� �G�G!2�$ !A&0    ��    � <�EA��yߚ�HA� KD�3��(	AN<Zox[���LB3�C�hT0 k� �D�D!2�$ !A&0    �    � <�IA��yך�D@�KD�3��(	AN4YotY�#��HB3�C�hT0 k� �$A�(A!2�$ !A&0    ��    � <�MA��zϚ�@?�KD�/��(	AN,XopX�'��HB3�C�dT0 k� �,>�0>!2�$ !A&0   ��    � <�QA��z�ǚ	�8>�KD�/��(	AN$WolW�+��DB3�C�`T0 k� �4;�8;!2�$ !A&0   ��    � <�UA��z	�4=��KD�+�|(	GnVodV�/��@B3�C�\T0 k� �@8�D8!2�$ !A&0   ��    � <�YA��z	�0;��KD�+�|(	GnVo`T�/��<B3�C�XT0 k� �H5�L5!2�$ !A&0   ��    � <�]A��{	�,:��KD�'�|(	GnUo\S�3��8B3�C�XT0 k� �P2�T2!2�$ !A&0   ��    � <�a                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��N ]�']'\ ` �� p�          � ڟ     p�� ڟ    ��                   �          ��     ���   0		!          �ݴm          ���'    �ݤ���     ���                 � ��        �     ���   8           ��Ip          �WZ    ��a��Wa&    ����                �         Ӡ  �  ���    	
	
�  	          Jt           ��b-     I�2���    "��   	            A�$                ���   (
	          �         .�H��     3��HZ�    �G�              ���$          ��     ���   X		          ��  ��	      B���    �����                              ���;              �  ���    0

 
2
 
            1�� � �
     V�y��     1h��x�8    j�             Z��          *��    ��`  
	           t�V  Q *	      j��p     t����dg    	Z          
 Z��          ��b     ��@ 8
          �      ~ �F      y    � �             # Z��         �      ��H   0	&          ?��  R R
     �����     ?���<�    6�              	
 Z��         	 ���   
  ��@  8
	           � ��     � �ݩ     � �ݩ                              ���n       
      �  ��@     

 0             UĐ � �	   �����     U�����I    ��	              s	 Z��         � �  (  ��`   @	                ��      �                                                                           �                               ��        ���          ��                                                                 �                          !o  ��        � ��     y �a    � � "                 x                j  �       �                              ��       �                      "                                                 �                          ��W���H��y�� �� �����          	        
 
  I   ��K #��       9$ �r@ :$  s@ :d s� ;� s` ˤ x� �� y  �D q` �D s� �d s����< ����J ����X ����  ����. ����< ����J ����X � � �t� �  u� �� �r@ �� s@ 
�< V� 
�< V� 
�\ W  
�< W� 
� W� 
�\ W� �� 0�  �� 0 �( 0�  �� 0�� �h 0� ���� � � }`���� � 
�| W����� � 
�< W� 
�� W� 
�| W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������� (�� Z  ������  
�fD
��L���"����D" � j  "  B   J jF�"   "�j  ���
��
��"     
�j ��   
 �
� �  �  
�      ��     �        p    ��     �            ��     �           � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �&!&      ��H �  ��        � � �  ��        �        ��        �        ��        �    ��    ��; ��        ��                         �$ (  ����                                    �                 ����              ���%��   (���� F �            2 Alexei Zhitnik      0:01                                                                        7  5     � �
"�; �
� �7K. �O K6 �(C �= C |kV k\ � �	k` � �
C C"! �c� �c�" � c� �k�) �k�! �k�1 �k�1 � k�1 � k�B �cjE � cr= � cs= x � � w � � cc~ � { c� � `J�= x J�M �"� � � "� � v � � v!
� � �""�< � #"�N r$"�8 r%*�G �&"� � � '"� � v(� � v)
� �6  *�6  *�> )�x � -*Fx.*8x.  *Gx0*8x.  *Gx � 2*Fx3*8x.  *Gx>  *Ax �  *As � 7*Os �  *Ks �  *Ks< )�s@ )�s �  *GZ �  *HZ � >)�B �  *HZ                                                                                                                                                                                                                         �� R         �     @ 
        A     k P E m  ���� @               
 �������������������������������������� ���������	�
��������                                                                                          ��    ���   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, ;� < F�  ]� g@���@� @��@������ ��~� ����                                                                                                                                                                                                                                                                                                              t@��A�                                                                                                                                                                                                                                         d    +    ��   R�J    
  "�  	                           ������������������������������������������������������                                                                                                                                         �    �      ��              �     �          	 	 
  	 	 	  ��  ������ ����������������������������������� � ���������������������������� ��������������������� ������� ����������������������� ������� ���������������� �������������������������� ��������������� �������� �� ��� �������� �� �           �                    �   " 3     �  :�J      �                             ������������������������������������������������������                                                                                                                                 �    �    �        e      �� u       �          
     �������������������� �� �������������� �������������������������������������������� ���������������������  ������������ ������������� �� �� ��������    ��������������� ��� � ����� ��������� ����������������������������������� ��� ��������� ��           x                                                                                                                                                                                                                                                                                       	                   �             


             �  }�         ������������  '�������������  +&   $����������������������������  N�����    ����������������������������                     R�                           'x  R�  'x                        ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""  L @               
                  � ��T� �r@                                                                                                                                                                                                                                                                                      )n)n
  1n)�        m            m            `            k      l                                                                                                                                                                                                                                                                                                                                                                        j                               > �  >�  @�  J�  C#�  J`�  ������̞����������]�F2��̎���� �������        <        �� G         
 
 �   & AG� �  O   
           �:�                                                                                                                                                                                                                                                                                                                                      J K    �     	                !��                                                                                                                                                                                                                            Y     �� �~ ��      �� D 
   
 ��  ������ ����������������������������������� � ���������������������������� ��������������������� ������� ����������������������� ������� ���������������� �������������������������� ��������������� �������� �� ��� �������� �� ��������������������� �� �������������� �������������������������������������������� ���������������������  ������������ ������������� �� �� ��������    ��������������� ��� � ����� ��������� ����������������������������������� ��� ��������� ��   �� �     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    >   !   I   !                          D     �  ����������      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$ ^h  ��   p   	 ��     �           �� �   6   
���(��   �   �  x���� ��  x  � ��� ��  � ��� n 
a�     �      �=  r@ 9$ ��  r@ 9$ �$ "  ��"        �   d   r���� e�����   g��� 	  �     f ^�          �� L (      r      ��Nz���2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                                      ���        ������������������ݭ�        �������ݪ������������        �               �                            �             �   �  ��  ͬ 
������������-Ѭ�����!-��!-��-̬����������!�"�-�����!��-�������������-�-��!����������-��,���,����-���-����ܭ��ܭ���� ̪� ʡ  ��  ��   �� ���
���ڪ��            !�-��!���ݪ���         
����-�����ͬ��ͬ��Ѭ̭Ѭ��ͪ���-�����������������̭�������������ʬ���         ��  �   �   �   �                                                                        �     Ѭ�� Ѫ�  Ѫ   �   
            ��ʡ̬Ѡ�Ѡ ݠ  �                                                                         �    wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "" "  """ ""   "! " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """               "  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """ ""   "! " ""  !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                   �   �                      �������  ���    �                    ��� ���� �� �   ��  ��  ��  �  �   ��  ��      � ���� ��   � � �                                                                                                                                                         	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                                   ��                  �                        ���� ��� ����            �   �   �   D   E�  U�  UO                         "  "  "                                                                                                                                                                �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        T   S   C   3   30  30  ;�  ��  ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �   �  �  �� �� �   �                            � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��   �  �   �   ��  �            ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    ���� �  ��     �                                    �  �� �                         ����     �   �  �  �  ��  �   �                                                                                                        �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����            �  �  ��  �   �   �        �   ��  ��  ��  �  �   ��  ��                                                                                                                                                                       �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �   �"!�����                            �  �� Ș ��  ��  �                              �  ��    �       �   �   �                                                                                                                                                                           ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                      ��� ���� ��                  ���                                                                                                                                                                                                 
   �   �  ��  �� ������-�� "��  �  
�  �C 
UU US �UD TE0 �� 
�� ʐ �  ̻  "�  "   " �� ����   �  �˰ ̻� �ݰ �w� ��� ����������˹�̹���ڙ��ٻ��ݰ̻� ˘  ��  3D  TD� 340 340 3D0 30 
��  ��  "/  "/  �� ���� �    ��                  "      �           �  �   �   ��  �             ��  ��  �                            �   �    �   �       �   �   �                .      �   "   "   "  �  �   �   ���                                                                                                                                                                                                           �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                /���"/�  ��                    �                                                                            �               �  �  ��  �   �   �                               ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                            �  	�  ˹ ˹ �̹ ��� ̽� ̽�̽�	�ͺ������J�CT�T UJ� UT� EU� T� J�  ��  ��  ʩ ̰ �  "" "" ""    ��   ��  ��  ��  �w  �p  ��  ��  ��  ̰  Ȱ  ��  ��  ��  ��  "�  0"� 3 � 30�C0 �C  Ƞ  ��  ��  ݻ ��"/""""""/"��� ��� ��             �� ������ ����  �   �  �   �  �     �                                       ��  "   /�  �  �              � ��         �� �� �� g} �� vw                     ��  ��  ��� ���                                                                                                                                                                                                                     �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                     �                             �   �   �   �   �   �                                                                                                                                       �  ��� ݻ� g�� bm� ggz�'w���������������˛������ˊۼ�����˻������H�DH�@U�DPT�E X�T H�P H�@ Ȥ� ̻� ˘ "�� � ���/�"" �""/���               �   �                                                     �  �                      � �                       ���           �                      �  �  �          ����  �   �             ����                         � "            � "�",�"+� ",                       "  .���"    �     �                              �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""wwwwwwwwwwwww""""wwwwwwwGwqGwGwDGwG""""wwwwwwqAqwAwG""""wwwwwwwwDDwwwwwwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwqDDDG""""wwwwwqqADAqq""""wwwwwwqwwwqwqwq""""wwwwqDDDwGq"""$www4ww4Gw4DGw4www4ww4wwwwwwwwwwtwww333DDDGwGGwqwDDwtwwww3333DDDDwGtqGwADqDGwDwwww3333DDDDwwqwwwwDwwDGwwwwww3333DDDDADAGqGqtGwDwwww3333DDDDGqGqGqGqtGwDwwww3333DDDDGqqqwwtDDwwww3333DDDDDDqwqqqwAwtDGwwww3333DDDDwqwqwGqDDGwwwww3333DDDDDGwAwwwwDDtDwwww3333DDDDww4Gw4Gw4Gw4Dww4www43334DDDD"""������������������""""������������������������""""��������������������""""������DDM�D��""""�������MM�M�M""""��������DD�A��""""�������MAA�MA""""��������AA�A""""����������M�MA""""������������M���M���M���"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUQUUQUUUUUUQUUUUUUUU3333DDDDUUUUDEEDDTEUUUU3333DDDDAEAEQQUDTDUUUU3333DDDDQUQUQDUDDUUUU3333DDDDAADAUAUEDUTUUUU3333DDDDADAEAQAUEDUTUUUU3333DDDDUDUQEUQUUQUEUDUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=LL����������D����3333DDDD    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����������A������ x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx""""�������I�I������ w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww""""�������I��D���I�������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(�D�M�D���M������3333DDDD �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""�����AMAD������ M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M""""������������������ � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
"�; �
� �7K. �O K6 �(C �= C |	kVk\ � �	k` � �
C C"! �c� �c�" � c� �k�) �k�! �k�1 �k�1 � k�1 � k�B �cjE � cr= � cs= x � � w � � cc~ � { c� � `J�= x J�M �"� � � "� � v � � v!
� � �""�< � #"�N r$"�8 r%*�G �&"� � � '"� � v(� � v)
� �6  *�6  *�> )�x � -*Fx.*8x.  *Gx0*8x.  *Gx � 2*Fx3*8x.  *Gx>  *Ax �  *As � 7*Os �  *Ks �  *Ks< )�s@ )�s �  *GZ �  *HZ � >)�B �  *HZ3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������ �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������=�N�K�U�X�K�T��0�R�K�[�X�_� � � � � � �-�1�B�����������������������������������������!��;�U�H�K�X�Z��;�K�O�I�N�K�R� � � � � � �-�1�B�������������������������������������������+�R�K�^�K�O��C�N�O�Z�T�O�Q� � � � � � �6�+� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������-�1�B� ��"�������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������6�+� � ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            