GST@�                                                           @h�                                                                ��             :`  2�������ʱ���������    ����        ��      #    ����                                d8<n    �  ?     F����  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    "�j��,  " ��
  �                                                                               ����������������������������������      ��    bb QQb  114 44c c   c      		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������=  0b  4  11                                         �  �  �  �                  F  
1          = �����������������������������������������������������������������������������                                ��  �       w�   @  #   �   �                          �                                                     'w w  )n)n1n  
1F    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    E�_���B�T0�(O-0W�$��E��tQ;�;��-TQs�T0 k� ��]��]%�0d  U8D"!  ��O    � 8�8E�_���B�X0�0N-0W�$��E��vQ;�;��,TOs�T0 k� ��^��^%�0d  U8D"!  ��O    � 9�9E�^��B�\0�4M-0X� ��E��wQ;�:��,TNs�T0 k� ��`��`%�0d  U8D"!  ��G    � :�:E��]��B�\0�<M-0Y� �#�E��yQ;�:��,TMs�T0 k� <�d� d%�0d  U8D"!  ��G    � ;�;E��\��B�d1�HL-0Z� }'�E��{Q;�9��,XJs�T0 k� =h�h%�0d  U8D"!  ��G    � <�<E��[��B�h1	LK-0Z� }+�E� |Q;�8��,XIs�T0 k� =j�j%�0d  U8D"!  ��G    � <�=E��Z�'�B�l1	TK-0[� }/�E�~Q;�8��,XHs�T0 k� =l� l%�0d  U8D"!  ��G    � <�>E��Z�/�B�p1	XK-0[� }3�E�Q;�7��,\Fs�T0 k� �$m�(m%�0d  U8D"!  ��G    � <�?E��X�?�B�x1	dJ0\� }7�E��Q;�6��,`Ds�T0 k� �,o�0o%�0d  U8D"!  ��G    � <�@E��W�G�B�x1	hJ0]� };�E��Q;�6��,�`Bs�T0 k� �4o�8o%�0d  U8D"!  ��G    � <�AE��V�O�B�|1	,lJ0]� };�E� �Q;�5��,�dAs�T0 k� �8o�<o%�0d  U8D"!  ��G    � <�BE��U�W�E��1	,tI4^� }?�E�$�Q;�5��,�d@s�T0 k� �<n�@n%�0d  U8D"!  ��G    � <�BE��T�_�E��1	,xI4^� }?�E�,�Q;�4��+�h>s�T0 k� �Dn�Hn%�0d  U8D"!  ��G    � <�BE,�R�o�E��1	,�I8_� }G�E�4Q;�4��+�l<s�T0 k� �@l�Dl%�0d  U8D"!  ��G    � <�BE,�Q�w�E��1	�I8_� mG�E�<~Q;�3��+�p;s�T0 k� �@k�Dk%�0d  U8D"!  ��G    � <�BE,�P��E��2	�I<`� mK�E�@~Q;�3��*�t9s�T0 k� �@i�Di%�0d  U8D"!  ��G    � <�BE-O���E��2	�I<`� mK�E�D}Q;�2��*�t8s�T0 k� �@h�Dh%�0d  U8D"!  ��G    � <�BE-N���E~�2	�I�@`� mO�E�H|Q;�2��*�x7s�T0 k� �Df�Hf%�0d  U8D"!  ��G    � <�BE-M���E~�3	�I�Da� mO�E�P|Q;�2��)�|6s�T0 k� �De�He%�0d  U8D"!  ��G    � <�BE-K���E~�3	,�I�Hb� mS�E�XzQ;�1��(��3s�T0 k� �Ld�Pd%�0d  U8D"!  ��G    � <�BE$J���E~�4	,�I�Lb� mS�E�\yQ;�0(��2s�T0 k� �Pc�Tc%�0d  U8D"!  ��G    � <�BE(I���E~�4	,�I�Pb� mS�E�`xQ;�0'��1s�T0 k� �Tb�Xb%�0d  U8D"!  ��G    � <�BE0H�ÈE~�5	,�I�Tc� mS�E�hwQ;�0'��0s�T0 k� �Xa�\a%�0d  U8D"!  ��G    � <�BE8G�ˈE~�6	,�I�Xc� mS�E�lvQ;�/&��/s�T0 k� �\`�``%�0d  U8D"!  ��G    � <�BE<F�ӉE~�6	�I�\c� ]S�E�puQ;�/%��.s�T0 k� �\a�`a%�0d  U8D"!  ��G    � <�BELD��En�8	�I�dd� ]S�E�puQ< . $��-s�T0 k� �``�d`%�0d  U8D"!  �G    � <�CEPC��En�8	�I�dd� ]S�E�tuQ< .$#��,s�T0 k� �da�ha%�0d  U8D"!  ��G    � <�DEXB��En�9	�I�hc� ]S�E�xtQ< -("��+s�T0 k� �db�hb%�0d  U8D"!  ��G    � <�DE`A���En�:	,�I�lc� ]S�E=|tQ< -0!��*s�T0 k� �l`�p`%�0d  U8D"!  ��G    � <�EEh@��En�;	,�I�pc� ]O�E=�sQ< -4 ��*s�T0 k� �t_�x_%�0d  U8D"!  ��G    � <�FEt>��En�=	,�I�|b� ]O�E=�rQL ,o<��)s�T0 k� ��^��^%�0d  U8D"!  ��G    � <�GE�|=��En�=	,�I��b� ]K�E=�rQL ,o@��(s�T0 k� ��]��]%�0d  U8D"!  ��G    � <�HE��=��En�>	�I��b� ]K�E=�rQL +oD��(!��T0 k� ��]��]%�0d  U8D"!  ��G    � <�IE��<�'�E^�?	�I��a� ]G�E=�qQL +oH��'!��T0 k� ��\��\%�0d  U8D"!  ��G    � <�JE��;�+�E^�@	�I��a� ]C�E=�qQL+oH��'!��T0 k� ��\��\%�0d  U8D"!  ��G    � <�KE��:�3�E^�A	�I��`� MC�E=�pQL+oL��'!��T0 k� ��[��[%�0d  U8D"!  ��G    � <�KE��9�?�E^�C	,�I�_� M?~E=�oQL*oT��'!��T0 k� ��Z��Z%�0d  U8D"!  ��G    � <�LE��9�C�C��D	,�I�_� M;E=�oU*?T��&!��T0 k� ��Y��Y%�0d  U8D"!  ��G    � <�ME��8�K�C��E	,�I�^� M7E=�nU)?X��&!��T0 k� ��X��X%�0d  U8D"!  ��G    � <�NE��8�O�C��F	,�I�]� M3E=�nU)?X��&!��T0 k� ��X��X%�0d  U8D"!  ��G    � <�OE��8�S�C��F	,�I�]� �/�E-�mU)?\��'!��T0 k� ��Y��Y%�0d  U8D"!  ��G    � <�PE}�7�W�C��G �I-�\� �/�E-�lU(?\��'!��T0 k� ��Y��Y%�0d  U8D"!  ��G    � <�QE}�7�[�C��H �I-�\� �+�E-�lU(?`��'s�T0 k� ��Y��Y%�0d  U8D"!  ��G    � <�RE}�7�_�C��I �I-�[� �'�E-�lU(?`� 's�T0 k� ��Z��Z%�0d  U8D"!  ��G    � <�SE}�7�g�C��J �I-�Z� ��E-�jU'?d�(s�T0 k� ��Y��Y%�0d  U8D"!  ��G    � <�TE}�7�k�C��K �I-�Y� ��E-�i@'?d
�(s�T0 k� ��X��X%�0d  U8D"!  ��    � <�UE}�7�o�C��L �I�Y� ��E-�i@'?d�(s�T0 k� ��X��X%�0d  U8D"!  ��    � <�VE}�7�s�C��M �I�X� ��E-�i@'?d�)s�T0 k� ��X��X%�0d  U8D"!  ��    � <�WE~7�s�C��M �I�W� ��E-�h@&Od�)s�T0 k� ��W��W%�0d  U8D"!  ��    � <�XD�7�w�C��N �I�W� ��E-�g@&Od�)s�T0 k� ��V��V%�0d  U8D"!  ��    � <�YD�7�w�C��O �I�V� ��E-�fE�&Od�*s�T0 k� ��U��U%�0d  U8D"!  ��    � <�ZD�8�{�C��O �I�U� ��E�eE�%Od�*s�T0 k� ��Y��Y%�0d  U8D"!  ��    � <�[D�$8�{�C��Q �I�T�$���E�dE�%og��+!��T0 k� � \�\%�0d  U8D"!  ��    � <�\E~,9��C��R �I�T�$��E�cE�$og��+!��T0 k� �^�^%�0d  U8D"!  ��    � <�]E~09��E^�R �I�S�$��E bE�$og��+!��T0 k� �_�_%�0d  U8D"!  ��    � <�^E~8:��E^�S �I�S�$	|�EaB�#og��,!��T0 k� �`�`%�0d  U8D"!  ��    � <�_E~<:��E^�S �I�R�$	|�EaB�"og��,!��T0 k� �a� a%�0d  U8D"!  ��'    � <�`E~@;��E^�T �I�R�$	|�E`B� "oc��,!��T0 k� �$b�(b%�0d  U8D"!  ��'    � <�aEnL<��EޜU �I�R�$	|ۏE ^B�$!oc��-!��T0 k� �0a�4a%�0d  U8D"!  �'    � <�aEnP=^�EޔV �I �Q�$LאE(^E( oc��-!��T0 k� �8a�<a%�0d  U8D"!  �'    � <�aEnX=^�EސW �I �Q�$LӑE,]E( o_��-!��T0 k� �@a�Da%�0d  U8D"!  ��'    � <�aEn\>^{�EތW �I �Q�$L˒E4\E, o_��.s�T0 k� �H`�L`%�0d  U8D"!  ��'    � <�aEn`?^{�EވX �I �P�$LǒE�<[E0 _[��.s�T0 k� �Lc�Pc%�0d  U8D"!  ��'    � <�aA�d?^{�E�Y �I �P�$LÓE�D[E4 _[��.s�T0 k� �Tf�Xf%�0d  U8D"!  ��'    � <�aA�p@^{�E�Y �I �P�$L��E�D[E<_W��/s�T0 k� �dd�hd%�0d  U8D"!  �/    � <�aA�tA^{�E�Z �I �O�$L��E�D[E<_S��/s�T0 k� �lg�pg%�0d  U8D"!  ��"    � <�aA�xB^{�E�Z �I �O�$L��R�@[E�@_O��/s�T0 k� �li�pi%�0d  U8D"!  ��"    � <�aA�|B^{�P��[ �I �O�$L��R�@[E�D_O��0s�T0 k� �hj�lj%�0d  U8D"!  ��"    � <�aA��C^{�P��[ �I �O�$<��R�@[E�H_K��0s�T0 k� �`k�dk%�0d  U8D"!  ��"    � <�aA��C^{�P��\ �I �N�$<��R�<[E�P_G��0s�T0 k� �\k�`k%�0d  U8D"!  ��"    � <�aA��D^{�P��\ �I �N�$<��R�<[E�T_C��0s�T0 k� �\l�`l%�0d  U8D"!  ��"    � <�aA��D^{�P��] �I �N�$<��R�<[D�X_?��1s�T0 k� �\l�`l%�0d  U8D"!  ��"    � <�aA��E^{�P�|] �I  N�$<��R�8[D�\_;��1s�T0 k� �Po�To%�0d  U8D"!  ��"    � <�aA��E^{�P�|^ �I  N�$<��R�8[D�`O7�� 1s�T0 k� �Hq�Lq%�0d  U8D"!  ��"    � <�aA��F^{�P�|_ �I  M�$<��R�8[D�dO3��1s�T0 k� �Ds�Hs%�0d  U8D"!  ��"    � <�aA��F^w�P�|_ �I  M�$<��R�8[D�hO/��2s�T0 k� �@t�Dt%�0d  U8D"!  ��"    � <�aA��G^w�P�x` �I M�$<��R�4[D�lO+��2s�T0 k� �8v�<v%�0d  U8D"!  ��"    � <�aA��G^w�P�x` �I M�$<{�R�4[D�tO'��2s�T0 k� �4w�8w%�0d  U8D"!  ��"    � <�aA��H^w�P�xa �I M�$Lw�R�4[D�xO#��2s�T0 k� �4x�8x%�0d  U8D"!  ��"    � <�aA��H^w�P�xa �I L�$Ls�R�0[D�|O��3s�T0 k� �<v�@v%�0d  U8D"!  ��"    � <�aA��H^w�P�ta �I L�$Lo�R�0[D����3s�T0 k� �<u�@u%�0d  U8D"!  ��"    � <�aA��I^w�P�tb �I L�$Lk�R�0[D� ���3s�T0 k� �@t�Dt%�0d  U8D"!  ��"    � <�aA��I^w�P�tb �I L�$Lg�R�0\D� ���3s�T0 k� �Dt�Ht%�0d  U8D"!  ��"    � <�aA��J^w�P�tc �I L�$<c�R�,\D� ���3s�T0 k� �Dt�Ht%�0d  U8D"!  ��"    � <�aA��J^w�E�tc �I K�$<_�R�,\D�!���4s�T0 k� �Dv�Hv%�0d  U8D"!  ��"    � <�aA��K^w�E�pd �I K�$<[�R�,\D�!���4s�T0 k� �Hw�Lw%�0d  U8D"!  ��"    � <�aA��K^w�E�pd �I K�$<W�R�,\D�"����4s�T0 k� �Lx�Px%�0d  U8D"!  ��"    � <�aA��K^w�E�pe �I K�$<W�R�,\D�"����4s�T0 k� �Lx�Px%�0d  U8D"!  ��"    � <�aA��L^w�E�lf �I K�$�S�R�(\D�#����4s�T0 k� �Hy�Ly%�0d  U8D"!  ��"    � <�aA��L^w�E�lf �I K�$�O�R�(\D�#����5s�T0 k� �Tz�Xz%�0d  U8D"!  ��"    � <�aA��M^w�E�lg �I J�$�K�R�(\D�$����5s�T0 k� �\z�`z%�0d  U8D"!  ��"    � <�aA��M^w�E�hh �I J�$�G�R�(\D��%����5s�T0 k� �d{�h{%�0d  U8D"!  ��"    � <�aA��M^w�E�hh �I J�$�C�R�$\D��%����5s�T0 k� �h|�l|%�0d  U8D"!  ��"    � <�aA��N^w�E�hi �I J�$
�?�R�$\D��&����5s�T0 k� �h}�l}%�0d  U8D"!  ��"    � <�aA��N^s�E�dj �I J�$
�;�R�$\D��'����6s�T0 k� �l}�p}%�0d  U8D"!  ��"    � <�aA��N^s�E�dk �I J�$
�;�R�$\D��'����6s�T0 k� �p~�t~%�0d  U8D"!  ��"    � <�aA��O^s�E�dk �I I�$
�7�R�$\D��(����6s�T0 k� �p�t%�0d  U8D"!  ��"    � <�aA��O^s�E�`l �I I�$
�3�R� \D��)N���6s�T0 k� �p��t�%�0d  U8D"!  ��"    � <�aA��O^s�E�`m �I I�$
�/�R� \D��*N���6s�T0 k� �p��t�%�0d  U8D"!  ��"    � <�aA��P^s�E�`n �I I�$
�+�R� \D��+N���x6s�T0 k� �l��p�%�0d  U8D"!  ��"    � <�aA��P^s�E�\o �I I�$
�+�R� \D��,N���t7s�T0 k� �l��p�%�0d  U8D"!  ��"    � <�aA��P^s�E�\p �I I�$	�'�R� \D��,N���l7s�T0 k� �l��p�%�0d  U8D"!  ��"    � <�aA��Q^s�E�\p �I  I�$	�#�R� \E ->���d7s�T0 k� �h��l�%�0d  U8D"!  ��"    � <�aA��Q^s�E�Xq �I  H�$	�#�R�\E.>���\7s�T0 k� �h��l�%�0d  U8D"!  ��"    � <�aA��Q^o�A�Xq �I  H�$	��R�\E/>���X7s�T0 k� �`��d�%�0d  U8D"!  ��"    � <�aA� R^k�A�Xq �I  H�$	��R�\E0>���P7s�T0 k� �X��\�%�0d  U8D"!  ��"    � <�aA� R^k�A�Tq �I  H�$	��R�\E1>���H7s�T0 k� �P�T%�0d  U8D"!  ��"    � <�aA�R^g�A�Tp �I $H�$	��R�\E� 2N���@8s�T0 k� �L~�P~%�0d  U8D"!  ��"    � <�aA�S^g�A�Tp �I $H�$	��R�\E�(3N��88s�T0 k� �H}�L}%�0d  U8D"!  ��"    � <�aA�S^c�A�Tp �I $H�$	��R�\E�04N��08s�T0 k� �D|�H|%�0d  U8D"!  ��"    � <�aA�S^c�A�Pp �I $H�$��R�]E�45N��,8s�T0 k� �D|�H|%�0d  U8D"!  ��"    � <�aA�S^_�A�Po �I $G�$��R�]E�<6N��$8s�T0 k� �D|�H|%�0d  U8D"!  ��"    � <�aA�T^_�A�Po �I (G�$��R�]E�D8N��8s�T0 k� �D|�H|%�0d  U8D"!  ��"    � <�aA�T^[�A�Po �I (G�$��R�]E�H9N��8s�T0 k� �@|�D|%�0d  U8D"!  ��"    � <�aA�T^[�A�Lo �I (G�$��R�]E}P:N��9s�T0 k� �@{�D{%�0d  U8D"!  ��"    � <�aA�U^W�A�Ln �I (G�$��R�]E}X;^��9s�T0 k� �@{�D{%�0d  U8D"!  ��"    � <�aA�U^W�A�Ln �I (G�$���R�]E}\<^�� 9s�T0 k� �@{�D{%�0d  U8D"!  ��"   � <�aA�U^S�A�Ln �I (G�$���R�]E}d>^���9s�T0 k� �<{�@{%�0d  U8D"!  ��"    � <�aA�U^S�A�Hn �I ,G�$���R�]E}h?^���9s�T0 k� �<z�@z%�0d  U8D"!  ��"    � <�aA� V^O�A�Hn �I ,G�$���R�]E}p@^���9s�T0 k� �<z�@z%�0d  U8D"!  ��"    � <�aA� V^O�A�Hm �I ,F�$���R�]E}xB^���9s�T0 k� �<z�@z%�0d  U8D"!  ��"    � <�aA�$V^O�A�Hm �I ,F�$���R�]E}|C^��9s�T0 k� �<z�@z%�0d  U8D"!  ��"    � <�aA�$V^K�A�Hm �I ,F�$���R�]E}�D^�.�:s�T0 k� �8z�<z%�0d  U8D"!  ��"    � <�aA�(V^K�A�Dm �I ,F�$���R�]E}�F^{�.�:s�T0 k� �8y�<y%�0d  U8D"!  ��"    � <�aA�(W^G�A�Dm �I 0F�$���R�]E}�G^{�.�:s�T0 k� �8y�<y%�0d  U8D"!  ��"    � <�aA�,W^G�A�Dm �I 0F�$���R�]E}�I^w�.�:s�T0 k� �8y�<y%�0d  U8D"!  ��"    � <�aA�,W^G�A�Dl �I 0F�$���R�]E}�Jnw�.�:s�T0 k� �8y�<y%�0d  U8D"!  ��"    � <�aA�0W^C�A�Dl �I 0F�$���R�]Em�Lns�.�:s�T0 k� �4y�8y%�0d  U8D"!  ��"    � <�aA�0X^C�A�@l �I 0F�$���R�]Em�Mns�.�:s�T0 k� �4y�8y%�0d  U8D"!  ��"    � <�aA�0X^?�A�@l �I 0F�$���R�]Em�Ono�.�:s�T0 k� �4x�8x%�0d  U8D"!  ��"    � <�aA�4X^?�A�@l �I 0F�$���R�]Em�Pno�.�:s�T0 k� �4x�8x%�0d  U8D"!  ��"    � <�aA�4X^?�A�@k �I 4F�$���R�]Em�R�k�.�;s�T0 k� �4x�8x%�0d  U8D"!  ��"    � <�aA�8X^;�A�@k �I 4E�$���R�]Em�T�g�.�;s�T0 k� �0x�4x%�0d  U8D"!  ��"    � <�aA�8Y^;�A�<k �I 4E�$���R�]Em�U�g�.�;s�T0 k� �0x�4x%�0d  U8D"!  ��"    � <�aA�<Y^;�A�<k �I 4E�$���R�]Em�W�c�.�;s�T0 k� �0x�4x%�0d  U8D"!  ��"   � <�aA�<Y^7�A�<k �I 4E�$���R�]Em�X�c�.�;s�T0 k� �0w�4w%�0d  U8D"!  ��"    � <�aA�<Y^7�A�<k �I 4E�$���R�]Em�Z�_�.�;s�T0 k� �0w�4w%�0d  U8D"!  ��"    � <�aA�@Y^3�A�<k �I 4E�$���R�]Em�\�_�.�;s�T0 k� �,w�0w%�0d  U8D"!  ��"    � <�aA�@Z^3�A�<j �I 8E�$���R�]Em�\�[�.�;s�T0 k� �,w�0w%�0d  U8D"!  ��"    � <�aA�@Z^3�A�8j �I 8E�$���R�]E]�^�[�.�;s�T0 k� �,w�0w%�0d  U8D"!  ��"    � <�aA�DZ^3�A�8j �I 8E�$���R�]E]�`�[�.�;s�T0 k� �,w�0w%�0d  U8D"!  ��"    � <�aA�DZ^/�A�8j �I 8E�$���R�]E]�a�W�.|;s�T0 k� �,w�0w%�0d  U8D"!  ��"    � <�aA�HZ^/�A�8j �I 8E�$���R�]E]�c�W�.x<s�T0 k� �,v�0v%�0d  U8D"!  ��"    � <�aA�HZ^/�A�8j �I 8E�$���R�]E]�d�S�.t<s�T0 k� �,v�0v%�0d  U8D"!  ��"    � <�aA�H[^+�A�8j �I 8E�$���R�]E]�f�S�.p<s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�L[^+�A�8j �I 8D�$���R�]E]�gO�.p<s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�L[^+�A�4j �I 8E�$���R�]E]�iO�.l<s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�L[^'�A�4j �I 8E�$���R�]E]�jK�.l;s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�P[^'�A�4k �I 8E�$���R�]E]�lK�.h;s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�P[^'�A�4k �I 4E�$ ���R�]E]�mK�.h;s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�P\^'�A�4k �I 4E�$ ���R�]EM�nG�.h;s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�T\^#�A�4k �I 4F�$ ���R�]EM�pG�.d;s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�T\^#�A�4k �I 0F�$ ���R�\EM�qC�.d;s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�T\^#�A�4k �I 0F�$ ���R�\EM�rC�.`:s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�T\^#�A�4k �I 0F�$ k��R�\EM�s@ .`:s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�X\^�A�4k �I 0F�$ k��R�\EM�t<.\:s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�X\^�A�4k �I 0F�$ k��R�\EM�u<.\:s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�X]^�A�4k �I ,F�$ k��R�\EM�v<.X:s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�\]^�A�4k �I ,G�$ k��R�\EM�w8.X:s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�\]^�A�4k �I ,G�$ ��R�\EM�x8.X:s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�\]^�A�4k �I ,G�$ ��R�\EM�y8.T9s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�\]^�A�4k �I (G�$ ��R�\E=�y4.T9s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�`]^�A�4k �I (G�$ ��R�\E=�z4.P9s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�`]^�A�4k �I (G�$ ��R�[E=�{4P9s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�`^^�A�4k �I (G�$���R�[E=�{0	P9s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�`^^�A�4k �I (H�$���R�[E=�|0
L9s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�d^^�A�4k �I $H�$���R�[Kݨ|0L9s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�d^^�A�4k �I $H�$���R� [Kݨ},L8s�T0 k� �(v�,v%�0d  U8D"!  ��"   � <�aA�d^^�A�4k �I $H�$���R� [Kݤ},H8s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�d^^�A�4k �I $H�$���R� [Kݤ~,�H8s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�h^^�A�4k �I $H�$���R� [Kݠ~(�D8s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�h^^�A�4k �I  H�$���R� [Kݠ(�D8s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�h^^�A�4k �I  H�$���R� [Kݜ(�@8s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�h_^�A�4k �I  I�$���R� [Kݜ�(�@8s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�l_^�A�4k �I  I�$���R� [Kݘ$�<8s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�l_^�A�4k �I  I�$���R� ZKݘ$�87s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�l_^�A�4k �I I�$���R�$ZKݔ$�87s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�l_^�A�4k �I I�$���R�$ZKݔ$�47s�T0 k� �(v�,v%�0d  U8D"!  ��"    � <�aA�l_^�A�4k �I I�$���R�$ZKݐ~ N07s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�p_^�A�4k �I I�$���R�$ZK�~ N,7s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�p_^�A�4k �I I�$���S$ZK�~ N,7s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�p_^�A�4k �I I�$���S$ZK�~ N(7s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�p_^�A�4k �I J�$���S$ZK�}N$7s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�p`^�A�4k �I J�$���S$ZK�}N 7s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�t`^�A�4k �I J�$���S$ZK�}N8s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�t`^�A�4k �I J�$���S$ZK�}N8s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�t`^�A�4k �I J�$���S$ZK�}�N8s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�t`^�A�4k �I J�$���S(ZK�|�N8s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�t`^�A�4k �I J�$���S(ZK�|��9s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�t`^�A�4k �I J�$���U�(ZK�|��9s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�x`^�A�4k �I J�$���U�(ZK�|��9s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�x`^�A�4k �I J�$���U�(ZK�||�� :s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�x`^�A�4k �I K�$��U�(ZK�|{���:s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�x`^�A�4k �I K�$��U�(ZK�|{���:s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�xa^�A�4k �I K�$��U�(ZK�x{���;s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�xa^�A�4k �I K�$��U�(ZK�x{���;s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�|a^�A�4k �I K�$��U�(ZK�x{���<s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�|a^�A�4k �I K�$��U�(ZK�tz���=s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�|a^�A�4k �I K�$��BN(ZK�tz���=s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�|a]��A�4k �I K�$��BN,ZK�tz� ��>s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�|a]��A�4k �I K�$��BN,ZK�pz�!��>s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�|a]��A�4k �I K�$��BN,ZK�pz�"��?s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA�|a]��A�4k �I K�$��BN,ZK�pz�#��@s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��a]��A�4k �I K�$��BN,ZK�ly� $��As�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��a]��A�4k �I K�$��BN,ZK�ly��%M�Bs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��a]��A�4k �I K�$��BN,ZK�ly��&M�Cs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��a]��A�4k �I K�$��BN,ZK�hy��'M�Ds�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I K�$��BN,ZK�hy��(M�Es�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I K�$��BN,ZK�hy��)M�Es�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I K"$��BN,ZK�hx��*M�Fs�T0 k� �(w�,w%�0d  U8D"!  ��"   � <�aA��b]��A�4k �I L"$��BN,ZK�dx��+M�Gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L"$��BN,ZK�dx��,M�Hs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L"$��BN0ZK�dx��-=�Is�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L"$��BN0ZK�dx=�/=�Js�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L"$��BN0ZK�`x=�0=�Ks�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L"$��BN0ZK�`x=�1=|Ls�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L"$��BN0ZK�`w=�2=xNs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L"$��BN0ZK�`w=�3=tOs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L"$��BN0ZK�`w=�5=lPs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L"$��BN0ZK�\w=�6=hQs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L�$��BN0ZK�\w=�7=dRs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L�$��BN0ZK�\w=�9=`Ts�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��b]��A�4k �I L�$��BN0ZK�\w=�:-XUs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L�$��BN0ZK�XwM�<-TVs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L�$��BN0ZK�XwM�=-PXs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L�$��BN0Z@�XvM�?-LYs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L�$��BN0Z@�XvM�@-H[s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L�$��BN0Z@�XvM�A-D\s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L�$��BN0Z@�Tv	]�B-@]s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L�$��BN4Z@�Tu	]�D-@_s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L�$��BN4ZE-Tu	]�E-<`s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L!�$��BN4ZE-Tt	]�F-8bs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L!�$�#�BN4ZE-Tt	]�G-8cs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I L!�$�#�BN4ZE-Tt	m�H4es�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I M!�$�'�BN4ZE-Ts	m�I4es�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I M!�$�'�BN4ZE-Xs	m�J0fs�T0 k� �(w�,w%�0d  U8D"!  ��"   � <�aA��c]��A�4k �I M!�$�+�BN4ZE-Xs	m�J0gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I M!�$�+�BN4ZE�Xs	m�K,hs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I  M!�$�/�BN4ZE�\s	]�L�(hs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I  M!�$3�M~4ZE�\r	]�M�$is�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I  M!�$3�M~4ZE�`r	]�M� j!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I  M!�$7�M~4ZE�`r	]�N� k!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I  M�$;�M~4ZE�dr	]�N�l!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��c]��A�4k �I  M�$?�M~4ZE�dq	m�O�l!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$?�M~4ZE�dq	m�O�m!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$C�M~4ZE�hp	m�O�n!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$G�M~4ZE�hp	m�P�o!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$K�M~4ZCMlo	m�P�o!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$O�M~4ZCMln	]�P�p!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$S�M�4ZCMln	]�Q�q!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$W�M�4ZCMpm	]�Q�r!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$[�M�8ZCMpm	]�Q� rs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$_�M�8ZCMpl	]�Q� ss�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$c�M�8ZCMpl	m�Q��ts�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$g�M�8ZCMpl	m�Q��ts�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I  M�$k�M�8ZCMpk	m�Q��us�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$o�M�8ZCMtk	m�Q��us�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$s�M�8ZCMtk	m�Q��vs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$w�M~8ZCMtk ��Q��ws�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�${�M~8ZC]tk ��Q��ws�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$�M~8ZC]tk ��Q��xs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$,��M~8ZC]tj ��Q��xs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$,��M~8ZC]tj ��Q��y!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$,��M~8ZC]tj m�Q��z!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$,��M~8ZC]tj m�Q��z!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$,��M~8ZC]ti m�Q��{!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$,��M~8ZC]ti m�Q��{!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �M�$,��BN8ZC]th m�Q��|!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �N�$,��BN8ZC]th m�Q��|!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �N�$,��BN8ZC]tg m�Q��}!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �N�$,� BN8ZCmtg m�Q��}!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �N�$,�BN8ZCmtf m�Q��~!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��d]��A�4k �I �N�$��BN8ZCmtf m�Q��~!��T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BN8ZCmte m�Q��s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BN8ZCmtd m�Q��s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BN8ZCmtd m�Q�̀s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BN8ZCmtc m�Q��s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��
BN8ZCmtc m�Q��s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BN8ZCmtc m�Q��s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BN8ZCmtb m�Q��s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BN8ZCmtb m�Q��s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BN8ZC}tb��Q��~s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BN<ZC}tb��Q��~s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$� BN<ZC}ta��Q��~s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$�BN<ZC}ta��Q��~s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$�BN<ZC}ta��Q��}s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$�BN<ZC}ta��Q��}s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$�BN<ZC}ta��Q��}s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$�BN<ZC}ta��Q��}s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$� BN<Z@�ta��Q��}s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$�(BN<Z@�ta��Q��|s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$�,BN<Z@�ta��Q��|s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$�0!BN<Z@�ta��Q��|s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$�8#BN<Z@�ta��Q��|s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$M<$BN<Z@�ta��Q��|s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$M@&BN<Z@�taͬQ��{s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$MH(BN<Z@�taͬQ�{s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$ML*BN<Z@mtaͬQ�{s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$MP+BN<Z@mtaͬQ�{s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$MT-BN<Z@mtaͬQ�{s�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$MX/BN<Z@mtaͬQ�zs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$M`1BN<Z@mtaͬQL�zs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$Md3BN<Z@mtaͬQL�zs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$Mh5BN<Z@mtaͬQL�zs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$Ml6BN<Z@mtaͬQL�ys�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$Mp8BN<Z@mtaͬQL�ys�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$]t:BN<Z@mtaͬQL�xs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$]x<BN<Z@mtaͬQL�xs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$]|>BN<Z@mtaͬQܰxs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$]�@BN<Z@taͬQܰws�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$]�BBN<Z@taͬQܰws�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BBN<Z@taͬRܰvs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��e]��A�4k �I �N�$��BBN<Z@taͰSܴvs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �N�$��CBN<Z@taͰS��us�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �N�$��DBN<ZK�taʹT��us�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �N�$��FBN<ZK�ta͸U��ts�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �N�$��GBN<ZK�ta͸U��ts�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �N�$��HBN<ZK�taͼV��ss�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �N�$͌IBN<ZK�taͼW��ss�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �N�$͐JBN<ZK�taͼX��ss�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �N�$͐KBN<ZK�ta��X��rs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �N�$͐MBN<ZK�ta��Y��rs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �N�$͐NBN<ZK�ta��Z��qs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$	}�OBN<ZK�ta��Z��qs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$	}�PBN<ZK�ta��[��qs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$	}�QBN<ZK�ta��\��ps�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$	}�RBN<ZK�ta��\��ps�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$	}�RBN<ZK�pa��]��os�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��RBN@ZK�pb��]��os�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��SBN@ZK�pb��^��os�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��SBN@ZK�pb��_��ns�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��TBN@ZK�pc��_��ns�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��TBN@ZK�pc��`��ns�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��UBN@ZK�lc��`��ms�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��UBN@ZK�ld��a� ms�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��VBN@ZK�ld��a�ms�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��VBN@ZK�ld��b�ls�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��WBN@ZK�le��b�ls�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��WBN@ZK�le��c�ks�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��XBN@ZK�le��c�ks�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�XBN@ZK�he��d� js�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�YBN@ZK�hf��d�(js�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�YBN@ZK�hf��e�(js�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�YBN@ZK�lf��e�,js�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�ZBN@ZK�lf��f�,is�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�ZBN@ZK�pf��f�0is�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�ZBN@ZK�pg��f�0is�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�ZBN@ZK�tg��f�4hs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�ZBN@ZK�tg��g�4hs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�ZBN@ZK�xg��g�8hs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�ZBN@ZK�xh��g�8gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�ZBN@ZK�|h��g�8gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�[BN@ZK�|h��g�<gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�[BN@ZK�|h��g�<gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�[BN@ZK��i ��g�<gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�[BN@ZK��i ��g�<gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�[BN@ZK��i ��g�<gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�[BN@ZK��i ��g�<gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZK��j ��g�@gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZK��j�g�@gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZK��j�g�@gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZK��j�g�@gs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZK��k�g�@fs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZK��k�g�Dfs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��k]�g�Dfs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��k]�g�Dfs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��k]�g�Hes�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��l]�g�Hes�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��l]�g�Les�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��l=�g�Lds�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��l=�g�Lds�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��l=�g�Pcs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��l=�g�Pcs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��l=�g�Pcs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��m=�g�Tcs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��m=�g�Tcs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��m=�g�Tcs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]BN@ZK��m=�g�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]M~@ZK��m=�gTbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]M~@Z@�m=�gTbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]M~@Z@�m=�gTbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��]M~@Z@�m=�gTbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��]M~@Z@�mM�gTbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��]M~@Z@�mM�g Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��]M~@Z@�mM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��]M~@Z@�mM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��]M~@Z@m�mM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��]M~@Z@m�mM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$��]M�@Z@m�mM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]M�@Z@m�mM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]M�@Z@m�mM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]M�@Z@��mM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]M�@Z@��lM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]M�@Z@��lM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�]M�@Z@��lM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��]M�@Z@��lM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��]M�@ZCM�lM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��]M~@ZCM�lM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��]M~@ZCM�lM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��]M~@ZCM�lM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��]M~@ZCM�lM�h Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��]M~@ZCM�lM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��]M~@ZCM�lM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��\M~@ZCM�lM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��\M~@ZC]�kM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��\M~@ZC]�kM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��\BN@ZC]�kM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��\BN@ZC]�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��\BN@ZC]�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$ ��\BN@ZC]�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZC]�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZC]�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZC]�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZC]�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZC]�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@Z@��jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@Z@��jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@Z@��jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@Z@��jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@Z@��jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZCM�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZCM�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$�\BN@ZCM�jM�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$�\BN@ZCM�j=�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$�\BN@ZCM�j=�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$]�\BN@ZCM�j=�i�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$]�\BN@ZCM�j=�i�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$]�\BN@ZCM�j=�i�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$]�\BN@ZCM�j=�i�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$]�\BN@ZKݔj=�i�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$]�\BN@ZKݔj=�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$]�\BN@ZKݔj=�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$]�\BN@ZKݔj=�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$]�\BN@ZKݐj=�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@ZKݐj=�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@ZKݐj=�h�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@ZKݐj=�g�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@ZKݐj=�g�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@ZKݐj=�g�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@ZKݐj=�f�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\BN@ZK݌j=�f�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�\M~@ZK݌jM�f�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�[M~@ZK݌jM�e�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�[M~@ZK�jM�e�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O�$]�[M~@ZK�jM�e�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aA��f]��A�4k �I �O!�$]�[M~@ZK�jM�e�Tbs�T0 k� �(w�,w%�0d  U8D"!  ��"    � <�aEXj���B�(.��WM(H�$���F�YQ;�D��*�P_s�T0 k� L�P��P%�0d  U8D"!  ��O    � 8�8E`i���B�4.��VM(J�$���F�]Q;�C��+�P]s�T0 k� ��Q��Q%�0d  U8D"!  .�O    � 8�8E`h���B�8.��VM(K�$���F�_Q;�B��,�P]s�T0 k� ��R��R%�0d  U8D"!  ��O    � 8�8Edg���B�<.��UM(L�$���E��aQ;�A��,�P\s�T0 k� ��S��S%�0d  U8D"!  ��O    � 8�8Ehf���B�D.��T=,M�$���E��cQ;�A��,�P[s�T0 k� ��T��T%�0d  U8D"!  ��O    � 8�8E�lf�×B�D/��T=,N�$���E��dQ;�@�-�PZs�T0 k� ��U��U%�0d  U8D"!  ��O    � 8�8E�td�˕B�D/�R=,P�$��E��hQ;�?�-�PXs�T0 k� ,�W��W%�0d  U8D"!  ��O    � 8�8E�xc�ӕB�D/�R=,Q�$��E��jQ;�?�-�PWs�T0 k� ,�W��W%�0d  U8D"! ��O    � 8�8E�|c�הB�H/�Q-,R�$��E��lQ;�>�-�PVs�T0 k� ,�X��X%�0d  U8D"! ��O    � 8�8E�b�ߔB�H/�Q-0S�$��E��mQ;�=�-�PUs�T0 k� ,�Y��Y%�0d  U8D"! ��O    � 8�8E�a��B�L/�P-0T�$��E��oQ;�=�-�PTs�T0 k� ,�Z��Z%�0d  U8D"! ��O    � 8�8E�a��B�P0� P-0U�$��E��qQ;�<��-�PSs�T0 k� ��[��[%�0d  U8D"! ��O    � 8�8                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \���Z ]�(^(^ h �� f��         ���
�     f����
�           	        	 
  ���          9�  �  ���   0
% 	          ��C�          ��y�+    ��C��y�+           	           @��          �  �  ���   0
 
          k�t          ��ܡ     k�t��ܡ                      ���          /�     ���  8

           IO�            �+��     IO��+��                      
	 A�$           0     ���   8          O;�            .�}��     O;��}��                         �$           ��      ���   P
	
          ��        B�	9�     ���	9�                             ���_             	  ���   P              []c    	   V�m%     [�$�mC�    ���            	 Z�a                 ��@   (
          Z�� � �
	     j���P     Z�����P                    N  Z�a         B`�     ��h   8�           j�� � �	   ~�ca�     j��cm�    ���L            t Z�a         ���  %  ��`  	@
           e.�  D D 
    ��z�F     eV��z�|    ���[             B Z�a         	 ڰb     ��@  H
$
          bږ  � �
     ��U�y     b���U�W    ���             \	 Z�a         
  �@�  	  ��`   H!	          �� ��	     � ��     �� ��                          	  ���$         �   C  ��@      0                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          w?�  ��        �����     w?�����                           x                j  �       �                          w    ��        ���       w  ��           "                                                �                         ���y���+�}�	�m���c�z�U �������                	 

   �    � �� ;�H       �� @h@ � @h� ��  i@ �D  p� ��  p� �� n� �D q` (� `r@ )D  s  �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0� ���� � � }`���� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����a�� <�� �  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    "�j�� , " �
� �  �  
�  k    ��     ���       k    ��     ���       Z    ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �"�      �� � �  ���        �t �  ���        �        ��        �        ��        �    ��    T�����        ��                         �$ (  ���                                     �                 ����             k�����%��   <�a��           �    18/41 (43%) e uk th    5:26                                                                        3  3     �C� �C� �=CB �-CF �2CJ �C �c� �c� �	c�- �
k~- �k�% � k�, �k�% �k�" �cV � c^ �B� � � B� � �c� � c�+ �C. � �8 � �7 �K( � K8 �kj � kr! � ks � kt PJ� h J�/ � "�# � !"�5 �"� �#
�. �$"�# � %"�5 �&"� �'*�. �("� � )"�$ �*� �+
� � ,*>| � -*l) .*LdA /*RdI  *lI  *lA 2*RdI  *l94*<dA5*2tY6*
lY *6tY *
lA9*2tY *6tY *6tY *
lY *
lY>*
lY *6t@�! 
�0 
�0                                                                                                                                                                                                 �� R @       �    @ 
        �     \ P E ^  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��    �H~�L� ��������������������������������������������������������   �4, 2   X� �����m� ���	����                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                         
      3    (    ��  D�J    	  4                             ������������������������������������������������������                                                                         
                                                              	      �      �      N                �  �          	  
 	 
 	 	 ��������������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� �                            
      F    )    ��	  H�J      �  	                           ������������������������������������������������������                                                                      
                                                                     �       �      �        �    ��              
 	  
	 
 	 	 ����� ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� �������������            �                                                                                                                                                                                                                                       
                                                                     �             


           �   }�         wwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwww N @ 0 
              	                  � W��( �h@                                                                                                                                                                                                                                                                                   )n)n1n  
1F                            d      m            `                                                                                                                                                                                                                                                                                                                                                                                                                     � � �  � ��  � ��  � @��  � #��  � ��  �����n����������n�����������9�����'����������y�                 u�> :�~ y        	 	 �   & AG� �  �   
              �                                                                                                                                                                                                                                                                                                                                      p B C   �     p                !��                                                                                                                                                                                                                            Y��   �� �� ��      �� B 	     ��������������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ������ ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� �������������             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    4      9      w                       B     �   ���������J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��    �   p���� ��     ! f  �  !l >     �f ��     �f �$ ^$ �@      ����� ��   �����    ����X ��   ����X �$ ^$     �  ��              +   ���X���� 
���������������h# Hj �  ��  �         ��   ���P h@ �� �� h@ �� �$ ^$         ��  <             ������          D��  �*  ��  yf  y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                                                �����   �   �   �   ����                                     
�  

  
 � 
 
 
   
   
   
   
  ��                  ��   
   
   
   
   
   
 
 
 � 

  
�                 �   
    �   
    �   
    �   
   
   �  
   �  
   �  
   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "  ""   "! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  ""   "! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "! ""! " "" """ "!   " ""            """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��� ���� ��    �     �                                                                                                                                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��     �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �    �  �  ��  �   �   �         �       �                        �   ��  ���  � �    �                                                                                                                                      �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        T   S   C   3   30  30  ;�  ��  ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                �   �               �  ��� ݼ� w{� �װ vw�           �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                          �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   2 1220!2 #!0 #      �  �   �   ��  �            ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �              �  �� ��  �    � ���                                                                                                                                                                                              �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �               �   �       �       Ț  ��  ��" �"��"/��"���  �     �   �   �   �      �  �                         �  ���          ���� ��� ����                �  ��  �                                      "  "  "      � �������������  �                                                                                                                                        UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �           J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"�  �             �   � �� ����ɪ�ܙ��� ��� ��� ��� ��� ��� ��� H��    �   ��  ��  ��  ט  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��                           � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �   �" �!  �  �� �   �                �  �� Ș ��  ��  �      �     �                                      � ����ݼ� ����                                                                                 �  �  ��  �                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                      �   �   �                           � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���      � �������������  �                                                                                                                                         �          �   �      "  �+ ɻ������̚� ��                        � U  X  �   �   �   �   � "� +���""�" �   ��  ��� ��� }�� w�z�w������������̽��̽��̽ۼ̽���л����������3X�DCX�T3�TC0�D30�M���K��� �������*�����"/��/���/  �              �  �  �  �  �  �   �     /�      �                           �   �   �   �   �   �   "  "  ""  "+� �� � ��   �  "   "�  +�  
�� ��� D�D 4ETO3    �   �   �   D   E�  U�  UO                         "  "  "                            ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                                  � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �        �  �  �   �   ��  �                            �   ���                            �   �                                                                                                   ̰ ˻ ���wݛk}�gz� w��  ��  ��  ��  ��  ,�  "�  �  ,�  "�  ..  ..  �  �   �                        �   �   ̰  ��  ��  ��� ��� �ܘ �ل@�؊@�4�@�H�@�D �@ �H� "H�""C�"ˋ" �" ��" "��� �  �                     ��  �                            �         �           �       �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                             �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                  ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                      ��  ��  ���                   ���                                      ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                     �  ��  ̽  ��  �w �
������������̽�̍������� ���  4� 4E    �   �   �   ڨ  ��� ��� ��ɨ�ͪ������˽��˽ۻ���������UUJ �  ��� ��  ��  ��  �  ��      �4DE�33E��;D����� �������� +�� �)�� ���                T�  UJ� UT� ET� D[� �� ��� ͻ�𽹀 �����ͻ� ��������/  �  �            /   �                    � ��� ��� ��  �                �   �     �   �           �  ��  ��  ��  ��� ��� ��� ��˰ɜ˰��˻�̻���������3���DDD�                                                                                                                                                                                                             �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(����������������� � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(����������������� 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5���������������� x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x���������������� w w x y�������H���������������������������������H������yxww����������������  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(���������������� , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,���������������� +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC� �C� �=CB �-CF �2CJ �C �c� �c� �	c�- �
k~- �k�% � k�, �k�% �k�" �cV � c^ �B� � � B� � �c� � c�+ �C. � �8 � �7 �K( � K8 �kj � kr! � ks � kt PJ� h J�/ � "�# � !"�5 �"� �#
�. �$"�# � %"�5 �&"� �'*�. �("� � )"�$ �*� �+
� � ,*>| � -*l) .*LdA /*RdI  *lI  *lA 2*RdI  *l94*<dA5*2tY6*
lY *6tY *
lA9*2tY *6tY *6tY *
lY *
lY>*
lY *6t3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������� ��5�K�\�O�T��=�U�J�J� � � � � � � � � � �/�.�7�������������������������������������������3�M�U�X��5�X�G�\�I�N�[�Q� � � � � � � �/�.�7����������������������������������������� ��=�K�X�X�_��B�G�Q�K� � � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������/�.�7� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�A�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                