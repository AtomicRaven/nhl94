GST@�                                                            \     �                                               � ���      �  �           ����e $�	 J�����������x�������        �g      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"��   " `  J  jF��    "�j "����
��
��     �j�� 
   ��
  �                                                                               ����������������������������������      ��    bb? QQ0 5 118 44                		 


     
               ��� 4    �                 nnY ))         88:�����������������������������������������������������������������������������������������������������������������������������==  00  44  11                                             ��  ��  ��  ��                  EE             �����������������������������������������������������������������������������                                D   P           @  &   z   �                                                                                 '      )n)nY  EE    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE P �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    XsA^O�A���]�+A��Y�7� �#�͔yC���G�!43��T0 k� �@��D�&�1D"3Q	24#Q  /�     ����ETsA^K�A���]�+A��Y�7� �#�͐yC���?�!03��T0 k� �<��@�&�1D"3Q	24#Q  ��     ����EPrA^K�A���]�+A��Y�7� �#�͌yI���7�!(3��T0 k� �8��<�&�1D"3Q	24#Q  ��     ����EPrA^G�A���]�+A��Y�7� �#�͌yI��/�!$3��T0 k� �8�<&�1D"3Q	24#Q  ��     ����ELrA^G�A���]�+A��Y�7� �#�͈yI�{�'�! 3��T0 k� �4�8&�1D"3Q	24#Q  ��     ����EHrA^C�A���]�+A��Y�7� �#�̈́yI�s��!3��T0 k� �0�4&�1D"3Q	24#Q  ��     ����EDqA^?�A���]�+A��Y�7� �#�̀yI�o��!3��T0 k� �,~�0~&�1D"3Q	24#Q  ��     ����E@qA^?�A���]�+A��Y�;� �#��|yI�g��!3��T0 k� �(~�,~&�1D"3Q	24#Q  ��     ����E<qA^;�A���]�+A��Y�;� �#��xyI�c��!3��T0 k� �$~�(~&�1D"3Q	24#Q  ��     ����E8pA^;�A���]�+A��Y�;��#��txI�_��!3��T0 k� � ~�$~&�1D"3Q	24#Q  ��     ����E4pA^7�A���]�+A��Y�;��#��pxI�[���!3��T0 k� �}� }&�1D"3Q	24#Q  ��     ����E0pA^7�A���]�+A��Y�;��#��lxI�[��� �3��T0 k� �}�}&�1D"3Q	24#Q  ��     ����E0pA^3�A���]�+A��Y�;��#��hxI�[��� �3��T0 k� �}�}&�1D"3Q	24#Q  ��     ����E,oA^3�A���]�+A��Y�;����dxI�[��� �3��T0 k� �|�|&�1D"3Q	24#Q  ��     ����E(oA^/�A���]�+A��Y�;����`xI�W��� �3��T0 k� �|�|&�1D"3Q	24#Q  ��     ����E$oA^/�A���]�+A��Y�;����`xI�W��� �3��T0 k� �|�|&�1D"3Q	24#Q  ��     ����E nA^+�A���]�+A��Y�?����\wI�S��� �3��T0 k� �|�|&�1D"3Q	24#Q  ��     ����E nA^+�A���]�+A��Y�?����XwLS� �� �3��T0 k� �{�{&�1D"3Q	24#Q  ��     ����EnA^'�A���]�+A��Y�?����TwLS� �� �3��T0 k� �{�{&�1D"3Q	24#Q  ��     ����EnA^'�A���]�+A��Y�?���PwLS� �� �3��T0 k� � {�{&�1D"3Q	24#Q  ��     ����EmA^#�A���]�+A��Y�?���PwLO� �� �3��T0 k� ��{� {&�1D"3Q	24#Q  ��     ����EmA^#�A���]�+A��Y�?���LwLO� �� �3��T0 k� ��z��z&�1D"3Q	24#Q  ��     ����EmA^#�A���]�+A��Y�?���HwLO� �� �3��T0 k� ��z��z&�1D"3Q	24#Q  ��     ����EmA^�A���]�+A��Y�?���DvLK� �� �3��T0 k� ��z��z&�1D"3Q	24#Q  ��     ����EmA^�A���]�+A��Y�?���DvLK� �� �3��T0 k� ��z��z&�1D"3Q	24#Q  ��     ����ElA^�A���]�+A��Y�?���@vLK� �� �3��T0 k� ��y��y&�1D"3Q	24#Q  ��     ����ElA^�A���]�+A��Y�?���<vLG� �� �3��T0 k� ��y��y&�1D"3Q	24#Q  ��     ����ElA^�A���]�+A��Y�C���8vLG� ���3��T0 k� ��y��y&�1D"3Q	24#Q  ��     ����E lA^�A���]�+A��Y�C���8vLG� ���3��T0 k� ��y��y&�1D"3Q	24#Q  ��     ����E�kA^�A���]�+A��Y�C���4vLG� ���3��T0 k� ��y��y&�1D"3Q	24#Q  ��     ����E�kA^�A���]�+A��Y�C���0vL-C� ���3��T0 k� ��x��x&�1D"3Q	24#Q  ��     ����E�kA^�A���]�+A��Y�C���0vL-C� ��3��T0 k� ��x��x&�1D"3Q	24#Q  ��     ����E�kA^�A���]�+A��Y�C���,uL-C� {��3��T0 k� ��x��x&�1D"3Q	24#Q  ��     ����E�kA^�A���]�+A��Y�C���,uL-C� w��3��T0 k� ��x��x&�1D"3Q	24#Q  ��     ����E�jA^�A���]�+A��Y�C���(uL-?� s��3��T0 k� ��x��x&�1D"3Q	24#Q  ��     ����E�jA^�A���]�+A��Y�C���$uL-?� k��3��T0 k� ��w��w&�1D"3Q	24#Q  ��     ����E�jA^�A���]�+A��Y�C���$uL-?� g��3��T0 k� ��w��w&�1D"3Q	24#Q  ��     ����E�jA^�A���]�+A�Y�C��� uL-?� c���3��T0 k� ��w��w&�1D"3Q	24#Q  ��     ����E�jA^�A���]�+A�Y�C��� uL-;� _��3��T0 k� ��w��w&�1D"3Q	24#Q  ��     ����E�jA^�A���]�+A�Y�C���uL-;� [��3��T0 k� ��w��w&�1D"3Q	24#Q  ��     ����E�iA^�A���]�+A�Y�C����uL-;� W��3��T0 k� ��v��v&�1D"3Q	24#Q  ��     ����E�iA^�A���]�+A�Y�G����uL-;� S��3��T0 k� ��v��v&�1D"3Q	24#Q  ��     ����E�iA^�A���]�+A�Y�G����tL-7� O��3��T0 k� ��v��v&�1D"3Q	24#Q  ��     ����E�iA^�A���]�+A�Y�G����tL-7� K��3��T0 k� ��v��v&�1D"3Q	24#Q  ��     ����E�iA^�A���]�+A�Y�G����tL-7� G��3��T0 k� ��v��v&�1D"3Q	24#Q  ��     ����E�iA]��A���]�+A�Y�G����tL-7� C�|3��T0 k� ��v��v&�1D"3Q	24#Q  ��     ����E�hA]��A���]�+A�Y�G����tL-7� ?�|3��T0 k� ��u��u&�1D"3Q	24#Q  ��     ����E�hA]��A���]�+A�Y�G����tL-3� ;�x3��T0 k� ��u��u&�1D"3Q	24#Q  ��     ����E�hA]��A���]�+A�Y�G����tL-3� 7�t3��T0 k� ��u��u&�1D"3Q	24#Q  ��     ����E�hA]��A���]�+A�Y�G����tL-3� 3�p3��T0 k� ��u��u&�1D"3Q	24#Q  ��     ����E�hA]��A���]�+A�Y�G����tL-3� /�l3��T0 k� ��u��u&�1D"3Q	24#Q  ��     ����E�hA]��A���]�+A�Y�G����tL-3� +� l3��T0 k� ��u��u&�1D"3Q	24#Q  ��     ����E�hA]��A���]�+A�Y�G���� tL-/� '� h3��T0 k� ��u��u&�1D"3Q	24#Q  ��     ����E�gA]��A���]�+A�Y�G���� sL-/� #� d3��T0 k� ��t��t&�1D"3Q	24#Q  ��     ����E�gA]��A���]�+A�Y�G����sL-/� � `3��T0 k� ��t��t&�1D"3Q	24#Q  ��     ����E�gA]��A���]�+A�Y�G����sL-/� � `3��T0 k� ��t��t&�1D"3Q	24#Q  ��     ����E�gA]�A���]�+A�Y�G����sL-/� � \3��T0 k� ��t��t&�1D"3Q	24#Q  ��     ����E�gA]�A���]�+A�Y�K����sL-+� � X3��T0 k� ��t��t&�1D"3Q	24#Q  ��     ����E�gA]�A���]�+A�Y�K����sL-+�� T3��T0 k� ��t��t&�1D"3Q	24#Q  ��     ����E�gA]�A���]�+A�Y�K����sL-+�� T3��T0 k� ��t��t&�1D"3Q	24#Q  ��     ����E�fA]�A���]�+A�Y�K����sL-+�� P3��T0 k� ��s��s&�1D"3Q	24#Q  ��     ����E�fA]�A���]�+A�Y�K����sL-+�� L3��T0 k� ��s��s&�1D"3Q	24#Q  ��     ����E�fA]�A���]�+A�Y�K����sL-+�� L3��T0 k� ��s��s&�1D"3Q	24#Q  ��     ����E�fA]�A���]�+A�Y�K����sL-'�� H3��T0 k� ��s��s&�1D"3Q	24#Q  ��     ����E�fA]�A���]�+A�Y�K����sL-'���� H3��T0 k� ��s��s&�1D"3Q	24#Q  ��     ����E�fA]�A���]�+A�Y�K����sL-'���� D3��T0 k� ��s��s&�1D"3Q	24#Q  ��     ����E�fA]�A���]�+A�Y�K����sL-'���� @3��T0 k� ��s��s&�1D"3Q	24#Q  ��     ����E�fA]�A���]�+A�Y�K����sL-'���� @3��T0 k� ��s��s&�1D"3Q	24#Q  ��     ����E�fA]�A���]�+A�Y�K����rL-'���� <3��T0 k� ��s��s&�1D"3Q	24#Q  ��     ����E�eA]�A���]�+A�Y�K����rL-'���� <3��T0 k� ��r��r&�1D"3Q	24#Q  ��     ����E�eA]�A���]�+A�Y�K����rL-#���� 83��T0 k� ��r��r&�1D"3Q	24#Q  ��     ����E�eA]�A���]�+A�Y�K����rL#���� 43��T0 k� ��r��r&�1D"3Q	24#Q  ��     ����E�eA]�A���]�+A�Y�K����rL#���� 03��T0 k� ��r��r&�1D"3Q	24#Q  ��     ����E�eA]�A���]�+A�Y�K����rL#���� 03��T0 k� ��r��r&�1D"3Q	24#Q  ��     ����E�eA]�A���]�+A�Y�K� ���rL#���� ,3��T0 k� ��r��r&�1D"3Q	24#Q  ��     ����E�eA]�A���]�+A�Y�K� ���rL#���� ,3��T0 k� ��r��r&�1D"3Q	24#Q  ��     ����E�eA]�A���]�+A�Y�O� ���rL#���� (3��T0 k� ��r��r&�1D"3Q	24#Q  ��     ����E�eA]�A���]�+A�Y�O� ���rL#���� (3��T0 k� ��r��r&�1D"3Q	24#Q  ��     ����E�dA]�A���]�+A�Y�O� ���rL#���� $3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�dA]ߋA���]�+A�Y�O� ���rL#���� $3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�dA]ߋA���]�+A�Y�O� ���rA]#����  3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�dA]ߋA���]�+A�Y�O� l��rA]#����  3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�dA]ߋA���]�+A�Y�O� l��rA]#���� 3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�dA]ߋA���]�+A�Y�O� l��rA]#��� 3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�dA]ߋA���]�+A�Y�O� l��rA]#��� 3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�dA]ߋA���]�+A�Y�O� l��rA�#��� 3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�dA]ۋA���]�+A�Y�O����rA�#��� 3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�dA]ۋA���]�+A�Y�O����rA�#��� 3��T0 k� ��q��q&�1D"3Q	24#Q  ��    ����E�dA]ۋA���]�+A�Y�O����qA�#��� 3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�dA]ۊA���]�+A�Y�O����qA�#��{� 3��T0 k� ��q��q&�1D"3Q	24#Q  ��     ����E�cA]ۊA���]�+A�Y�O����qA�#��s� 3��T0 k� ��p��p&�1D"3Q	24#Q  ��     ����E�cA]ۊA���]�+A�Y�O����qA�#��k�3��T0 k� ��p��p&�1D"3Q	24#Q  ��     ����E�cA]ۊA���]�+A�Y�O����qA�#��g�3��T0 k� ��p��p&�1D"3Q	24#Q  ��     ����E�cA]׊A���]�+A�Y�O����qA�#�?_�3��T0 k� �|p��p&�1D"3Q	24#Q  ��     ����E�cA]׊A���]�+A�Y�O����qA�#�?W�3��T0 k� �|p��p&�1D"3Q	24#Q  ��     ����E�cA]׊A���]�+A�Y�O����qA�#�?S�3��T0 k� �|p��p&�1D"3Q	24#Q  ��     ����E�cA]׊A���]�+A�Y�O�����qA�#�?K�3��T0 k� �|p��p&�1D"3Q	24#Q  ��     ����E�cA]׊A���]�+A�Y�O�����qA�#�?C��3��T0 k� �xp�|p&�1D"3Q	24#Q  ��     ����E�cA]׊A���]�+A�Y�O�L���qA�#�??�� 3��T0 k� �xp�|p&�1D"3Q	24#Q  ��     ����E�cA]׊A���]�+A�Y�O�L���qA�#�?7�� 3��T0 k� �xp�|p&�1D"3Q	24#Q  ��     ����E�cA]ӊA���]�+A�Y�O�L���qA�#�?/���3��T0 k� �xp�|p&�1D"3Q	24#Q  ��     ����E�cA]ӊA���]�+A�Y�O�L���qA�'�?'���3��T0 k� �xp�|p&�1D"3Q	24#Q  ��    ����E�cA]ӊA���]�+A�Y�O�L���qA�'�?#���3��T0 k� �tp�xp&�1D"3Q	24#Q  ��     ����E�cA]ӊA���]�+A�Y�S�����qA�'�?���3��T0 k� �tp�xp&�1D"3Q	24#Q  ��    ����E�cA]ӊA���]�+A�Y�S����qA�'�?���3��T0 k� �tp�xp&�1D"3Q	24#Q  ��     ����E�bA]ӊA���]�+A�Y�S����qA�'�O���3��T0 k� �to�xo&�1D"3Q	24#Q  ��     ����E�bA]ӊA���]�+A�Y�S����qA�'�O���3��T0 k� �to�xo&�1D"3Q	24#Q  ��     ����E�bA]ӉA���]�+A�Y�S����qA�'�N����3��T0 k� �to�xo&�1D"3Q	24#Q  ��     ����E�bA]ӉA���]�+A�Y�S����qA�'�N����3��T0 k� �po�to&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�N����3��T0 k� �po�to&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�N����3��T0 k� �po�to&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�N����3��T0 k� �po�to&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�N����3��T0 k� �po�to&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�N����3��T0 k� �lo�po&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�N����3��T0 k� �lo�po&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�N����3��T0 k� �lo�po&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�^����3��T0 k� �lo�po&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�^����3��T0 k� �lo�po&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�^��?�3��T0 k� �lo�po&�1D"3Q	24#Q  ��     ����E�bA]ωA���]�+A�Y�S����qA�'�^��?�3��T0 k� �lo�po&�1D"3Q	24#Q  ��     ����E�bA]ˉA���]�+A�Y�S����pA�'�^��?�3��T0 k� �ho�lo&�1D"3Q	24#Q  ��     ����E�bA]ˉA���]�+A�Y�S����pA�'�^��?�3��T0 k� �ho�lo&�1D"3Q	24#Q  ��     ����E�bA]ˉA���]�+A�Y�S����pA�'�^��?�
3��T0 k� �ho�lo&�1D"3Q	24#Q  ��     ����E�bA]ˉA���]�+A�Y�S����pA�'�^��?�	3��T0 k� �ho�lo&�1D"3Q	24#Q  ��     ����E�bA]ˉA���]�+A�Y�S����pA�'�^��?�	3��T0 k� �ho�lo&�1D"3Q	24#Q  ��     ����E�bA]ˉA���]�+A�Y�S����pA�'�^�?�3��T0 k� �hn�ln&�1D"3Q	24#Q  ��     ����E�aA]ˉA���]�+A�Y�S����pA�'�^w�?�3��T0 k� �hn�ln&�1D"3Q	24#Q  ��     ����E�aA]ˉA���]�+A�Y�S����pA�'�ns�?�3��T0 k� �dn�hn&�1D"3Q	24#Q  ��    ����E�aA]ˉA���]�+A�Y�S����pA�'�nk�?�3��T0 k� �dn�hn&�1D"3Q	24#Q  ��     ����E�aA]ˉA���]�+A�Y�S����pA�'�nc�?�3��T0 k� �dn�hn&�1D"3Q	24#Q  ��     ����E�aA]ˉA���]�+A�Y�S����pA�'�n[�O�3��T0 k� �dn�hn&�1D"3Q	24#Q  ��     ����E�aA]ˉA���]�+A�Y�S����pA�'�nW�O|3��T0 k� �dn�hn&�1D"3Q	24#Q  ��     ����E�aA]ˉA���]�+A�Y�S����pA�'�^O�Ot3��T0 k� �dn�hn&�1D"3Q	24#Q  ��     ����E�aA]ǉA���]�+A�Y�S����pA�'�^G�Op3��T0 k� �dn�hn&�1D"3Q	24#Q  ��     ����E|aA]ǉA���]�+A�Y�S����pA�'�^C�Ol3��T0 k� �dn�hn&�1D"3Q	24#Q  ��     ����E|aA]ǈA���]�+A�Y�S����pA�'�^;�?h3��T0 k� �`n�dn&�1D"3Q	24#Q  ��     ����E|aA]ǈA���]�+A�Y�S����pA�'�^3�?` 3��T0 k� �`n�dn&�1D"3Q	24#Q  ��     ����E|aA]ǈA���]�+A�Y�S����pA�'�^+�?\ 3��T0 k� �`n�dn&�1D"3Q	24#Q  ��     ����E|aA]ǈA���]�+A�Y�S����pA�'�^'�?[�3��T0 k� �`n�dn&�1D"3Q	24#Q  ��     ����E|aA]ǈA���]�+A�Y�S����pA�'�^�?W�3��T0 k� �`n�dn&�1D"3Q	24#Q  ��     ����E|aA]ǈA���]�+A�Y�W����pA�'�^�?O�3��T0 k� �`n�dn&�1D"3Q	24#Q  ��     ����E|aA]ǈA���]�+A�Y�W����pA�'���?K�3��T0 k� �`n�dn&�1D"3Q	24#Q  ��     ����E|aA]ǈA���]�+A�Y�W����pA�'���?G�3��T0 k� �`n�dn&�1D"3Q	24#Q  ��     ����ExaA]ǈA���]�+A�Y�W����pA�'���?C�3��T0 k� �`n�dn&�1D"3Q	24#Q  ��     ����ExaA]ǈA���]�+A�Y�W����pA�'����??�3��T0 k� �`n�dn&�1D"3Q	24#Q  ��     ����ExaA]ǈA���]�+A�Y�W����pA�'����?;�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��     ����ExaA]ǈA���]�+A�Y�W��ߣ�pA�'����O7�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��     ����ExaA]ǈA���]�+A�Y�W��ߣ�pA�'����O3�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��    ����ExaA]ǈA���]�+A�Y�W��ߣ�pA�'����O/�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��     ����ExaA]ǈA���]�+A�Y�W��ߣ�pA�'����O+�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��     ����ExaA]ÈA���]�+A�Y�W��ߣ�pA�'��ϿO'�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��     ����ExaA]ÈA���]�+A�Y�W��ߤ�pA�'��˾O#�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��     ����ExaA]ÈA���]�+A�Y�W��ߤ�pA�'��ýO�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��     ����ExaA]ÈA���]�+A�Y�W��ߤ�pA�'�=��O�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��     ����EtaA]ÈA���]�+A�Y�W��ߤ�pA�'�=��O�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��     ����EtaA]ÈA���]�+A�Y�W��ߤ�pA�'�=��O�3��T0 k� �\n�`n&�1D"3Q	24#Q  ��     ����EtaA]ÈA���]�+A�Y�W��ߤ�pA�'�=��O�3��T0 k� �Xn�\n&�1D"3Q	24#Q  ��     ����EtaA]ÈA���]�+A�Y�W��ۥ�pA�'�=��O�"s��T0 k� �Xn�\n&�1D"3Q	24#Q  ��     ����EtaA]ÈA���]�+A�Y�W��ۥ�pA�'�	���O�"s��T0 k� �Xn�\n&�1D"3Q	24#Q  ��    ����EtaA]ÈA���]�+A�Y�W��ۥ�pA�'�	���O�"s��T0 k� �Xn�\n&�1D"3Q	24#Q  ��     ����EtaA]ÈA���]�+A�Y�W��ۥ�pA�'�	���N��"s��T0 k� �Xm�\m&�1D"3Q	24#Q  ��     ����EtaA]ÈA���]�+A�Y�W� lۥ�pA�'�	���N��"s��T0 k� �Xm�\m&�1D"3Q	24#Q  ��     ����Et`A]ÈA���]�+A�Y�W� lۦ�pA�'�	���N��"s��T0 k� �Xm�\m&�1D"3Q	24#Q  ��     ����Et`A]ÈA���]�+A�Y�W� lۦ�pA�'�	̓�N��"s��T0 k� �Xm�\m&�1D"3Q	24#Q  ��     ����Et`A]ÈA���]�+A�Y�W� lۦ�pA�'�	�{�N��"s��T0 k� �Xm�\m&�1D"3Q	24#Q  ��     ����Et`A]ÈA���]�+A�Y�W� lߧ�pA�'�	�w�N��"s��T0 k� �Xm�\m&�1D"3Q	24#Q  ��     ����Et`A]ÈA���]�+A�Y�W�ߧ�pA�'�	�s�N��"s��T0 k� �Xm�\m&�1D"3Q	24#Q  ��     ����Et`A]ÈA���]�+A�Y�W�ߧ�pA�'�	�o�N��"s��T0 k� �Xm�\m&�1D"3Q	24#Q  ��     ����Ep`A]ÈA���]�+A�Y�W�ߨ�pA�'�=k�N��3��T0 k� �Xm�\m&�1D"3Q	24#Q  ��     ����Ep`A]ÈA���]�+A�Y�W���pL]'�=g�N��3��T0 k� �Xm�\m&�1D"3Q	24#Q  ��     ����Ep`A]ÈA���]�+A�Y�W���pL]'�=c�N��3��T0 k� �Tm�Xm&�1D"3Q	24#Q  ��     ����Ep`A]ÈA���]�+A�Y�W���pL]'�=_�N��3��T0 k� �Tm�Xm&�1D"3Q	24#Q  ��    ����Ep`A]ÈA���]�+A�Y�W���pL]'�=[�N��3��T0 k� �Tm�Xm&�1D"3Q	24#Q  ��     ����Ep`A]ÈA���]�+A�Y�W���pL]'�=W�N��3��T0 k� �Tm�Xm&�1D"3Q	24#Q  ��     ����Ep`A]ÈA���]�+A�Y�W���pL]'�=W�N��3��T0 k� �Tm�Xm&�1D"3Q	24#Q  ��     ����E�,KB�'�S��� E�Y|#�!7��4D"?��g��3�"s��T0 k� "�&�1D"3Q	24#Q �?    ��� ��8LB�+�S���E�
Y|#�!;��2D"C��g��/�"s��T0 k� "�&�1D"3Q	24#Q ��?    ��� ��@LB�3�U����E�	Y|#�!C��0D"D �g��+�"s��T0 k� "�&�1D"3Q	24#Q ��?    ��� ��HLB�7�U����B��Y|#�!G��.D"H�g��'�"s��T0 k� "�&�1D"3Q	24#Q ��?    ��� ��PLB�;�U����	B��Y|#�K��,D"L�c��#�3��T0 k� ��&�1D"3Q	24#Q ��?    ��� �`MB�G�U����B��Y|#�W��(ObT
�c�C�3��T0 k� ��&�1D"3Q	24#Q ��?    ��� �hMB�K�U����B��Y|#�_��&ObT�_�C�3��T0 k� ��&�1D"3Q	24#Q ��?    ��� �pMB�S�U����B�� Y|#�c��$ObX�_�C�3��T0 k� ��&�1D"3Q	24#Q ��?    ��� �|MB�W�U����B���Y|#�g��"Ob\3_�C�3��T0 k� 2�&�1D"3Q	24#Q ��?    ��� ��MB�_�U����B���Y|#�o��� Ob`3[�C�3��T0 k� 2�&�1D"3Q	24#Q ��?    ��� ��NB�_�A�� B���Y|#�w���Obd3[�C�3��T0 k� 2�&�1D"3Q	24#Q ��?    ��� ��NB�_�A��$B���Y|#�{���Obh3W�B��3��T0 k� 2�&�1D"3Q	24#Q ��?    ��� ��NB�g�A��(B���Y|#�����Obp3W�B�3��T0 k� 2�&�1D"3Q	24#Q ��?    ��� ��NB�k�A��,B���Y|#�����Obp3S�2�"���T0 k� ��&�1D"3Q	24#Q ��?    ��� ���NB�o�Eq���,B���Y|#�����Obt3S�2�"���T0 k� ��&�1D"3Q	24#Q ��?    ��� ���NB�s�Eq���0B���Y|#������Obx!3O�2�"���T0 k� ��&�1D"3Q	24#Q ��?    ��� ���OB�{�Eq���4B���Y|#������Ob|#3O�2�"���T0 k� �� &�1D"3Q	24#Q ��?    ��� ���OB�{�Eq���8 B���Y|#����� Ob�'CK�2�
"���T0 k� �� &�1D"3Q	24#Q ��?    ��� ���OB��Ea���8"B���Y|#�����Ob�)CK�2�"���T0 k� "� &�1D"3Q	24#Q ��?    ��� ���NBу�Ea���<#B���Y|#�����Ob�+CG�2�"���T0 k� "� &�1D"3Q	24#Q $�?    ��� ���NBы�Ea���@$B���Y|#�����
Ob�-CG�2�"���T0 k� " �$&�1D"3Q	24#Q ��?    ��� ��NBы�Eaê�D'B���Y|#�����Ob�0�C�2�"���T0 k� " �$&�1D"3Q	24#Q ��?    ��� ��NBя�D1ë�D(B���Y|#����� Ob�2�?�2�3��T0 k� " �$&�1D"3Q	24#Q ��?    ��� ��NBї�D1ì�H)B���Y|#�����(Eb�4�?�"�3��T0 k� "$�(&�1D"3Q	24#Q ��?    ��� ��NBћ�D1í�H*B���Y|#�����,Eb�6�;�"�3��T0 k� "$�(&�1D"3Q	24#Q ��?    ��� �r,MB���D1ï�P-B���Y|#�q���8 Eb�9�7�"�3��T0 k� �(�,&�1D"3Q	24#Q ��?    ��� �r4MB���D1ð�P.B���Y|#�q���C�Eb�;�3�"�3��T0 k� �(�,&�1D"3Q	24#Q ��?    ��� �r<LB���D1ñ�T/B���Y|#�r��G�ER�=�/�"�3��T0 k� �(�,&�1D"3Q	24#Q ��?    ��� �rDLB���D1ó�T0B��Y|#�r��O�ER�?�+�"�!3��T0 k� �,�0&�1D"3Q	24#Q ��?    ��� �rTKB�˜DAõ�X2B��Y|#�r��[�ER�C�'�"�%3��T0 k� B,�0&�1D"3Q	24#Q ��?    ��� �r\JB�ӜDAö�\3B��Y|#����c�ER�E3#�"�'3��T0 k� B,�0&�1D"3Q	24#Q ��?    ��� �rdJB�ۛDA÷�\5B��Y|#����k�ER�F3�"�(3��T0 k� B8�<&�1D"3Q	24#Q ��7    ��� �rdJB��DA���`7B�+�Y|#��'��w�ER�J3�"�,3��T0 k� BL�P&�1D"3Q	24#Q ��7    ��� �rdJB��DA���d8B�/�Y|#��/��{�ER�K3�"�.3��T0 k� �X
�\
&�1D"3Q	24#Q ��7    ��� �rhIB���DA���d9B�7�Y|#��3����ER�M3��.3��T0 k� �`
�d
&�1D"3Q	24#Q ��'    ��� �rhIB��Ea���d9E?�Y|#��7����ER�N3��.3��T0 k� �l
�p
&�1D"3Q	24#Q ��'    ��� �rlIB��Ea���d9EK�Y|#��C����ER�QC��13��T0 k� �|	��	&�1D"3Q	24#Q  ��'    ��� �rpIB��Ea���d9ES�Y|#�rK����ER�SC��23��T0 k� "�	��	&�1D"3Q	24#Q  ��'    ��� �rpJB��Ea���`9E[�Y|#�rO����EB�TC���33��T0 k� "�	��	&�1D"3Q	24#Q  -�'    ��� �rtJI/�Ea���`:Eg�Y|#�r[����EB�WC���63��T0 k� "�	��	&�1D"3Q	24#Q  ��'    ��� �rxJI7�Ea���`:Eo�Y|#�r_����EB�X2����73��T0 k� "�	��	&�1D"3Q	24#Q  ��'    ��� �rxKI;�Ea���`;Ew�Y|#�rc�·�EB�Z2����83��T0 k� ����&�1D"3Q	24#Q  ��'   ��� �r|KIC�Ea���`;E�Y|#�rk�»�C��[2����93��T0 k� ����&�1D"3Q	24#Q ��'    ��� �r�KI"O�Ea���`;E��a�#�rs�»�C��]2� ��<3��T0 k� ����&�1D"3Q	24#Q ��'    ��� �r�KI"S�EQ���\<E���a�#�r{�»�C��^2���=3��T0 k� ����&�1D"3Q	24#Q ��'    ��� �r�LI"[�EQ���\<E���a�#�r{�¿�C��_2���>3��T0 k� 2���&�1D"3Q	24#Q ��'    ��� �r�LI"c�EQ���\=E���a�#�r����C��`"���A3��T0 k� 2���&�1D"3Q	24#Q ��'    ��� �r�LIk�EQ���\=E���a�#�b�����C��a"�
��B3��T0 k� 2���&�1D"3Q	24#Q ��'    ��� �r�LIo�EQ���\=E���a�#�b�����C��b"���C3��T0 k� 2���&�1D"3Q	24#Q ��'    ��� �r�MIs�EQ���\=E���a�#�b�����C��b"���D3��T0 k� ����&�1D"3Q	24#Q ��'    ��� �r�MI{�EQw��\>E���a�#�b�����C��c"���F3��T0 k� �� �� &�1D"3Q	24#Q ��'    ��� �r�MI"�EQs��X>E���Y|#�b�����C��d"���G3��T0 k� ������&�1D"3Q	24#Q ��'    ��� �r�MI"��EQo��X>E���Y|#�b�����C��d"��H3��T0 k� ������&�1D"3Q	24#Q ��'    ��� �r�NI"��EQc��X?E���Y|#�2�����C��e"��J3��T0 k� "�����&�1D"3Q	24#Q  ��'    ��� �b�NI"��EQ[��X?E���Y|#�2��b��C��e"��K3��T0 k� "�����&�1D"3Q	24#Q  ��'    ��� �b�NE���EQW��X?E��Y|#�2��b��C��e"�L3��T0 k� "�����&�1D"3Q	24#Q  ��'    ��� �b�NE���EAG��X@Ep�Y|#�2��b��C��e"�!N3��T0 k� "�����&�1D"3Q	24#Q  /�'    ��� �b�NE���EAC��X@Ep�Y|#�b��b��C��e�#O3��T0 k� �����&�1D"3Q	24#Q  ��'    ��� ���NE���EA;��X@Ep�Y|#�b��b��C��e�%P3��T0 k� �����&�1D"3Q	24#Q  ��'    ��� ���NE���EA/��TAEp+�Y|#�b��b� C�|e�),R3��T0 k� �x �| &�1D"3Q	24#Q  ��'    ��� ���ME���EA'��TAEp3�a�#�b��b� C�xe�+0S3��T0 k� �t�x&�1D"3Q	24#Q  ��'    ��� ���ME���EA��TAEp;�a�#�b��b�C�te�-8T3��T0 k� �t�x&�1D"3Q	24#Q  ��'    ��� �R�ME�ßEA��TBEpG�a�#�b��b�C�hd�0�HU3��T0 k� �l�p&�1D"3Q	24#Q  ��'    ��� �R�MErˠEA��TBEpO�a�#�b��r�C�dd�2�PV3��T0 k� �l�p&�1D"3Q	24#Q  ��'    ��� �R�MErϠEA��TBEpS�a�#�b��r�C�`d 4�TW3��T0 k� �l�p&�1D"3Q	24#Q  ��'    ��� �R�MErӡE@���TBE`[�a�#�R��r�C�\c6�\X3��T0 k� �l�p&�1D"3Q	24#Q  ��'    ��� ��MErߣE@���TCE`g�a�#�R��r�C�Pb9�lY3��T0 k� �h�l&�1D"3Q	24#Q  ��'    ��� ��MEr�C����TCE`k�a�#�R��r�C�Lb;�tY3��T0 k� �d�h&�1D"3Q	24#Q  ��'    ��� ��MEr�C����PCE`s�a�#�R��r�C�Da�<�|Z3��T0 k� �`�d&�1D"3Q	24#Q  ��'    ��� ��MEr�C����PCE`w�Y|#�R��ҤC�@a�>��Z3��T0 k� �d�h&�1D"3Q	24#Q  ��'    ��� ��NEr��C����LCE`�Y|#�R��ҜC�4_�A��[3��T0 k� �d�h&�1D"3Q	24#Q  ��    ��� ��NEr��Ip���LCE`��Y|#���ҘC�,^�B��[3��T0 k� �d�h&�1D"3Q	24#Q  ��    ��� ��NEr��Ip���LCE`��Y|#��{�ҔC�(^� Cs�\3��T0 k� �d�h&�1D"3Q	24#Q  ��    ��� ��|NEs�Ip���HCE`��Y|#��w�҈C�\�(Fs�\3��T0 k� �\�`&�1D"3Q	24#Q  ��    ��� ��xNEc�Ip���HCE`��Y|#��o�҄C�[�0Gs�\3��T0 k� �\�`&�1D"3Q	24#Q  ��    ��� ~�xNEc�I����DCE`��Y|#��k�Ҁ	C�Z�4Hs�\3��T0 k� �X�\&�1D"3Q	24#Q  ��    ��� {RtNEc�I����DCEP��Y|#��g��x	C�Y�8Is�\3��T0 k� �P�T&�1D"3Q	24#Q  ��    ��� xRtNEc�I����@CEP��Y|#��_��l
C��W�@Ks�\3��T0 k� �H�L&�1D"3Q	24#Q  ��    ��� tRpNEc�I����<CEP��Y|#��[��h
C��VsDLs�\3��T0 k� �G��K�&�1D"3Q	24#Q  ��    ��� qRpNEc�E���<CEP��Y|#��S��d
EA�UsHMs�\3��T0 k� �C��G�&�1D"3Q	24#Q  ��    ��� nRlNEc#�E�{��<BEP��Y|#��O��\
EA�TsLNs�[3��T0 k� �?��C�&�1D"3Q	24#Q  ��    ��� kRlNEc'�E�k��8BEP��Y|#��C��PEA�RsTOs�[3��T0 k� �3��7�&�1D"3Q	24#Q  ��    ��� hRlNEc'�E�g��4BC��Y|#��?��HEA�Ps\Ot Z3��T0 k� �+��/�&�1D"3Q	24#Q  ��    ��� eRhOEc+�E�_��4BC��Y|#��7��DEA�Os`PdZ3��T0 k� �'��+�&�1D"3Q	24#Q  ��    ��� b�dOEc+�E�W��0AC��Y|#��/��<EA�NsdPdY3��T0 k� ���#�&�1D"3Q	24#Q  ��   ��� _�\OEc/�E�K��,AC��Y|#��#��0
EA�KslQdX3��T0 k� ����&�1D"3Q	24#Q  ��    ��� \�XOEc/�E�C��,AC��Y|#����(
EA�J�pQd W3��T0 k� ����&�1D"3Q	24#Q  ��    ��� Y�TOD3/�Ip?��(AC��Y|#����$
EA�I�tRd$W3��T0 k� ������&�1D"3Q	24#Q  ��    ��� V�POD3/�Ip7��(AC��Y|#����
EA�G�tRd,V3��T0 k� ������&�1D"3Q	24#Q  ��    ��� S�HOD3/�Ip3��$@C��Y|#����
E1�F�xRd0U3��T0 k� ������&�1D"3Q	24#Q  �   ��� O�@OD3/�Ip'�� @C��Y|#���"	E1�C��Rd8T3��T0 k� ������&�1D"3Q	24#Q ��    ��� K�<OD3/�Ip#�� @C��Y|#��"	E1|B��Rd<S3��T0 k� ������&�1D"3Q	24#Q ��    ��� G�<OEc/�I��� @C��Y|#��!�	E1t@��R4@R3��T0 k� ������&�1D"3Q	24#Q ��    ��� C�8OEc/�I���?C��Y|#��!�E1l?��Q4DR3��T0 k� ������&�1D"3Q	24#Q ��    ��� ?�8OEc/�I���>C��Y|#�ۢ!�E1d=��Q4HQ3��T0 k� ������&�1D"3Q	24#Q ��    ��� ;"0NEc+�I���>C��Y|#�ӡ!�E1`<��Q4LP3��T0 k� ������&�1D"3Q	24#Q ��    ��� 7"(NEc+�I���=C��Y|#�Ϡ1�E1X:��Q4PO3��T0 k� ������&�1D"3Q	24#Q ��    ��� 3" NES+�E@��<C��Y|#�ǟ1�E1P9��P4TN3��T0 k� ������&�1D"3Q	24#Q ��   ��� /"MES'�E@��;C��Y|#���1�E1L7��P4TM3��T0 k� ������&�1D"3Q	24#Q ��    ��� ,"MES'�EO���:C��Y|#���1�E1D5��O4XL3��T0 k� ������&�1D"3Q	24#Q ��    ��� )" LES�EO���9C���Y|#���1�E182��N4\J3��T0 k� �����&�1D"3Q	24#Q ��    ��� &!�LC��EO���8C���Y|#���A�E100��Md`I3��T0 k� �w��{�&�1D"3Q	24#Q ��    ��� #!�KC��EO��27D ��Y|#���A�E1,.��Md`H3��T0 k� �o��s�&�1D"3Q	24#Q ��    ���  !�KC��EO��2 6D ��Y|#���A�E1$-��Ld`G3��T0 k� �g��k�&�1D"3Q	24#Q ��    ��� !�KC��EO��2 5D �Y|#���A�E1 +��KddF3��T0 k� �_��c�&�1D"3Q	24#Q ��    ��� !�JC��EO��1�5D {�Y|#���A�CA)s�KddE3��T0 k� �W��[�&�1D"3Q	24#Q ��    ��� !�JES�E?��1�4D s�Y|#�{�A�CA's�JTdD3��T0 k� �O��S�&�1D"3Q	24#Q ��    ��� !�IES�E?��1�3D o�Y|#�w�A�CA%s�IThC3��T0 k� �G��K�&�1D"3Q	24#Q ��    ��� !�IES�E?��1�3D k�Y|#�o�A�CA#s�HThB3��T0 k� �?��C�&�1D"3Q	24#Q ��    ��� !�HER��E?��1�1D c�Y|#�_�A�C@� s�FTh@3��T0 k� �/��3�&�1D"3Q	24#Q ��    ��� !�HER��E?����1D [�Y|#��W�A�C@�s�E�h?3��T0 k� �'��+�&�1D"3Q	24#Q ��    ��� !�HER��E?����0D W�Y|#��O�A�E��s�D�h>3��T0 k� ����&�1D"3Q	24#Q ��    ��� !�HER��E?����0DO�Y|#��G�A�E��s�C�h=3��T0 k� ����&�1D"3Q	24#Q ��    ��� !�GEB��E?����/DK�Y|#��?�A�E��c�A�d<3��T0 k� ����&�1D"3Q	24#Q  ��    �����!�GEB��E?����/DC�Y|#��;�A|E��c�@�d;3��T0 k� ����&�1D"3Q	24#Q  ��    �����!�GEB��E?����/D?�Y|#�Q3�AxE��c�?�d:3��T0 k� ������&�1D"3Q	24#Q  /�    �����!�FEB��E/����.D7�Y|#�Q+�AtE��c�>�d93��T0 k� �����&�1D"3Q	24#Q  ��    �����!�FEB��E/����.D3�Y|#�Q#�ApE��c�=�`83��T0 k� ����&�1D"3Q	24#Q  ��    �����Q|EEB��E/����.D'�Y|#�Q�AhE��3�:�\63��T0 k� �۔�ߔ&�1D"3Q	24#Q  ��    �����QtEEB��E/����.D�Y|#�Q�AdE��
3�9�\5c��T0 k� �ې�ߐ&�1D"3Q	24#Q  ��    �����QpEEB��E/����.D�Y|#�A�A`E��3�7�X5c��T0 k� �א�ې&�1D"3Q	24#Q  ��    �����QhEC�� E/����.D�Y|#�@��Q\E��3�6�T4c��T0 k� �Ӑ�א&�1D"3Q	24#Q  ��    �����Q\DC��E/����-C��Y|#�@�QPE��3�3�P2c��T0 k� �ǐ�ː&�1D"3Q	24#Q  ��    �����QTDC��E�����-C�� Y|#�@�QLE��3�2�L1c��T0 k� ����Ð&�1D"3Q	24#Q  ��    �����QLCC��E����-C�� Y|#�@ہQHE���C�0�L1c��T0 k� ������&�1D"3Q	24#Q  ��    �����QDCC��E�{���-C��Y|#�@ӀQDE���C�/�H0c��T0 k� ������&�1D"3Q	24#Q  ��    �����Q<CC��E�w���-C��Y|#�@ˀQ<E���C�.�D/c��T0 k� ������&�1D"3Q	24#Q  ��    �����Q0BC�|E�o�Ѹ-C��Y|#�@��Q4E���C�+�<.c��T0 k� ������&�1D"3Q	24#Q  ��    ������(BC�tE�o��-C��Y|#���Q,E���C�)�8-c��T0 k� ������&�1D"3Q	24#Q  ��    ������ AC�pE�k��-C��Y|#���Q(E���C�(�4,c��T0 k� �{���&�1D"3Q	24#Q  ��    ������AC�hE�c��-C�Y|#���Q E���C�&0+c��T0 k� �o��s�&�1D"3Q	24#Q  ��    ������@C�`E�_��-C�Y|#���AE���C�$,+c��T0 k� �c��g�&�1D"3Q	24#Q  ��&    ������@C�XE�[��-C�Y|#���AE��C�#(*c��T0 k� �[��_�&�1D"3Q	24#Q  ��&    �����P�?C�LE�W��-C��Y|#��AE�s�C�  )c��T0 k� �G��K�&�1D"3Q	24#Q  ��&    �����P�?C�DE�S��-C��Y|#�w�A E�o�S�(3��T0 k� �?��C�&�1D"3Q	24#Q  ��&    �����P�>C�<E�O��-C��Y|#�o�@�E�g�S�'3��T0 k� �7��;�&�1D"3Q	24#Q  ��&    �����P�>C�4E�K��-C��Y|#�g�@�E�c�S�'3��T0 k� �/��3�&�1D"3Q	24#Q  ��&    �����P�=C�,E�K��-C�|Y|#�_�@�C�[�S�&3��T0 k� �'��+�&�1D"3Q	24#Q  ��&    �����P�=C�$E�G��x-C�tY|#�W���C�W�S�%3��T0 k� ���#�&�1D"3Q	24#Q  ��&    �����P�<C�E�C��t-C�lY|#� O���C�O�S�%3��T0 k� ����&�1D"3Q	24#Q  ��&    �����P�<C�E�C��l-C�dY|#� G���C�K�S�$3��T0 k� ����&�1D"3Q	24#Q  ��&    �����P�;C�E�?��`-C�TY|#� 7���C�;�S��#3��T0 k� ����&�1D"3Q	24#Q  ��&    �����P�;C��E�;��X-DL	Y|#� /���E�7�S��"3��T0 k� ������&�1D"3Q	24#Q  ��&    �����@�;C��E/;��P-DH	Y|#� '���E�/�S��"3��T0 k� �����&�1D"3Q	24#Q  ��&    �����@�:C��E/7��L-D@	Y|#� ���E�'�c��!3��T0 k� ����&�1D"3Q	24#Q  ��&    �����@�:C��E/7��D-D8
Y|#� ���E�#�c��!3��T0 k� ����&�1D"3Q	24#Q  ��&    �����@�:C��E/7��<,D0
Y|#� ���E��c�� 3��T0 k� �ۜ�ߜ&�1D"3Q	24#Q  ��&    �����@x:C��E/7��4,D(
Y|'� ���E��c��3��T0 k� �ӝ�ם&�1D"3Q	24#Q  ��&    �����@p9C�� E/3��,,D 
Y|'�/����E��c�	�3��T0 k� �˝�ϝ&�1D"3Q	24#Q  ��&    �����@`9C���E/3� ,DY|'�?���	E���c��3��T0 k� ������&�1D"3Q	24#Q  ��&    �����@T9C���E/3�,E_Y|'�?���	E���c��3��T0 k� ������&�1D"3Q	24#Q  ��&    �����@L9C���B�3�,E_ Y|'�?ߑ�|
E���c��3��T0 k� ������&�1D"3Q	24#Q  ��&    �����@D9C���B�3�,E^�Y|'�?ג�tE���c��3��T0 k� ������&�1D"3Q	24#Q  ��&    �����@<9C���B�3� ,E^�Y|'�?ϓ�lE���c��3��T0 k� ������&�1D"3Q	24#Q  ��&    �����049C���B�3� �,E^�Y|'��ǔ�dE���c��3��T0 k� ������&�1D"3Q	24#Q  ��&    �����0$:C���B�7� �,E^�Y|+�߷��TE���c��3��T0 k� ������&�1D"3Q	24#Q  ��&    �����0:C�{�B�7� �,E^�Y|+�߯��LE���c��3��T0 k� ������&�1D"3Q	24#Q  ��&    �����0:C�s�B�7� �,E^�Y|+�ߧ��DE��c��3��T0 k� �����&�1D"3Q	24#Q  ��&    �����0;C�k�B�?��,E^�Y|+�ߛ��<E��c��3��T0 k� �w��{�&�1D"3Q	24#Q  ��&    �����0;C�c�B�C��,E^�Y|+�ߓ��4E��c��3��T0 k� �o��s�&�1D"3Q	24#Q  ��&    �����O�<C�[�B�K��,EN�Y|+�ߋ��,Ec��3��T0 k� �g��k�&�1D"3Q	24#Q  ��&    �����O�<C�S�B�O��,EN�Y|+�߃��$Ec��3��T0 k� �_��c�&�1D"3Q	24#Q  ��&    �����O�=C�C�B�O��,EN�Y|+����E���c��3��T0 k� �S��W�&�1D"3Q	24#Q  �&    �����O�>C�;�O/K��,EN�Y|+��{�@E���c��3��T0 k� �S��W�&�1D"3Q	24#Q  ��&    �����O�?C�3�O/K��,EN�Y|+��{�@E�{�c��3��T0 k� �S��W�&�1D"3Q	24#Q  ��&    �����O�@C�+�O/K��,EN�Y|+��w�@ E�s�c��3��T0 k� �S��W�&�1D"3Q	24#Q  ��&    �����O�AC��O/K�x,ENtY|+��o�O�E�c�c��3��T0 k� �K��O�&�1D"3Q	24#Q  ��&    �����O�BC��O/K��p,ENlY�+��k�O�E�[�c��3��T0 k� �G��K�&�1D"3Q	24#Q  ��&    �����O�CC��O/G��d,ENdY�+��g�O�D�S�c��3��T0 k� �C��G�&�1D"3Q	24#Q  ��F    �����O�DC��O/G��\,E�\Y�+��c�O�D�K�c��3��T0 k� �?��C�&�1D"3Q	24#Q   �F    �����_�EC���O/G��T,E�TY�+��_�O�D�G�c��3��T0 k� �;��?�&�1D"3Q	24#Q  ��F    �����_�HC���O/G��D,E�DY�+��S�O�!D�7�c��3��T0 k� �3��7�&�1D"3Q	24#Q  ��F    �����_�IC���O/G�%�<,E�<Y�+��O�O�"D�3�c��3��T0 k� �/~�3~&�1D"3Q	24#Q  ��F    �����_�JC���O/C�%�4,E�4Y�+��K�?�#E�+�c��3��T0 k� �+}�/}&�1D"3Q	24#Q  ��F    �����	_�KC���O/C�%�,,E�,Y�+��G�?�$E�#�c��3��T0 k� �#|�'|&�1D"3Q	24#Q  ��F    �����	_�MC���O/C�%�$,E�$Y�+��?�?�%E��c��3��T0 k� �{�#{&�1D"3Q	24#Q  ��F    �����	_|NC���O/C�%�,E�Y�+��;�?�&E��c��3��T0 k� �z�z&�1D"3Q	24#Q  ��F    �����	_pPC���O/C�%�,E�Y�+��/�?�(E��c��3��T0 k� �|�|&�1D"3Q	24#Q  ��F    �����	_lQC���O/?�%�,E�Y�+��+�?�*E��c��3��T0 k� �}�}&�1D"3Q	24#Q  ��F    �����	ohRC���O/?�%��,E��Y�+��#�?�+E���c��3��T0 k� ��~��~&�1D"3Q	24#Q  ��F    �����	odSC���O/?�%��,E��Y�+���?|-E���c��3��T0 k� ����&�1D"3Q	24#Q  ��F    �����	o`SC���O/?�%��,E��Y�+���Ox.E���c��3��T0 k� ����&�1D"3Q	24#Q  ��F    �����	oXTC���O/?�%��,E��Y�+�_�Op/E���c��3��T0 k� ����&�1D"3Q	24#Q  ��F    �����	oXUC���O/;�%��,E��Y�+�_�Oh1F��c��3��T0 k� ����&�1D"3Q	24#Q  ��F    ����~	_TVC��O/;�%��,E��Y�+�_�Od2F��c��3��T0 k� �ߌ��&�1D"3Q	24#Q  ��F    ����|	_PVC�w�O/;�%��,E��Y�+�^��O\4F��c��3��T0 k� �ێ�ߎ&�1D"3Q	24#Q  ��F    ����z	_HXC�g�E�7�%��,E��Y�+�^�OP7F��c�|3��T0 k� �Ϗ�ӏ&�1D"3Q	24#Q  ��F    ����x	_DYC�c�E�7�%��,E�Y�+�^�OL9F��c�x3��T0 k� �Ǒ�ˑ&�1D"3Q	24#Q  ��F    ����u�@YC�[�E�7�%��,E�Y�+�^�OH:F��c�x3��T0 k� ����Ò&�1D"3Q	24#Q  ��F    ����s�8ZC�S�E�7�%��,E�Y�+�^ۍO@<F��c�t3��T0 k� ������&�1D"3Q	24#Q  ��F    ����p�4[C�K�E�7�%��,E�Y�+�^ӍO<=F��c�t3��T0 k� ������&�1D"3Q	24#Q  ��F    ����m�0\C�C�E�3�%��,E]�Y�+�^ˍO4?F��c�t3��T0 k� ������&�1D"3Q	24#Q  ��F    ����k�,]C�;�E�3�%��,E]�Y�+�NÍ_0AF��c�p3��T0 k� ������&�1D"3Q	24#Q  ��F    ����h�(^C�3�E�3�%��,E]�Y�+�N��_,BE���c�p3��T0 k� ������&�1D"3Q	24#Q  ��F    ����f�$_C�/�E�3�%��+E]�Y�+�N��_$DE���c�l3��T0 k� ������&�1D"3Q	24#Q  ��F    ����c�`C�'�E�/�%��+E]xY�+�N��_ FE���c�l3��T0 k� ������&�1D"3Q	24#Q  ��F    ����a�aC��E�/�%��+E]pY�+�N��_HE���c�l3��T0 k� �����&�1D"3Q	24#Q  ��F    ����^�bC��E�+�%��+E]hY�+�N��?IE���c��h3��T0 k� �w��{�&�1D"3Q	24#Q  ��F    ����[�dE��E�+�%�t+E]XY�+���?ME���c|�d3��T0 k� �_��c�&�1D"3Q	24#Q  ��F    ����X� eE��E�'�%�p+E]PY�+��?NE���c|�d3��T0 k� �O��S�&�1D"3Q	24#Q  ��F    ����V��fE���E�#�%�l+E]HY�+�w�?PE���cx�`3��T0 k� �C��G�&�1D"3Q	24#Q  ��F    ����T��gE���E�#��d+E]@Y�+�o�? RE���Sx�\3��T0 k� �7��;�&�1D"3Q	24#Q  ��F    ����R��gE���E���`+E]<Y�+�g�>�TE���St�\3��T0 k� �/��3�&�1D"3Q	24#Q  ��F    ����P��hE���E���X+E]4
Y�+�_�.�VE���Sp�X3��T0 k� �'��+�&�1D"3Q	24#Q  ��F    ����N��iE���E���T+E],
Y�+�W�.�XE���Sp�T3��T0 k� ���#�&�1D"3Q	24#Q  ��F    ����L��jE���E���L+EM$
Y�+�K�.�YE���Sl �P3��T0 k� ����&�1D"3Q	24#Q  ��F    ����J��lE���E���@+EM
Y�+�;�.�]E����d �L3��T0 k� ����&�1D"3Q	24#Q  ��&    ����H��mC��E_��<+EM
Y�+�3���]E����` �H3��T0 k� ����&�1D"3Q	24#Q  �&    ����G��nC��E_��4+EM
Y�+�n+���_E����c��D3��T0 k� �����&�1D"3Q	24#Q ��/    ����F�oC��E_��,+EL�
Y�+�n#���`@����_��@3��T0 k� ������&�1D"3Q	24#Q ��/    ����E�pC��E^���(+EL�
Y�+�n���a@����[��83��T0 k� ������&�1D"3Q	24#Q �/    ����E^�qCE^��_ +EL�
Y�+�n���c@����W��43��T0 k� ������&�1D"3Q	24#Q �/    ����E^�sA_��E^�_+EL�	Y�+�n�	^�e@����K��,3��T0 k� �����&�1D"3Q	24#Q ��/    ����E^�tA_��E^�_+EL�	Y�+�]��	^�fE����G��(3��T0 k� �����&�1D"3Q	24#Q ��/    ����E^�uA_�E^�_+EL�	Y�+�]�	^�gE����C��$3��T0 k� ����&�1D"3Q	24#Q ��/    ����E^�vA_w�I�߆_ +EL�	Y�+�]�	^�iE����?��3��T0 k� ������&�1D"3Q	24#Q ��/    ����E^|wA_s�I�ۅ^�+EL�	Y�+�]�	^�jE����;��3��T0 k� ������&�1D"3Q	24#Q ��/    ����E^xwA_k�I�Ӆ^�+EL�	Y�+�]ߔ	n�kE����3�3��T0 k� ������&�1D"3Q	24#Q ��/    ����E^pxA_c�I�τ^�+A�Y�+�Mה	n�kEο��/�3��T0 k� ������&�1D"3Q	24#Q ��/    ����E^hyA_[�I�˄^�+A�Y�+�Mӕ	n�lEο��'�3��T0 k� ������&�1D"3Q	24#Q ��/   ����E^dzA_W�I�ǃ^�+A�Y�+�M˕	n�mEο��#� 3��T0 k� ������&�1D"3Q	24#Q ��/    ����E^\{A_O�I�Ã^�+A�Y�+�MÕ	n�nEο����3��T0 k� ������&�1D"3Q	24#Q	 ��/    ����E^X|A_K�I���^�+A�Y�+�M��	^�oEο����3��T0 k� ������&�1D"3Q	24#Q	 ��/    ����E^P}A_C�I���^�+A�Y�+�M��	^�oC������3��T0 k� ������&�1D"3Q	24#Q	 ��/    ����E^L~A_;�I���^�+A�Y�+�M��	^�pC������3��T0 k� ������&�1D"3Q	24#Q
 ��/    ����E^D~A_7�I���^�+A�Y�+�M��	^�qC������3��T0 k� ������&�1D"3Q	24#Q
 ��/   ����E^@A_/�I���^�+A|Y�+�M��	^�rC������3��T0 k� ������&�1D"3Q	24#Q
 ��/    ����E^8�A_+�I���^�+Axa�+�M����rC������"���T0 k� ������&�1D"3Q	24#Q
 ��/    ����E^4�A_#�I���^�+Apa�+�M����sC������"���T0 k� ������&�1D"3Q	24#Q
 ��/    ����E^,A_�I���^�+Ala�+�M����sC������"���T0 k� ������&�1D"3Q	24#Q ��/    ����E^(A_�I���^�+Ada�+�M����sC������"���T0 k� ������&�1D"3Q	24#Q ��/    ����E^$A_�I���^�+A`a�+�M����rC������"���T0 k� ������&�1D"3Q	24#Q ��/    ����E^A_�I���^�+AXa�+�M���rC������"���T0 k� ������&�1D"3Q	24#Q ��/    ����E^~A_�I���^�+ATa�+�M{���rC������"���T0 k� ������&�1D"3Q	24#Q ��/    ����E^~A_�I���^�+APa�+�Mw���rC������"���T0 k� ����&�1D"3Q	24#Q ��/    ����E^~A^��I���^�+AHa�+�Mo���qC������"���T0 k� ����&�1D"3Q	24#Q ��/    ����E^~A^��I���^�+ADa�+�Mk���qC������"���T0 k� ��	��	&�1D"3Q	24#Q ��/    ����E^~A^�I���^�+A@a�+�Mg���qC������"���T0 k� ����&�1D"3Q	24#Q ��/    ����E^ }A^�I���^�+A8Y�+�M_���qC������3��T0 k� ����&�1D"3Q	24#Q ��/   ����E]�}A^�I���^�+A4Y�+�	}[���qC������|3��T0 k� ����&�1D"3Q	24#Q ��/    ����E]�}A^�I���^�+A0Y�+�	}W���pC������t3��T0 k� ����&�1D"3Q	24#Q ��/    ����E]�}A^ߩI���^x+A,Y�+�	}S��|pC������l3��T0 k� ����&�1D"3Q	24#Q ��/    ����E]�|A^ۨI���^t+A(Y�+�	}O��xpC������`3��T0 k� ����&�1D"3Q	24#Q
 ��/    ����E]�|A^קI���^p+A Y�+�	}K��ppC������X3��T0 k� ��!��!&�1D"3Q	24#Q
 ��/    ����E]�|A^ӧI���^l+AY�+�	}G��loC���{��P3��T0 k� ��$��$&�1D"3Q	24#Q
 ��/    ����E]�|A^ϦI���^h+AY�+�	�C��hoC���s��H3��T0 k� ��(��(&�1D"3Q	24#Q
 ��/    ����E]�|A^˦A���^d+AY�+�	�?��doC��k��@3��T0 k� ��+��+&�1D"3Q	24#Q	 ��/    ����E]�|A^åA���^d+AY�+�	�;��`oC�{�c��83��T0 k� ��/��/&�1D"3Q	24#Q	 ��/    ����E]�{A^��A���^`+AY�+�	�;��XoC�w��[��03��T0 k� ��2��2&�1D"3Q	24#Q	 ��/    ����E]�{A^��A���^\+Aa�+�	�7��TnC�s��S��$"s��T0 k� ��6��6&�1D"3Q	24#Q ��/    ����E]�{A^��A���^X+Aa�+�	}3��PnC�o��K��"s��T0 k� ��9��9&�1D"3Q	24#Q ��/    ����E]�{A^��A���^T+Aa�+�	}3��LnC�k��C��"s��T0 k� ��<��<&�1D"3Q	24#Q ��/    ����E]�{A^��A���^P+Aa�+�	}/��HnC�c��;��"s��T0 k� ��@��@&�1D"3Q	24#Q ��/    ����E]�zA^��A���^L+Aa�+�	}/��DnC�_��3��"s��T0 k� ��C��C&�1D"3Q	24#Q ��/    ����E]�zA^��A���^H+Aa�+�	}+��@nC�[��+���"s��T0 k� ��G��G&�1D"3Q	24#Q ��/   ����E]�zA^��A���^D+Aa�+�	�+��<mC�S��#���"s��T0 k� ��J��J&�1D"3Q	24#Q ��    ����EM�zA^��A���^D+A a�+�	�'��8mC�O����"s��T0 k� ��N��N&�1D"3Q	24#Q ��    ����EM�zA^��A���^@+A a�/�	�'��4mC�K����"s��T0 k� ��Q��Q&�1D"3Q	24#Q ��    ����EM�yA^��A���^<+A�a�/�	�'�0mE�C����"s��T0 k� ��U��U&�1D"3Q	24#Q ��    ����EM�yA^��A���^8+A�a�/�	�'�,mE�?����"s��T0 k� ��X��X&�1D"3Q	24#Q ��    ����EM�yA^��A���^4+A�Y�/�	}#�(mE�7�����3��T0 k� ��[��[&�1D"3Q	24#Q ��    ����EM�yA^��A���^4+A�Y�/�	}#� nE�3�����3��T0 k� ��_��_&�1D"3Q	24#Q ��    ����EM�xA^��A���^0+A�Y�/�	}#�oE�/�����3��T0 k� ��b��b&�1D"3Q	24#Q ��    ����EM�xA^��A���^,+A�Y�/�	}#��oE�'�����3��T0 k� �|f��f&�1D"3Q	24#Q  ��    ����EM�xA^��A���^,+A��Y�/�	}#��pE������3��T0 k� �|i��i&�1D"3Q	24#Q  ��   ����EM�xA^��A���^(+A��Y�/�	�#�� qE������3��T0 k� �xm�|m&�1D"3Q	24#Q  ,�    ����E�wA^�A���^$+A��Y�/�	�#���rE������3��T0 k� �xp�|p&�1D"3Q	24#Q  ��    ����E�wA^{�A���^ +A��Y�/�	�#���sE������3��T0 k� �ts�xs&�1D"3Q	24#Q  ��    ����E�wA^w�A���^ +A��Y�/�	�#���tE�����3��T0 k� �tw�xw&�1D"3Q	24#Q ��    ����E�wA^s�A���^+A��Y�/�	�#���uE�����!�3��T0 k� �pz�tz&�1D"3Q	24#Q ��    ����E�vA^s�A���^+A��Y�3�#���vE�����!�3��T0 k� �l~�p~&�1D"3Q	24#Q ��    ����E�vA^o�A���^+A��Y�3�#���wC����!|3��T0 k� �l��p�&�1D"3Q	24#Q ��    ����E�vA^k�A���^+A��Y�3�#���wC����!t3��T0 k� �h��l�&�1D"3Q	24#Q (�    ����E|vA^g�A���^+A��Y�3�#���xC����!p3��T0 k� �h��l�&�1D"3Q	24#Q ��    ����ExvA^g�A���^+A��Y�3�#���yC�۶��!h3��T0 k� �`��d�&�1D"3Q	24#Q ��     ����ExuA^c�A���^+A��Y�3� �#���yC�ӵ��!d3��T0 k� �`��d�&�1D"3Q	24#Q ��     ����EtuA^_�A���^+A��Y�3� �#�͸zC�˳�!\3��T0 k� �\��`�&�1D"3Q	24#Q ��     ����EpuA^_�A���^+A��Y�3� �#�ʹ{C�òw�!X3��T0 k� �X��\�&�1D"3Q	24#Q ��     ����EltA^[�A���^+A��Y�3� �#�ͬzC�o�!P3��T0 k� �T��X�&�1D"3Q	24#Q ��     ����EhtA^W�A���^+A��Y�3� �#�ͨzC�g�!L3��T0 k� �P��T�&�1D"3Q	24#Q  ��     ����EdtA^W�A���^ +A��Y�3� �#�ͤzC���_�!D3��T0 k� �L��P�&�1D"3Q	24#Q  ��     ����E`tA^S�A���^ +A��Y�7� �#�͠zC���W�!@3��T0 k� �H��L�&�1D"3Q	24#Q  ��     ����E\sA^S�A���]�+A��Y�7� �#�͘yC���O�!83��T0 k� �D��H�&�1D"3Q	24#Q  ��     ����E                                                                                                                                                                            � � �  �  �  d A�  �K����   �      � \��B� ]�":"9 � �! `�3    �	  ���     `�����    ���#             
    ��         �     ���   0
&


         ��K          ��p    ��N�p,    ����                 	 ^ �         ��      ���   (
 
          ��RE          ��+    ��RE��+                          �         �     ���   0	
           +��           �`ho     +���`oy      ��   
                �$          �      ���   H	$
         ��E�        /� �    ��I�� �    ��                   �$          �p     ���   03 
          ��R+ ��     C��5    ��R+���       2                     ���u             )  ���   P		 5             ���  Q Q   W�9�%    ���g�9N�    ��               1		���E          ��       ��@   (
	           pU�   S	    k�(�     pW!�(�    ���               ���E          �     ��J   8	 

         ��g� � �	   �I�    ��v��IŜ    �<��             
	���E         ���     ��`   
	          ���  � �
   ��U?�    ��U��U>�    ���               o	���E         	 ��     ��`  0
3
         ���H  � �	    ���c    ��8)����    �/��              D ���E         
 ��    ��`   H


         ���  ��     � �Ρ    ���  �Ρ                            ���[               ��@    		 5 	                 ��      �                                                                           �                               ��        ���          ��                                                                 �                          m��  ��        ����     m�{���    ���# "                  x                j  �        �                          m    ��        ��       m  �           "                                                 �                         ��p���`���9�(�I�U�� �����    
      	       
  /   �] �L�B       � @o� ʄ  p` �� 0p� �$ @q  ˤ q� �� q� �D l� ɤ  v@ �� v����J ����X � '� d@ � �w` � 0x` �d  x� פ y  Z� x� ?� v   s@ 
�| W  
�\ W  
�< W� 
�� W� 
�\ X  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �D �Q����� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����E������ �  ������  
�fD
��L���"����D"� �  " `   J jF��    "�j "���
��
���     �j��  
  �
� �  �  
�  `    ��     ��       `    ��     ��       p    ��     ��(          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  � &&       ��t  ��        �t  ��        �        ��        �        ��        �    ��    ���� f�        ��                         T�) ,  �����                                      �                 ����              `� ���&��  ���E���� ;            35 Bob Essensa le                                                                                   4  4      �
"�b
�b'�$'�;K/3K7	 KC
KD" 	KJ

KK �	cW � �c] � �k � �k� � �k� � �k� � � k� � � k� � �c� � �c� � � c� � � c� � �c� � �C_ � C#g �J� � � J� � wK � � K � bc�# � c�) Y c� I!c�$ I "c�, }#* | �$!� | �%"9 � � &"F � � '"H �(* | )"Q �*" � +"G �,!� |=-"7 |E ."E �]  "D � � 0"J � 1"' �2"- |H 3"E �`  "S � �5"; � 6"Q �7!� �D8"+ |\ "= � z  "D t �;!� x <"K �W  "! x �>"* �  *J � 
�                                                                                                                                                                                                                 �� P        �     @ 
        �     _ P E a  ��                     ������������������������������������� ���������	�
���������                                                                                          ��    ��W�� ��������������������������������������������������������   �4, >    �@<�@��A�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     C    2    �� �:�J                                      ������������������������������������������������������                                                                                                                                             ����  ��                                             �������������������������� ����������� ��������� ��� ����� ��� ��� ������������� ����� ���� �� ����� �� ��� ������������� � �������� ���������� �������������������������� ����������� ���� ������� ���������������������������� ���                                    B   ! 2    �� �R�J      P  	                           ������������������������������������������������������                                                                                                                                         ����  �  �                                           ��� ����������������������������������������� ����������������� ��������� ���� ��������� ����������������������������� ���  �������������������������������� ��   ��� ��������������������������� ���� ��  ���������������������������� ������� � ��� �������                                                                                                                                                                                                                                                                                                                   	         �              


             �   }�         ���}  �  2�  �����  I��������������������������������������������������������������������������������      2�             R     [                                                      ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � �8�5 �\                                                                                                                                                                                                                                                                                            )n)nY  EE     r       k      l      k                        `                                                                                                                                                                                                                                                                                                                                                                                                        > �  >�  �  
�  � ��  J`�  ���Q����u��� u��H�S�̞�����������������0                      �� |        $   �   &  QW  �   �                    �                                                                                                                                                                                                                                                                                                                                        K K   �                      !��                                                                                                                                                                                                                            Z   �� �� Ѱ�      �� \      �������������������������� ����������� ��������� ��� ����� ��� ��� ������������� ����� ���� �� ����� �� ��� ������������� � �������� ���������� �������������������������� ����������� ���� ������� ���������������������������� ������ ����������������������������������������� ����������������� ��������� ���� ��������� ����������������������������� ���  �������������������������������� ��   ��� ��������������������������� ���� ��  ���������������������������� ������� � ��� �������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ?      @   �  m                       f     �  ���������J'      ��     F�   �      �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ��  � ��     � ��  � ��   p �� �� �z   p����  ��  �� ��  [� �� �� �z  [� � �$ ^$&  ��  ��   ��     ��  m �� �� �z  m�� ��  � ��  �� ��   ��  �� �� �  �� �� �z � ��� �$  � �  �� �  �      �       !���� e����� g���       f ^�         �� c��      !      ��B����2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                                                  U  T   T   T     T UDUDDUDDDDDDDDDDDDDDDP   E�  DU� DDU�DDDUDDDDDDDDDDDD                UP  E�  E   E                                           ���U�UTD�DDDDDDTDD TDD   �   U_ DEU�DDDUDDDDD��DZT�DDDDDDDDDDDDTDDDDDDDDUTU�����DDDDDDDDDDDEDDDEDDDDTUTU�Ԫ���Z_   P   � �U�UTDUDDDDUTD�DT��D        U_��DEU_DDD_DDDPDDE�DDE  �DD DD DD �DD �UD  �U       DZTDEDDDDE�DDE�DDE�TDDT�DE�TE���DDTU�ZD���������DDTDD��ZT�T���ZTDDE��D��T�T��DUTTT��Z��TQTDDUTD�DDDTDDD�DDDDDDE�DD_TDE�DD_ DDP DDP DD_ DU_ U�  �                                       TE�DDD�UUU                    ���DDDUUUTD  D  D  D  D  U��D�TDDDDEUUDP  DP  DP  DP  UP  TDE�DDDPUUU_                                                    wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwtwwwCwwt1wwCwt1wC�t1��C1����������""""���������������!���""!����,���ww��7����������������wwwwwwwwwwwwwwwwwwww7wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwws��w1wt1�wC�t1��s��s��s������"$��Gw�!������������L���q��"r��������!�����!ww�r�w�ww!�wwrwwwwwwqwwwrwwww�7ww�ww�ww��7w��w���G��'!wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                                    �����   �   �   �   ����                                     	�  		  	 � 	 	 	   	   	   	   	  ��                  ��   	   	   	   	   	   	 	 	 � 		  	�                 �   	    �   	    �   	    �   	   	   �  	   �  	   �  	   �                                                       �����   �   �   �   ����                                     
�  

  
 � 
 
 
   
   
   
   
  ��                  ��   
   
   
   
   
   
 
 
 � 

  
�                 �   
    �   
    �   
    �   
   
   �  
   �  
   �  
   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    "!  "" "  """ ""   "! " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ ""   "! " ""  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """ "!    " ""            """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                 �   �  
� 
�� ���	���    �   ��  ��  �ڠ bj� gj��w���������������˽,̲" �""  "  
�  
�   �   �   J   
           ����̻ۻ�˽��˽�̻��뻽���K���RDD>�UD4NUDD�T4�K 3˸ Ȣ   "" �   �   �   �   �   �   "   "   "   "   ".  C � ;� �ˊ  ��  
�"  0  0 2#  3 "# 0 0     " �/����      �             "�"�����   �� �          ����   �       �                                   �    ��"  �"                    ".  ".  ���   ��                                 � "�"  �    � � �                                                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��  ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  &'  vv  w                �                        ��"� �"� ����        �   �   �"  �""��� �   �     �   "  "  "   �                                                                                                                                                                             �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���        �/  ��  �                          �   � � /  �"" �"  �       �    � �  �                     �         "   "   �       �   �   �   D   E�  U�  UO                         "  "  "      � "�"  �    � � �                                                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��                        �          �   � � /  �"" �"  �                     � �� ���H���     ̰ �˻���ݹ��w���&ɧvvɪ�p              �  "� "� "/ "�                         ����                               ���                          ����                  �   �� �       �  �  "�  "   "                                                          �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp��& ��vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �" �"" �"   �                    .   .   �                   �   ��  �ڛ�}ک�"   "   "  �� ��                   �".��".���                   �  �  �  �               �   ��  ���   �                 ���������������������  ��  ��  ��  �   �    �          �         �                                �  �  "�  "   "                                                            �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �      �              �   �                                    �  .   .     �   �  ��  �                                                                                                                    �  �  "   "                                                                    �U  EU  U  3 � �   �  �   �   �   �                   U�  U�@ EZ� 4Z� 3ZS U� E����" ��� 
��  �" ""�"" �"!  �  �                        "  "/  "��� "  !��  ���  �       �  ��  ̽  ��  �w  �� 
�� ��� ��� ��� ��� ��� ��� ��� �� ���    �   �   �   �   �   ˰  ˙  ɪ  ��� ټ� �̰ �̰ ��� ��  ��     �                                                                            �               �     "   "                   ��   �  ��  �  �  �         � ".��".��/����  �                                                                                                                                         	�  �� �� ���ܙܽɪ�͚�����͙ͼ̨��̄DC"�D32�C33�333�33P330X̽ 
�� ˪  "   ""/"""�����vv ��p ��  ��  ̽  ˸  ɚ  ��  ؛  -�� .ܰ .��  �"  �   .   "�                   � �  ��            Z   Z   Z   Z  Z  �� �� �� "� "" "" ""/ ����   �   � .�". �" ����                    �� ��������p��r`  .  " "" ��� "                       �   �    �                                                                       � ��       "   "   "�  �                            �   ���                            �   "                                                                                                      �  ��� ݻ� g�� bm� ggz�'w���������������˛������ˊۼ�����˻������H�DH�@U�DPT�E X�T H�P H�@ Ȥ� ̻� ˘ "�� � ���/�"" �""/���               �   �                                                     �  �                      � �                       ���           �                      "  "             ��.�  .                 ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                               ���                          ����                  �   �� �       �  �  "�  "   "                                            �w
���̩ۚ,���+��   �   �   �   �  �  9  D3  D2 T2 DB DB �@ ��  ��  ��  �  "" ""�"!��" ��       �                w�  ��� ��� ��� ˼����ɀ�؊�˽ـ��˰��̰�̻@"���"+H�"$X�"$�@"E� U� E� D� ,˸  ��  ��  ,� "" �"" """�"!���� � �              �         �           �       �                                      "  ."  �"    �          �� ̻� ��� ww� &'� vvw    �   �     �     �  �  "   "   "   "�  �                                  ���                                                                                                                                                                             �  �� �� wȠb���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 " "" "  �   �   �           �   �   �           �  "�  "                                       ����                               ���                          ����                  �   �� �       �  �  "�  "   "                                                                    �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ���������""��""��""�����        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                                               �         �  "� "  �  ��                                                                                                                                                 2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�GwDGwqwDDwtwwww3333DDDD �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�""""����������A��I��I = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=""""�����A�DA�I��I�    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"��������I���I���I���I��� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(XxMAMAMMMM�M�M����3333DDDD w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xwwD�����MD��M����3333DDDD  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���4���4���4���4���4���43334DDDD �  + � � � � � � � � � � ��	� � � ��� � � � � � � � � � � ��	� � � ��� �� ����(+((�""""wwwwqqqqwGwGGG ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""wwwwwwqqDAwG M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M������������������333DDD � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�M��M��D��M����������3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DD��D�M��D����3333DDDD 5 6  X � �F � � � � � ����� � ����������� � ����� � � � � ��	F ��(X((6(5""""wwwwwwDGqGq x �  l � �G � � � � � � � � � � ������������� � � � � � � � � � ��	G ��l((�x""""wwwwwwwGqGqqD w w x y ������H���������������������������������H�����yxww""""wwwwwwwwGwwGwwGwwGw  � + w�������I�J�K�L�M�N�O � � � � � � � � � � � � � � � � � � � ��O�N�M�L�K�J�I������w(+�(DDwwwqwwGwtDGwwww3333DDDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A e ��A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,GwAqAADqtDGwwwww3333DDDD +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�] � ځ]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+www4www4www4Gww4Gww4www43334DDDD 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U �h�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5""""���������M�MMM =  U ,     !d�P���e�f�g�!�!�!�k�!�!�!�l�!�!�!�!�k�!�!�!�l�!�!�!�g�f�e���P)d((( ((,(U((=""""�������A��AA     =  U , N ,�-�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�-(,(N(,(U((=((( ��������������333DDD � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � �I��I����������������3333DDDD  � �!�AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((���A���I��I���I�����3333DDDD m � �!�A�A� � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""������������������������  � �!�AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M""""������D�D��� 
 � �!�AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�""""������������������������ - � �!�!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�wqwwqwwwwwqwwwDwwww3333DDDD 69�:���  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5qqwwwDDwtGwwww3333DDDD x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xwww4www4www4www4www4www43334DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwqwwwqwqwq + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""wwwwwwwDwGwA � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(��A�L�L�L��L���333DDDLDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDD
"�b
�b'�$'�;K/3K7	 KC
KD" 	KJ

KK �	cW � �c] � �k � �k� � �k� � �k� � � k� � � k� � �c� � �c� � � c� � � c� � �c� � �C_ � C#g �J� � � J� � wK � � K � bc�# � c�) Y c� I!c�$ I "c�, }#* | �$!� | �%"9 � � &"F � � '"H �(* | )"Q �*" � +"G �,!� |=-"7 |E ."E �]  "D � � 0"J � 1"' �2"- |H 3"E �`  "S � �5"; � 6"Q �7!� �D8"+ |\ "= � z  "D t �;!� x <"K �W  "! x �>"* �  *J3333DDDDAqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD��������������������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ��������������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ��������������������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE��������������������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD��������������������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD��������������������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD��������������������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� ��%��:�L�S�S�L��0�R�S�\�U�K���������8�>�7���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� ����7�\�J��<�V�I�P�[�H�P�S�S�L�������8�>�7���""""������A�D��I��""""�������D����� ��!��-�V�I��0�Z�Z�L�U�Z�H����������8�>�7���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �8�>�7��� ���A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �>��<�����""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,�����������DDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �����<�L�Z�\�T�L��2�H�T�L����������������� ����4�U�Z�[�H�U�[��<�L�W�S�H�`��������������� ����.�O�H�U�N�L��2�V�H�S�P�L���������������� ������0�K�P�[��7�P�U�L�Z���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            