GST@�                                                           @c�                                                      W��       �  d   %   	      ����e ����ʱ����������X�������        Vi     #    ����                                d8<n    �  ?     b_����  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    B�jl �   B ��
                                                                                 ����������������������������������      ��    oo? 0 go5  8  +     '         ��  
    
          	� 74 V 	�                 �Y          8::�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             $F  ")          == �����������������������������������������������������������������������������                                �7  7       t�   @  #   �   �                                                                                '     �Y  "$)F    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    CO�/_��A�  8#�C�|( @`+�A (1�< @��P�#AP� T0 k� �| �� %�0d  e1�� Bb  ��/    �   CO�._��A�  o8#?C�|( @`+�A (1�< @�� �#AP� T0 k� �t �x %�0d  e1�� Bb  ��/    �   CO�._��A�  o8#?G�|, @`+�C�(1�< @�� �#AP� T0 k� �l �p %�0d  e1�� Bb  ��/    �   E��-_��A�  o8#?G�!�, @`+�C�$0�< 0�� �#J�� T0 k� �c��g�%�0d  e1�� Bb  ��D    �   E��,_��A�  o8#?G�!�, @`+�C�$0�< 0�� �#J�� T0 k� �c��g�%�0d  e1�� Bb  ��D    �   E��,?��C��  o8#?K�!�, @�+�C�$/�< 0�� �#J�� T0 k� �c��g�%�0d  e1�� Bb  ��D    �   E��+?��C��  �8#?K�!�, @�+�C� /�< 0�� ��#J�� T0 k� �g��k�%�0d  e1�� Bb  ��D    �   E��*?��C��  �8#OK�!�, @�+�C� /�< 0�� ��#J�� T0 k� �k��o�%�0d  e1�� Bb  ��D    �   E��)?��C��  �8#OO�!�, @�+�C� .p<  �� ��#J�� T0 k� �o��s�%�0d  e1�� Bb  ��D    �   E��(?��C��  �8#OO�!�, @�+�C�.p<  �� ��#J�� T0 k� �w��{�%�0d  e1�� Bb  ��D    �   E��'?��A��  �8#OO�!�, C�+�C�-p<  �� ��#J�� T0 k� �w��{�%�0d  e1�� Bb  ��D    �   E��&?��A��  �8#OS�!�, C�'�C�,p<  �� `�#J�� T0 k� �{���%�0d  e1�� Bb  ��D    �   E��%?��A�� 8#OS�!�, C�'�C�,p<  �� `�#J�� T0 k� �����%�0d  e1�� Bb  ��D    �   E��$?��A�� 8#OS�!�, C�'�C�+ < ��� `�#J�  T0 k� �����%�0d  e1�� Bb  ��D    �   E��$���A�� 8#OW�|, C�'�C�* < ��� `�#J�  T0 k� �����%�0d  e1�� Bb  ��D    �   E��#���A�� 8#OW�|, A '�E0) < ��� `�#J� T0 k� ������%�0d  e1�� Bb  ��D    �   E��"���A�� 8$?W�|, A #�E0) < ��� `�$J� T0 k� �����%�0d  e1�� Bb  ��D    �   E�� ���A�� O8$?[�|, A #�E0'P<  �� `�$J� T0 k� �{���%�0d  e1�� Bb  ��D    �   E�����A�� O8$?[�|, A #�E0&P<  �� `�$J� T0 k� �{���%�0d  e1�� Bb  ��D    �   E�����BO� O8%?[�|, E��E0%P<  �� �%J� T0 k� �w��{�%�0d  e1�� Bb  ��D    �   E�����BO� O8%�_�|, E��E $P<  �� �%J� T0 k� �w��{�%�0d  e1�� Bb  ��D    �   E�����BO� O8&�_�|, E��E $P8  �� �%J� T0 k� �{���%�0d  e1�� Bb  ��D    �   	E�����BO� O8'�c�|, E��E "�8 �� �&J� T0 k� �{���%�0d  e1�� Bb  ��D    �   
E�����@� O4'�c�|, E��E !�4 ���&J� T0 k� �����%�0d  e1�� Bb  ��D    �   E�����@� O4(�g�|, E��E  �4 ���&J� T0 k� �s��w�%�0d  e1�� Bb  ��D    �   E�����@� �4)�g�|, E��E �4 ���&J� T0 k� �o��s�%�0d  e1�� Bb  ��D    �   E����@� �4*�k�|, E��E �, ���'J� T0 k� �k��o�%�0d  e1�� Bb  ��D    �   E����B�� �4+�k�|, E��E �, ����'J�T0 k� �g��k�%�0d  e1�� Bb  ��D    �   E����B�� �0,�o�|, E���E �( ����'J�T0 k� �c��g�%�0d  e1�� Bb  ��D    �   E����B�� �0,�o�|, E���E�$ �����'J�T0 k� �c��g�%�0d  e1�� Bb  ��D    �   E����B�� �0-�o�|, E���E�  �����'J�T0 k� �` �d %�0d  e1�� Bb  ��D    �   E����B�� �,/�s�|, E���E� �����'J�T0 k� �` �d %�0d  e1�� Bb  ��D    �   E����B�� �,0�s�|, D?��E� �����'J�T0 k� �\ �` %�0d  e1�� Bb  ��D    �   E����B�� �(1�w�|, D?��J@� �����'J�T0 k� �` �d %�0d  e1�� Bb  ��D    �   E����B�� �$2�w�|, D?��J@� �����'J�T0 k� �` �d %�0d  e1�� Bb  ��D    �   E����B�� � 3�w�|, D?��J@ � ����&J�T0 k� �`�d%�0d  e1�� Bb  ��D    �   E�����B�� �4�w�|, E_��J@$� ����&J�T0 k� �`�d%�0d  e1�� Bb  ��D    �   E�����B�� �5�w�|, E_��E0$� ����&J�T0 k� �`�d%�0d  e1�� Bb  ��D    �   A_����B�� �6�w�|, E_��E0$P ����&J�T0 k� �`�d%�0d  e1�� Bb  ��D    �   A_����B�� �6�w�|, E_��E0(P ���%J�T0 k� �`�d%�0d  e1�� Bb  ��D    �   A_����B�� �7�w�|, E_��E0(P����%J�T0 k� �`�d%�0d  e1�� Bb  ��D    �   A_����B�� �9�w�|, E_��E�(P���� $J�T0 k� �`	�d	%�0d  e1�� Bb  ��D    �   A_����B�� �9�w�|, E_��E�,@����$$J�T0 k� �X�\%�0d  e1�� Bb  ��D    �   A�����B�� � :�s�|, E_��E�,@����(#J�T0 k� �T�X%�0d  e1�� Bb  ��D    �   A�����B�� ��;�s�|, E_��E�,@����,#J�T0 k� �T�X%�0d  e1�� Bb  ��D    �   A�����B�� ��<�l|, EO��E�0@���4"J�T0 k� �P�T%�0d  e1�� Bb  ��D    �   A�����B�� ��=ol|, EO��E�0p���8!J� T0 k� �@�D%�0d  e1�� Bb  ��D    �   A�����B�� ��=oh|, EO��E�0p���<!J� T0 k� �0�4%�0d  e1�� Bb  �D    �   
A���àQ� ��>oh|, EO��E�4p��#�@ J� T0 k� �$�(%�0d  e1�� Bb  ��D    �   	A���ǞQ� ��?od|, EO�E�4p��#�D J� T0 k� � �$%�0d  e1�� Bb  ��D    �   A���ϜQ� ��@�`|, EOo�E�4���+�H J�$T0 k� � �$%�0d  e1�� Bb  ��D    �   A���ӛQ� ��A�\|, EOg�E�4���/�L J�(T0 k� �$�(%�0d  e1�� Bb  ��D    �   A���ךQ� �A�X	|, EOc�E�4���/��PJ�(T0 k� �(�,%�0d  e1�� Bb  ��D    �   A���ߙQ� �B�T
|, EO[�E�4
���3��TJ�,T0 k� �(�,%�0d  e1�� Bb  ��D    �   A����Q� �C�L|, EOK�E�4
���;��XJ�0T0 k� �$
�(
%�0d  e1�� Bb  ��D    �   A����Q/� �D�H|, EOC�P�4
���?��\J�0T0 k� � �$%�0d  e1�� Bb  ��D    �  ��A����Q/� �D�D|, E??�P�4
p��C��\ J�4T0 k� �� %�0d  e1�� Bb  ��D    �  ��A�����Q/� �E�@|, E?7�P�4	p��C��` J�4T0 k� ��%�0d  e1�� Bb  ��D    �  ��A�����Q/� �E�<|, E?/�P�4	p��C��d J�8T0 k� �	�	%�0d  e1�� Bb  ��D    �  ��A����Q/� �F�8|, E?'�P�4p��G��d J�8T0 k� ��%�0d  e1�� Bb  ��D    �  ��A����Q/� �G�,|, E��P�0p��O��l!J�<T0 k� ��%�0d  e1�� Bb  ��D    �  ��A����Q?� xH�(|, E��P�0@��S��l!J�<T0 k� ��%�0d  e1�� Bb  ��D    �  ��D?���Q?� pH_$|, E��P�0@��W��p!J�<T0 k� � 
�
%�0d  e1�� Bb  ��D    �  ��D?��#�Q?� hI_|, E��P�0@�
�[��t"J�@T0 k� ��� %�0d  e1�� Bb  ��D    �  ��D?��+�Q?� `I_|, E���P�0@�
�c��x"J�@T0 k� ����%�0d  e1�� Bb  ��D    �  ��D?��7�Q?� PJ_|, E��P�,@�
�k�р#J�@T0 k� ����%�0d  e1�� Bb  ��D    �  ��D?��?�Q?� HK_|, E��P�,@�
�o�ф$J�@T0 k� ����%�0d  e1�� Bb  ��D    �  ��D?��G�Q?� @Ko |, E��P�, ��
�s�ш$J�DT0 k� ����%�0d  e1�� Bb  ��D    �  ��D?��K�Q?� 8Ln�|, E�ۺP�, ��
�{�ь$J�DT0 k� ����%�0d  e1�� Bb  ��D    �  ��DO��S�Q?� 0Ln�|, E�ӹP�, ��
��ѐ%J�HT0 k� ����%�0d  e1�� Bb  ��D    �  ��DO��c�Q?� Mn�|,E�ǷP�, ��
ы�ј&J�LT0 k� ����%�0d  e1�� Bb  ��D    �  ��DO��k�Q?��Nn�|,Eο�P�, ��
я�
ќ&J�LT0 k� ����%�0d  e1�� Bb  ��D    �  ��DO��s�Q?��Nn�|,E޷�P�, `�
ѓ�
Ѡ&J�PT0 k� ����%�0d  e1�� Bb  ��D    �  ��DO��w�Q?��N��|,Eޯ�A�, `�
��
Ѩ'J�TT0 k� ����%�0d  e1�� Bb  ��D    �  ��DO���Q?��O��|,Eޫ�A�, `�
��
Ѭ'J�TT0 k� ����%�0d  e1�� Bb  ��D    �  ��DO����Q?���P�|,Eޛ�A�, `�
��
Ѹ(J�\T0 k� ����%�0d  e1�� Bb  ��D    �  ��DO� ���Q?���P�|,CA�, `�
��
Ѽ(J�`T0 k� ����%�0d  e1�� Bb  ��D    �  ��DO�!���Q?���Q� |,CA�, `�
��
��(J�dT0 k� ����%�0d  e1�� Bb  ��D    �  ��D_�!���Q?���Q� |,CAP,�
��
��)E�hT0 k� ����%�0d  e1�� Bb  ��D    �  ��D_�"���Q?���Q� |,C��AP,�
���
��)E�lT0 k� �|��%�0d  e1�� Bb  ��D    �  ��D_�#���Q?���R�!|,C�w�AP,�
���
��)E�pT0 k� �t�x%�0d  e1�� Bb  ��D    �  ��D_�$���Q?���R�!|,E�o�AP(�
���
��*E�tT0 k� �l�p%�0d  e1�� Bb  ��D    �  ��D_�%���Q?���S�!|,E�g�AP(�
���
��*E�xT0 k� �d�h%�0d  e1�� Bb  ��D    �  ��D_�'�ˊQ?���S�x!|,E�[�C�(
p�
���
��+E��T0 k� �T�X%�0d  e1�� Bb  ��D    �  ��D_�(�ӋQ?���T�p"|,E�S�C�(
p�
���
��+E��T0 k� �L�P%�0d  e1�� Bb  ��D    �  ��D_�)�׋Q?���T�h"|,E�K�C�$
p�
���
��+E��T0 k� �D�H%�0d  e1�� Bb  ��D    �  ��D_�*�ߌQ?�ݔU�`"|,E�C�C�$
p�
���
� ,E��T0 k� �<�@%�0d  e1�� Bb  ��D    �  ��D_|+��Q?�݌U�X!|,E�;�C� 
p�
��
�,E��T0 k� �4�8%�0d  e1�� Bb  ��D    �  ��Dox,��Q?�݄U�P!|,E�7�C� 
��
��
�,A�T0 k� �,�0%�0d  e1�� Bb  ��D    �  ��Dot-��Q?��|V�H!|,E�/�C� 
��
��
�-A�T0 k� �$�(%�0d  e1�� Bb  ��D    �  ��Dop.��Q?��tV�@!|,E�'�C� 
��
��
�-A�T0 k� �
� 
%�0d  e1�� Bb  ��D    �  ��Dod1���Q?��dW�0!|,E��C�
��
�'�
�,-A�T0 k� �
�
%�0d  e1�� Bb  ��D    �  ��Do`2���Q?��\W�( |,E��C�
��
�/�
�0.A�T0 k� �
� 
%�0d  e1�� Bb  ��D    �  ��Do\3��Q?��TW�  |,E��C�
��
�7�
�8.A�T0 k� �	� 	%�0d  e1�� Bb  ��D    �  ��DoT5��Q?��LX�|,E���C�
��
�?�
�@.A�T0 k� �	�	%�0d  e1�� Bb  ��D    �  ��DoP6��Q?��DX�|,E���C�	
��
�G�
�H/A�T0 k� ��%�0d  e1�� Bb  ��D    �  ��DoL7��Q?��<X�|,E��C�	
��
�O�
�P/A�T0 k� ��%�0d  e1�� Bb  ��D    �  ��DoH8��Q?��4X�|,E��C�	
��RW�
�X/A�T0 k� ��%�0d  e1�� Bb  ��D    �  ��D?@:��Q?��,X��|,E��C� 	
��R_�
�`/A�T0 k� ��%�0d  e1�� Bb  ��D    �  ��D?<;��Q?��$Y��|,A�ۣC� 	
��Rc�
�h0A�T0 k� � �%�0d  e1�� Bb  ��D    �  ��D?4=��Q?��Y��|,A�ӢD  

��Rk�
�p0A�T0 k� ��� %�0d  e1�� Bb  ��D    �  ��D?0>��Q?��Y��|,A�ˢD�

��Rs�
�x0A�T0 k� ����%�0d  e1�� Bb  ��D    �  ��D?,?��Q?��Y�|,A�âD�

��Rw�
Ҁ0A�T0 k� ����%�0d  e1�� Bb  ��D    �  ��D? B��Q?���Y�|,P���D�
��R��
�1A�T0 k� ����%�0d  e1�� Bb  ��D    �  ��D?D��Q?�<�Y�|,P���D�
�#�R��
�1A�T0 k� ����%�0d  e1�� Bb  ��D    �  ��D?E��Q?�<�Y�|,P���D�
�'�R��
�1A�T0 k� ����%�0d  e1�� Bb  ��D    �  ��I�F��Q?�<�X�|,P���D�
�+�R��
�1A�T0 k� ����%�0d  e1�� Bb  ��D    �  ��I�H��Q?�<�X�|,P���D�
�/���
�2JѼT0 k� ����%�0d  e1�� Bb  ��D    �  ��I�I��Q?�<�X�|,P���D�
�/����2JѼT0 k� ����%�0d  e1�� Bb  ��D    �  ��I� J��Q?���X�|,P͋�D�
�7����2JѼT0 k� ����%�0d  e1�� Bb  ��D    �  ��I��K��Q?���X�|,P͇�D�
�;�����2J��T0 k� ����%�0d  e1�� Bb  ��D   �  ��I��L��Q?��W�|,P��D�
�?�����2J��T0 k� �� �� %�0d  e1�� Bb  ��D    �  ��I��M��Q?��W�|,P�{�D�
�C�����3J��T0 k� ������%�0d  e1�� Bb  ��D    �  ��I��N��Q?��W�|,P�s�D�
�G�����3J��T0 k� ������%�0d  e1�� Bb  ��D    �  ��I��O��Q?��W�|,P�o�D�
�K�����3J��T0 k� ������%�0d  e1�� Bb  ��D    �  ��I��Q��Q?� �V�|0P�c�D�
�W�����3J��T0 k� ������%�0d  e1�� Bb  ��D    �  ��I��R��Q?� ��U�|0P�[�D�
�[�����4J��T0 k� ������%�0d  e1�� Bb  ��D    �  ��I��S��Q?� ��Uݐ
|4P�W�D�
�c�����4J��T0 k� ������%�0d  e1�� Bb  ��D    �  ��I��S��Q?� ��Tݐ	|4P�O�E�
�g�����4EQ�T0 k� ������%�0d  e1�� Bb  ��D    �  ��I��T�Q?� �xT݌|8P�K�E�
�o������4EQ�T0 k� ������%�0d  e1�� Bb  ��D    �  ��I��U�Q?� �pS݈|8P�G�E�
�w������4EQ�T0 k� ������%�0d  e1�� Bb  ��D    �  ��I��U�Q?���hR݄|<P�?�E�
�{����� 4EQ�T0 k� ������%�0d  e1�� Bb �D    �  ��I��V ��Q?���`R��|<E�;�E�
Ѓ�����4EQ�T0 k� ������%�0d  e1�� Bb ��O    �  ��I��V ��Q?���XQ�||<E�7�E�
Ћ�����4EQ�T0 k� ������%�0d  e1�� Bb ��O    �  ��I��W �Q?���LO�t|@E�+�E�
З�����4Ea�T0 k� ������%�0d  e1�� Bb ��O    �  ��I��W �Q?���DN�t|@E�'�E�
П�����4Ea�T0 k� ������%�0d  e1�� Bb ��O    �  ��I��X �Q?���@M	p|@ E��E�|
������4Ea�T0 k� ������%�0d  e1�� Bb
 ��O    �  ��I��X �Q?���8L	l |@ E��D?t
��2��34Ea�T0 k� ����%�0d  e1�� Bb ��O    �  ��I��X �Q?��0K	k�|@ E��D?l
��2��33Ea�T0 k� ����%�0d  e1�� Bb ��O    �  ��I��Y@ۭQ?��,J	g�|@ E��D?h
��2��33C��T0 k� �'��+�%�0d  e1�� Bb ��O    �  ��I��Y@׮Q?��$I	g�|@ E��D?`
���2��33C��T0 k� �3��7�%�0d  e1�� Bb ��O    �  ��I��Y@ӮQ?�� H	c�|@ E��D?X
���2��33C��T0 k� �C��G�%�0d  e1�� Bb ��O    �  ��I��Y@˯Q?��G	_�|@ F�D?P
���2��32C��T0 k� �P �T %�0d  e1�� Bb ��O    �  ��I��Y@ǰQ?��F	[�|@ F��D?H
���2��3 2C��T0 k� �\ �` %�0d  e1�� Bb ��O    �  ��I��Y@ðQ?��D	[�|@ F��D?D
���2��3 1C��T0 k� �l�p%�0d  e1�� Bb ��O    �  ��I��Y@��Q?���C	W�|@ F��D?<
���2��3 1C� T0 k� �x�|%�0d  e1�� Bb ��O    �  ��I��Y@��Q?���B	S�|@ F��D?4
���2��3$0C� T0 k� ����%�0d  e1�� Bb ��O    �  ��I��Y@��Q?���A	O�|@ F�D?, 
��2��3$0C� T0 k� ����%�0d  e1�� Bb �O    �  ��I��Y@��Q?��� ?	O�|@ F�A�$!
������$0AR T0 k� ����%�0d  e1�� Bb �O    �  ��I��Y@��Q?����>	K�|@ F�A�"
������$/AR T0 k� ����%�0d  e1�� Bb ��O    �  ��A��Y@��Q?��=	G�|@ F�A�#
������$/AR T0 k� ����%�0d  e1�� Bb ��O    �  ��A��Y@��Q?��;	G�|@ E��A�$
�'�����(.AR T0 k� ����%�0d  e1�� Bb ��O   �  ��A��Y@��Q?��:	C�|@ E��A�%
�/�����(.AR T0 k� ����%�0d  e1�� Bb ��O    �  ��A��Y@��Q?��9	C�|@ E��A� &
�7�����(-AR T0 k� ����%�0d  e1�� Bb ��O    �  ��A��Y@��Q?{��7	?�|@ E��A��'
�?�����(-AR T0 k� ��	� 	%�0d  e1�� Bb ��O    �  ��BN�Y@�Q?{��6	;�|@ E�ߩA��'
�G�����(,AR T0 k� �
�
%�0d  e1�� Bb  ��O    �  ��BN�Y@{�Q?{��4	;�|@ E�ߪA��(
�O�����(,AR T0 k� ��%�0d  e1�� Bb! ��O    �  ��BN�Y0s�Q?w��3M7�|@ E�ߪA��)
�W�����,+AR T0 k� �(�,%�0d  e1�� Bb! ��O    �  ��BN�Y0o�Q?w���2M7�|@ E�߫A��*
�_�����,+ART0 k� �4�8%�0d  e1�� Bb" ��O    �  ��BN�Y0g�Q?w���0M3�|@ E�߬A��+
�g�����,+ART0 k� �D�H%�0d  e1�� Bb# ��O    �  ��B��Y0c�Q?w���/M/�|@ E�߬A��,
�k�����,*ART0 k� �P�T%�0d  e1�� Bb$ ��O    �  ��B��Y0[�Q?s���-M/�|@ B�߭A��-
�s�����,*ART0 k� �`�d%�0d  e1�� Bb% ��O    �  ��B��Y@W�Q?s���,M+�|@ B�߭A��.
�{�����,)ART0 k� �p�t%�0d  e1�� Bb% ��O    �  ��B��Y@O�Q?s���+M+�|@ B�߮A��.
у�����,)ART0 k� �|��%�0d  e1�� Bb& ��O    �  ��B��Y@K�QOs���*M'�|@ B�߯A��/
ч�����0)ART0 k� ����%�0d  e1�� Bb' ��O    �  ��B��Y@G�QOo���(M'�|@ B�߯A��0
я�����0(ART0 k� ����%�0d  e1�� Bb' ��O    �  ��B��Y@?�QOo���'M#�|@ B��A��1
ї�����0(ART0 k� ����%�0d  e1�� Bb( ��O    �  ��B��Y@;�QOo���&M#�|@ B��A��2
ћ�����0(ART0 k� ����%�0d  e1�� Bb( ��O    �  ��B��Y@7�QOo���%M�|@ B��A��2
ѣ�����0'ART0 k� ����%�0d  e1�� Bb) ��O    �  ��B��Y@/�QOo���#M�|@ E��A��3
ѫ�����0'ART0 k� ����%�0d  e1�� Bb* ��O    �  ��B��Y@+�QOk���"M�|@ E��A��4
ѯ�����0'ART0 k� ����%�0d  e1�� Bb* ��O    �  ��B��YP'�QOk���!M�|@ E��A��5
ѷ�����4&ART0 k� ����%�0d  e1�� Bb+ ��O    �  ��B��YP#�QOk��� M�|@ E��A��5
ѻ�����4&ART0 k� � �%�0d  e1�� Bb+ ��O    �  ��B��YP�Uk���M�|@ E��A��6
�������4&ART0 k� ��%�0d  e1�� Bb+ ��O    �  ��B��YP�Ug���M�|@ E��A��7
�������4%ART0 k� �� %�0d  e1�� Bb, ��O    �  ��B��YP�Ug���M�|@ E��A��7
�������4%ART0 k� �(�,%�0d  e1�� Bb, ��O    �  ��B��YP�Ug���M�|@ E���A��8
�������4%ART0 k� �8�<%�0d  e1�� Bb- ��O    �  ��B��YP�Ug���M�|@ E���A�|9
�������4$ART0 k� �H�L%�0d  e1�� Bb- ��O    �  ��B��YP�Ug���M�|@ E���A�t9
�������4$ART0 k� �T�X%�0d  e1�� Bb- ��O    �  ��B��Y_��Uc���M�|@ E���A�p:
�������4$ART0 k� �d�h%�0d  e1�� Bb- ��O    �  ��B��Y_��Uc���M�|@ E��A�l;
�������8#ART0 k� �p�t%�0d  e1�� Bb. ��O    �  ��B��Y_��Uc���M�|@ E��A�h;
�������8#ART0 k� ����%�0d  e1�� Bb. ��O    �  ��B� Yo��BOc�� M�|@ E��A�d<
�������8#ART0 k� � �� %�0d  e1�� Bb. ��O    �  ��B�Yo��BOc��M�|@ E��A�`<
�������8#ART0 k� � �� %�0d  e1�� Bb. ��O    �  ��B�Yo��BOc��M�|@ E��A�\=
�������8"ART0 k� �!��!%�0d  e1�� Bb. ��O    �  ��B�Yo��BOc��M�|@ E��A�X>
�������8"ART0 k� �"��"%�0d  e1�� Bb. ��O    �  ��B�Yo��BOc��M�|@ E��A�T>
�������8"ART0 k� ��#��#%�0d  e1�� Bb/ ��O    �  ��B�Yo��A�c��L��|@ E��A�P?
�������8"ART0 k� ��$��$%�0d  e1�� Bb/ ��O    �  ��B�Yo��A�_��L��|@ E��A�L?
�������8!ART0 k� ��$��$%�0d  e1�� Bb/ ��O    �  ��B�$Yo��A�_��L��|@ BM�A�H@
�������<!ART0 k� ��%��%%�0d  e1�� Bb/ ��O    �  ��B�(Yo��A�_��L��|@ BM�A�D@
�������<!ART0 k� � &�&%�0d  e1�� Bb/ ��O    �  ��B�0Yo��A�_�� L��|@ BM�A�@A
������<!ART0 k� �'�'%�0d  e1�� Bb/ ��O    �  ��B�4Yo��D�_��$L��|@ BM#�A�<A
������< ART0 k� � (�$(%�0d  e1�� Bb/ ��O    �  ��B�<Y��D�_��(L��|@ BM#�A�8B
������< ART0 k� �,(�0(%�0d  e1�� Bb. ��O    �  ��B�@Y��D�_�(L��|@ BM'�A�4C
������< ART0 k� �<)�@)%�0d  e1�� Bb. ��O    �  ��B�HY��D�_�,L��|@ BM'�A�0C
������< ART0 k� �H*�L*%�0d  e1�� Bb. ��O    �  ��B�LY�D�_�4L��|@ BM+�A�0C
������<AR T0 k� �X+�\+%�0d  e1�� Bb. ��O    �  ��B�TY�D�_�8L��|G�BM+�A�,D
������<AR T0 k� �h,�l,%�0d  e1�� Bb. ��O    �  ��IXY�D�_�<L��|G�BM/�A�(D
������<AR T0 k� �t,�x,%�0d  e1�� Bb. ��O    �  ��I`Y�D�_�@L��|G�BM/�A�$E
������<AR T0 k� �-��-%�0d  e1�� Bb- ��O    �  ��IdY�	D�[�DL��|G�BM3�A� E
������@AR$T0 k� �.��.%�0d  e1�� Bb- ��O    �  ��IhY�D�X HL��|G�BM3�A�F
�#�����@AR$T0 k� �/��/%�0d  e1�� Bb- ��O    �  ��IlY�D�XPL��|G�BM7�A�F
�#�����@AR$	T0 k� �0��0%�0d  e1�� Bb, ��O    �  ��I/pY�D�XTL��|G�BM7�A�G
�'�����@AR$	T0 k� �0��0%�0d  e1�� Bb, ��O    �  ��I/tYO�D�XXL��|G�BM;�A�G
�+�����@AR(	T0 k� ��1��1%�0d  e1�� Bb, ��O    �  ��I/xYO�D�X`L��|G�BM;�A�H
�+�����@AR(	T0 k� ��2��2%�0d  e1�� Bb+ ��O    �  ��I/|YO�D�X�dL��|G�BM?�A�H
�/�����@AR(	T0 k� ��3��3%�0d  e1�� Bb+ ��O    �  ��I/�YO�D�X�lL��|G�BM?�A�H
�/�����@AR(
T0 k� ��4��4%�0d  e1�� Bb* ��O    �  ��K��YO�D�X�pL��|G�BMC�A�I
�3�����@AR,
T0 k� �4�4%�0d  e1�� Bb* ��O    �  ��K��YO�D�X�xL��|G�BMC�A�I
�7�����@AR,
T0 k� �5�5%�0d  e1�� Bb) ��O    �  ��K��YO�D�X�|L��|G�BMG�A�J
�7�����@AR,
T0 k� � 6�$6%�0d  e1�� Bb) ��O    �  ��K��YO�!D�X	��L��|K�BMG�A� J
�;�����@AR,
T0 k� �07�47%�0d  e1�� Bb( ��O    �  ��K��YO�#D�X
��L��|K�BMK�A� J
�;�����@AR,
T0 k� �<8�@8%�0d  e1�� Bb( ��O    �  ��K��YO�%D�X��L��|K�BMK�A��K
�?�����DAR0T0 k� �L8�P8%�0d  e1�� Bb' ��O    �  ��K��YO�'D�X��L��|K�BMK�A��K
�C�����DAR0T0 k� �\9�`9%�0d  e1�� Bb& ��O    �  ��K��YO�)D�T��L��|K�BMO�A��L
�C�����DAR0T0 k� �h:�l:%�0d  e1�� Bb& ��O    �  ��K��Y_�+D�T��L��|K�BMO�A��L
�G�����DAR0T0 k� �x;�|;%�0d  e1�� Bb% ��O    �  ��K��Y_�-D�T��L��|K�BMS�A��L
�G�����DAR0T0 k� �<��<%�0d  e1�� Bb$ ��O    �  ��K��Y_�/D�T��L��|K�BMS�A��M
�K�����DAR4T0 k� �<��<%�0d  e1�� Bb# ��O    �  ��K��Y_|2D�T��L��|K�BMS�A��M
�K�����DAR4T0 k� �=��=%�0d  e1�� Bb# ��O   �  ��K��Y_x4D�T��L��|K�BMW�A��M
�O�����DAR4T0 k� �>��>%�0d  e1�� Bb" ��O    �  ��K��Y�x6D�T��L��|K�BMW�A��N
�O�����DAR4T0 k� ��?��?%�0d  e1�� Bb! ��O    �  ��K��Y�t8D�T��L��|K�BM[�A��N
�S�����DAR4T0 k� ��@��@%�0d  e1�� Bb  ��O    �  ��K��Y�t:D�T��L��|K�BM[�A��N
�S�����DAR4T0 k� ��@��@%�0d  e1�� Bb ��O    �  ��K��Y�p<D�T��L��|K�BM[�A��O
�W�����DAR8T0 k� ��A��A%�0d  e1�� Bb ��O    �  ��K��Y�p=D�T��L��|K�BM_�A��O
�W�����DAR8T0 k� ��B��B%�0d  e1�� Bb ��O    �  ��K��Y�l?D�T��L��|K�BM_�A��O
�[�����DAR8T0 k� �C�C%�0d  e1�� Bb ��O    �  ��K��Y�lAD�T��L��|K�BM_�A��P
�[�����DAR8T0 k� �D�D%�0d  e1�� Bb ��O    �  ��K��Y�hCD�T!�L��|K�BMc�A��P
�_�����HAR8T0 k� �$D�(D%�0d  e1�� Bb ��O    �  ��K��Y�hED�T#�L��|O�BMc�A��P
�_�����HAR8T0 k� �4E�8E%�0d  e1�� Bb ��O    �  ��K��Y�dGD�T$�L��|O�BMc�A��P
�_�����HAR<T0 k� �@F�DF%�0d  e1�� Bb ��O    �  ��K��Y�dHD�T&�L��|O�BMg�A��Q
�c�����HAR<T0 k� �PG�TG%�0d  e1�� Bb ��O    �  ��K��Y�`JD�T(�$L��|O�BMg�A��Q
�c�����HAR<T0 k� �\H�`H%�0d  e1�� Bb ��O    �  ��K��Y�`LD�T*�,L��|O�BMg�A��Q
�g�����HAR<T0 k� �lH�pH%�0d  e1�� Bb ��O    �  ��K��Y�\MD�T,�4L��|O�BMk�A��R
�g�����HAR<T0 k� �|I��I%�0d  e1�� Bb ��O    �  ��K��Y�\OD�T-�<L��|O�BMk�A��R
�k�����HAR<T0 k� �J��J%�0d  e1�� Bb ��O    �  ��K��Y�XQD�P/�DL��|O�BMk�A��R
�k�����HAR@T0 k� �K��K%�0d  e1�� Bb ��O    �  ��K��Y�XRD�P1�LL��|O�BMk�A��R
�k�����HAR@T0 k� �L��L%�0d  e1�� Bb ��O   �  ��K��Y�TTD�P3�TL��|O�BMo�A��S
�o�����HAR@T0 k� �L��L%�0d  e1�� Bb ��O    �  ��K��Y�TUD�P5�\|��|O�BMo�A��S
�o�����HAR@T0 k� ��M��M%�0d  e1�� Bb ��O    �  ��K��Y�TWD�P7�d|��|O�BMo�A��S
�o�����HAR@T0 k� ��N��N%�0d  e1�� Bb ��O    �  ��K��Y�PXD�P9�l|��|O�BMs�A��S
�s�����HAR@T0 k� ��O��O%�0d  e1�� Bb ��O    �  ��K��Y�PZFP;�t|��|O�BMs�A��T
�s�����HAR@T0 k� ��P��P%�0d  e1�� Bb	 ��O    �  ��K��Y�L[FP=�||��|O�BMs�A��T
�w�����HAR@T0 k� ��Q� Q%�0d  e1�� Bb ��O    �  ��K��Y�L]FP?��|��|O�BMs�A��T
�w�����HARDT0 k� �Q�Q%�0d  e1�� Bb ��O    �  ��K��Y�L^FTA��|��|O�BMw�A��T
�w�����HARDT0 k� �R�R%�0d  e1�� Bb ��O    �  ��K��Y�H_FTC��|��|O�BMw�A��U
�{�����HARDT0 k� �(S�,S%�0d  e1�� Bb ��O   �  ��K��Y�HaFTE��|��!�O�BMw�A��U
�{�����HARDT0 k� �4T�8T%�0d  e1�� Bb ��O    �  ��K��Y�DbFTG��|��!�O�BMw�A��U
�{�����LARDT0 k� �DU�HU%�0d  e1�� Bb  ��O    �  ��K��Y�DcFTI�����!�O�BM{�A��U
������LARDT0 k� �TU�XU%�0d  e1�� Bb  ,�O    �  ��K��Y�DeFXK�����!�O�BM{�A��U
������LARDT0 k� �`V�dV%�0d  e1�� Bb  ��O    �  ��K� Y�@fFXM�����!�S�BM{�A��V
������LARDT0 k� �pW�tW%�0d  e1�� Bb ��O   �  ��K� Y�@gFXO�����!�S�BM{�A��V
҃�����LARHT0 k� �|X��X%�0d  e1�� Bb ��O    �  ��K�Y�@iE�\R�����!�S�BM�A��V
҃�����LARHT0 k� �Y��Y%�0d  e1�� Bb (�O    �  ��K�Y�<jE�\T�����!�S�BM�A��V
҃�����LARHT0 k� $�X��X%�0d  e1�� Bb ��O    �  ��K�Y�<kE�`U�����!�S�BM�A��V
҃�����LARHT0 k� $�W��W%�0d  e1�� Bb ��O    �  ��K�Y�<lE�`W�����!�S�BM�A��W
҇�����LARHT0 k� $�V��V%�0d  e1�� Bb ��O    �  ��K�Y�8mE�dY�����!�S�BM��A��W
҇�����LARHT0 k� $�V��V%�0d  e1�� Bb ��O    �  ��K�Y�8nE�d[��|��|S�BM��A��W
҇�����LARHT0 k� $|U��U%�0d  e1�� Bb ��O   �  ��K�Y�8pE�h]��|��|S�BM��A��W
ҋ�����LARHT0 k� $|T��T%�0d  e1�� Bb ��O    �  ��K�Y�8qE�l_��|��|S�BM��A��W
ҋ�����LARHT0 k� �xS�|S%�0d  e1�� Bb  ��O    �  ��K�Y�4rE�pa��|��|S�BM��A��X
ҋ�����LARLT0 k� �tS�xS%�0d  e1�� Bb  ��O    �  ��K�Y�4sE�pb��|��|S�BM��A��X
ҋ�����LARLT0 k� �pR�tR%�0d  e1�� Bb  .�O    �  ��K�Y�4tE�td� |��|S�BM��A��X
ҏ�����LARLT0 k� �pQ�tQ%�0d  e1�� Bb  ��O    �  ��K�Y�0uE�xf�|��|S�BM��A��X
ҏ�����LARLT0 k� �lQ�pQ%�0d  e1�� Bb  ��O    �  ��K�Y�0vE�|g�|��|S�BM��A��X
ҏ�����LARLT0 k� 4hP�lP%�0d  e1�� Bb  ��O    �  ��K�Y�0wE��i�|��|S�BM��A��X
ҏ�����LARLT0 k� 4dO�hO%�0d  e1�� Bb  ��O    �  ��K�Y�0xE��j�L��|S�BM��A��Y
ғ�����LARLT0 k� 4dN�hN%�0d  e1�� Bb  ��O    �  ��K�Y�,yE��l�L��|S�BM��A��Y
ғ�����LARLT0 k� 4`N�dN%�0d  e1�� Bb  ��O    �  ��K�Y�,zE��m�$L��!�S�BM��A��Y
ғ�����LARLT0 k� 4\M�`M%�0d  e1�� Bb  ��O    �  ��K� Y�,{E��n�(L��!�S�BM��A��Y
ғ�����LARLT0 k� �\L�`L%�0d  e1�� Bb  ��O    �  ��K� Y�(|E��p�,L��!�S�BM��A��Y
җ�����LARLT0 k� �XL�\L%�0d  e1�� Bb  ��O    �  ��K� Y�(}E��q�0|��!�S�BM��A��Y
җ�����LARPT0 k� �TK�XK%�0d  e1�� Bb  ��O   �  ��K� Y�(~E��r�8|��!�S�BM��A��Z
җ�����LARPT0 k� �PJ�TJ%�0d  e1�� Bb  ��O    �  ��K� Y�(~E��s�<|��!�S�BM��A��Z
җ�����PARPT0 k� �PJ�TJ%�0d  e1�� Bb  ��O    �  ��K� Y�$E��t�@|��!�S�BM��A��Z
қ�����PARPT0 k� �LI�PI%�0d  e1�� Bb  ��O    �  ��@` Y�$�E��u�D|��!�S�BM��A��Z
қ�����PARPT0 k� �HH�LH%�0d  e1�� Bb  ��O    �  ��@` Y�$�E��u�H|��!�S�BM��A��Z
қ�����PARPT0 k� �HG�LG%�0d  e1�� Bb  ��O    �  ��@` Y�$�E��v�P|��!�S�BM��A��Z
қ�����PARPT0 k� �DG�HG%�0d  e1�� Bb  ��O    �  ��@` Y�$E��w�T|��!�S�BM��A��Z
қ�����PARPT0 k� �@F�DF%�0d  e1�� Bb  ��O    �  ��@` YO E��w�X|��|S�BM��A��[
ҟ�����PARPT0 k� �@E�DE%�0d  e1�� Bb  ��O    �  ��@` YO E��x�\���|S�BM��A��[
ҟ�����PARPT0 k� �<E�@E%�0d  e1�� Bb  ��O    �  ��@� YO E��y�`���|W�BM��A��[
ҟ�����PARPT0 k� �8D�<D%�0d  e1�� Bb  ��O    �  ��@� YO E��y�d���|W�BM��A��[
ҟ�����PARPT0 k� �4C�8C%�0d  e1�� Bb  ��O    �  ��@� YO ~E��y�h���|W�BM��A��[
ҟ�����PARPT0 k� �4C�8C%�0d  e1�� Bb  ��O    �  ��@� Y �~E��z�l���|W�BM��A��[
ң�����PARTT0 k� �0B�4B%�0d  e1�� Bb  ��O    �  ��@� Y �~E��z�p���|W�BM��A��[
ң�����PARTT0 k� �,A�0A%�0d  e1�� Bb  ��O    �  ��A  Y �~E��z�t���|W�BM��A��[
ң�����PARTT0 k� �,A�0A%�0d  e1�� Bb  ��O    �  ��A  Y �}E��z�x���|W�BM��A��\
ң�����PARTT0 k� �(@�,@%�0d  e1�� Bb  ��O    �  ��A  Y �}E��z�|���|W�BM��A��\
ң�����PARTT0 k� �$?�(?%�0d  e1�� Bb  ��O    �  ��A  Y o}E��{΀|��|W�BM��A��\
ҧ�����PARTT0 k� �$?�(?%�0d  e1�� Bb  ��O    �  ��A  Y o}E��{΄|��|W�BM��A��\
ҧ�����PARTT0 k� � >�$>%�0d  e1�� Bb  ��O    �  ��AP Y o}C��{Έ|��|W�BM��A��\
ҧ�����PARTT0 k� �=� =%�0d  e1�� Bb  ��O    �  ��AP Y o |C��{ΐ|��|W�BM��A��\
ҧ�����PARTT0 k� �<�<%�0d  e1�� Bb  ��O    �  ��AP Y |C��{ΐ|��|W�BM��A��\
ҧ�����PARTT0 k� �;�;%�0d  e1�� Bb  ��O    �  ��APY |C��zΔ|��|W�BM��A��\
ҫ�����PARTT0 k� �;�;%�0d  e1�� Bb  ��O    �  ��C�Y${C��zΘ|��|W�BM��A��]
ҫ�����PARTT0 k� �:�:%�0d  e1�� Bb  ��O    �  ��C�Y${K��z��|��|W�BM��A��]
ҫ�����PARTT0 k� �9�9%�0d  e1�� Bb  ��O    �  ��C�Y({K��z��L��|W�BM��A��]
ҫ�����PARTT0 k� �9�9%�0d  e1�� Bb  ��O    �  ��C�Y�(zK��z�� L��|W�BM��A��]
ҫ�����PARXT0 k� �8�8%�0d  e1�� Bb  ��O    �  ��C�Y�,zK��z�� L��|W�BM��A��]
ҫ�����PARXT0 k� �7�7%�0d  e1�� Bb  ��O    �  ��C�Y�,yK��y�� L��|W�BM��A��]
ҫ�����PARXT0 k� � 7�7%�0d  e1�� Bb  ��O    �  ��C�Y�0yK��y�� L��|W�BM��A��]
ү�����PARXT0 k� � 6�6%�0d  e1�� Bb  ��O    �  ��C�Y�4xK��y�� L��|W�BM��A��]
ү�����PARXT0 k� ��5� 5%�0d  e1�� Bb  ��O   �  ��C�Y�4xK��y�� L��|W�BM��A�|]
ү�����PARXT0 k� ��5� 5%�0d  e1�� Bb  ��O    �  ��C�Y�8wK��y��!L��|W�BM��A�|^
ү�����PARXT0 k� ��4��4%�0d  e1�� Bb  ��O    �  ��C�Y�<wK��y��!L��|W�BM��A�|^
ү�����PARXT0 k� ��3��3%�0d  e1�� Bb  ��O    �  ��C�Y�@vK��y��!L��|W�BM��A�|^
ү�����PARXT0 k� ��3��3%�0d  e1�� Bb  ��O    �  ��C� Y�DuK��x��!L��|W�BM��A�|^
ү�����PARXT0 k� ��2��2%�0d  e1�� Bb  ��O    �  ��C��Y�DuK��x��"L��|W�BM��A�|^
ҳ�����PARXT0 k� ��1��1%�0d  e1�� Bb  ��O    �  ��K�Y�HtK��x��"L��|W�BM��A�|^
ҳ�����TARXT0 k� ��1��1%�0d  e1�� Bb  ��O    �  ��K�Y�LsL�x��#L��|W�BM��A�x^
ҳ�����TARXT0 k� ��0��0%�0d  e1�� Bb  ��O    �  ��K�Y�PrL�x��#L��|W�BM��A�x^
ҳ�����TARXT0 k� ��/��/%�0d  e1�� Bb  ��O    �  ��K�Y�TrL�x��$L��|W�BM��A�x^
ҳ�����TARXT0 k� ��/��/%�0d  e1�� Bb  ��O    �  ��K�Y�XqL�x��$L��|W�BM��A�x^
ҳ�����TARXT0 k� ��.��.%�0d  e1�� Bb  ��O    �  ��Eo�X�\pL�x�%L��|W�BM��A�x^
ҳ�����TARXT0 k� ��.��.%�0d  e1�� Bb  ��O    �  ��Eo�X�`oL�w�%L��|W�BM��A�x^
ҳ�����TARXT0 k� ��-��-%�0d  e1�� Bb  ��O    �  ��Eo�X�dnL�w�&L��|W�BM��A�x_
ҷ�����TARXT0 k� ��,��,%�0d  e1�� Bb  ��O    �  ��Eo�X�hmL  w�'L��|W�BM��A�x_
ҷ�����TARXT0 k� ��,��,%�0d  e1�� Bb  ��O    �  ��Eo�W�lmL  w�'L��|W�BM��A�t_
ҷ�����TAR\T0 k� ��+��+%�0d  e1�� Bb  ��O    �  ��E�W�llL  w�(L��|W�BM��A�t_
ҷ�����TAR\T0 k� ��*��*%�0d  e1�� Bb  ��O    �  ��E�V�plL  w�)L��|W�BM��A�t_
ҷ�����TAR\T0 k� ��*��*%�0d  e1�� Bb  ��O    �  ��E�V�tkL  w *L��|W�BM��A�t_
ҷ�����TAR\T0 k� ��)��)%�0d  e1�� Bb  ��O    �  ��E�U�tkL w+L��|W�BM��A�t_
ҷ�����TAR\T0 k� ��(��(%�0d  e1�� Bb  ��O    �  ��E�U�xjL w+L��|W�BM��A�t_
ҷ�����TAR\T0 k� ��(��(%�0d  e1�� Bb  ��O    �  ��L_�T�|jL v,L��|W�BM��A�t_
ҷ�����TAR\T0 k� ��'��'%�0d  e1�� Bb  ��O    �  ��L_�T�|iL v-L��|[�BM��A�t_
һ�����TAR\T0 k� ��'��'%�0d  e1�� Bb  ��O    �  ��L_�T�|iL v.L��|[�BM��A�t_
һ�����TAR\T0 k� ��&��&%�0d  e1�� Bb  ��O    �  ��L_�S��iL v /L��|[�BM��A�t_
һ�����TAR\T0 k� ��%��%%�0d  e1�� Bb  ��O    �  ��L_�S��iL v(0L��|[�BM��A�p_
һ�����TAR\T0 k� ��%��%%�0d  e1�� Bb  ��O    �  ��L_�R��hL v,1L��|[�BM��A�p_
һ�����TAR\T0 k� ��$��$%�0d  e1�� Bb  ��O    �  ��L_�R��hL v�42L��|[�BM��A�p`
һ�����TAR\T0 k� ��#��#%�0d  e1�� Bb  ��O    �  ��L_�Q��hL v�83L��|[�BM��A�p`
һ�����TAR\T0 k� ��#��#%�0d  e1�� Bb  ��O    �  ��L_�Q��hL v�<4L��|[�BM��A�p`
һ�����TAR\T0 k� ��"��"%�0d  e1�� Bb  ��O    �  ��L_�Q��hL v�D5L��|[�BM��A�p`
һ�����TAR\T0 k� ��"��"%�0d  e1�� Bb  ��O    �  ��L_�P��hL v�H6L��|[�BM��A�p`
һ�����TAR\T0 k� ��!��!%�0d  e1�� Bb  ��O    �  ��Lo�P��hL u�P8L��|[�BM��A�p`
ҿ�����TAR\T0 k� �� �� %�0d  e1�� Bb  ��O    �  ��Lo�P��hL u�X9L��|[�BM��A�p`
ҿ�����TAR\T0 k� �� �� %�0d  e1�� Bb  ��O   �  ��Lo�O�hL u�\:L��|[�BM��A�p`
ҿ�����TAR\T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�O�hL u�`;L��|[�BM��A�p`
ҿ�����TAR\T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�N�hL u�h<L��|[�BM��A�l`
ҿ�����TAR\T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�N�hL u�l>L��|[�BM��A�l`
ҿ�����TAR\T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�N�hL u	_t?L��|[�BM��A�l`
ҿ�����TAR\T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�M�hL u	_x@L��|[�BM��A�l`
ҿ�����TAR\T0 k� ����%�0d  e1�� Bb  ��O   �  ��Lo�M�hL u	_|AL��|[�BM��A�l`
ҿ�����TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�M�hL u	_�BL��|[�BM��A�l`
ҿ�����TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�L�hL u	_�BL��|[�BM��A�l`
ҿ�����TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�M�hL u	o�CL��|[�BM��A�l`
ҿ�����TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�M�hL u	o�CL��|[�BM��A�la
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�M�hL t	o�CL��|[�BM��A�la
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�M�hL t	o�CL��|[�BM��A�la
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�N�hL t	o�CL��|[�BM��A�la
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O   �  ��Lo�N�hK�tO�CL��|[�BM��A�la
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�N�hK�tO�DL��|[�BM��A�ha
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�N�hK�tO�DL��|[�BM��A�ha
�������TAR`T0 k� �|��%�0d  e1�� Bb  ��O    �  ��Lo�N�hK�tO�DL��|[�BM��A�ha
�������TAR`T0 k� �x�|%�0d  e1�� Bb  ��O    �  ��Lo�O�hK�tO�EL��|[�BM��A�ha
�������TAR`T0 k� �x�|%�0d  e1�� Bb  ��O    �  ��Lo�O��hK�tO�EL��|[�BM��A�ha
�������TAR`T0 k� �t�x%�0d  e1�� Bb  ��O    �  ��Lo�O��hC�tO�EL��|[�BM��A�ha
�������TAR`T0 k� �t�x%�0d  e1�� Bb  $�O   �  ��Lo�O��hC�tO�FL��|[�BM��A�ha
�������TAR`T0 k� 3t�x%�0d  e1�� Bb  ��O    �  ��Lo�O��hC�tO�FL��|[�BM��A�ha
�������TAR`T0 k� 3x�|%�0d  e1�� Bb  ��O    �  ��Lo�P��hC�sO�GL��|[�BM��A�ha
�������TAR`T0 k� 3x�|%�0d  e1�� Bb  ��O    �  ��Lo�P��hC�sO�HL��|[�BM��A�ha
�������TAR`T0 k� 3|��%�0d  e1�� Bb  ��O    �  ��Lo�P��hC�sO�HL��|[�BM��A�ha
�������TAR`T0 k� 3|��%�0d  e1�� Bb  ��O    �  ��Lo�P��hC�s_�IL��|[�BM��A�ha
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�P��hC�r_�JL��|[�BM��A�ha
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�Q��hC�r_�JL��|[�BM��A�ha
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�Q��hC�q_�KL��|[�BM��A�ha
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�Q��hC�q_�KL��|[�BM��A�ha
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�Q��hC�q_�LL��|[�BM��A�ha
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�Q��hC�p_�LL��|[�BM��A�hb
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�Q��hC�p_�LL��|[�BM��A�db
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�R��hC�o_�ML��|[�BM��A�db
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�R��hC�n_�ML��|[�BM��A�db
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�R��hC�n_�ML��|[�BM��A�db
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�R��hE�mo�ML��|[�BM��A�db
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��Lo�R��hE�lo�ML��|[�BM��A�db
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��L_�R��hE�lo�ML��|[�BM��A�db
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��L_�R��hE�ko�ML��|[�BM��A�db
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��L_�S��hE� jo�ML��|[�BM��A�db
�������TAR`T0 k� ����%�0d  e1�� Bb  ��O    �  ��L_�S��hE��j ��ML��|[�BM��A�db
�������TARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��L_�S��hE��i ��ML��|[�BM��A�db
�������TARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��L_�S��hE��h ��ML��|[�BM��A�db
�������TARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��K?�S��hE��g ��ML��|[�BM��A�db
�������TARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��K?�S��hE��g ��ML��|[�BM��A�db
�������TARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��K?�S��hEo�f ��ML��|[�BM��A�db
�������TARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��K?�S��hEo�e ��ML��|[�BM��A�db
�������TARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��K?�S��hEo�d ��ML��|[�BM��A�db
�������TARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��Ko�S��hEo�cO�ML��|[�BM��A�db
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��Ko�S��hEo�cO�NL��|[�BM��A�db
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��Ko�S��hE�cO�NL��|[�BM��A�db
�������XARdT0 k� ����%�0d  e1�� Bb  ��O   �  ��Ko�R��hE�bO�NL��|[�BM��A�db
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��Ko�R��hE�bO�NL��|[�BM��A�db
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��J�Q��hE�aO�OL��|[�BM��A�db
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��J�Q��hE�aO�OL��|[�BM��A�db
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��J�P��hE��`O�OL��|[�BM��A�db
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��J�P��hE��_O�PL��|[�BM��A�db
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��J�O��hE��_O�P|��|[�BM��A�db
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��J�O�hE��_O�Q|��|[�BM��A�`b
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��J�N�hE��^O�R|��|[�BM��A�`b
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��J�N�hE��]_�R|��|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E��M�hE�]_�S|��|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E��M�hE�\_�S|��|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E��M�hE�\_�T|��|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E��LO�hE�\_�T|��|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E��LO�hE�[߈U|��|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E��KO�hJ�[߈U|��|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E�KO�hJ�[߈V���|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E�KO�hJ�Z߈V���|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E�J��gJ�Z߈W���|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E�J��gJ�Z߈W���|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��E�J��gJ�Z߈W���|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��D��J��gJ�Z߈W���|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��D��J��gJ�Z߈W���|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��D��J��gJ/�Z߈W���|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��D��J��gJ/�Z߈W���|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��D��J��gJ/�Z߈W|��|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��D��J��gJ/�Z�W|��|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O   �  ��D��J��gJ/�Z�W|��|[�BM��A�`c
�������XARdT0 k� ����%�0d  e1�� Bb  ��O    �  ��C�d �K�(g$\O�W|(@�@� � ���;�Z3�T0 k� �C�#İ %�0d  e1�� B ��    �  C�d �K�(g$\O�W|(@�@� � ���;�Z3�T0 k� �C�#İ %�0d  e1�� B ��    �  C�d �K�(g$\N�W|(@�@� � ���;�Z3�T0 k� �C�#İ %�0d  e1�� B ��    �  C�d �K�(g$`N�W|(@�@� � ���;�Z3�T0 k� �C�#İ %�0d  e1�� B ��    �  @c�d �K�(g$`N�W|(@�@� � ���;�Z3�T0 k� �C�#İ %�0d  e1�� B ��    �  @c�d �K�(g$`N�W|(@�@� � ���;�Z3�T0 k� �C�#� %�0d  e1�� B ��    �  @c�d �K�(g$`N�W|(@�@� � ���;�Z3�T0 k� �C�#� %�0d  e1�� B ��    �  @c�d �K�(g$dM�W|(@�@� � ���;�Z3�T0 k� �C�#� %�0d  e1�� B ��    �  @c�d �K�(g$dM�W|(@�@� � ���;�Z3�T0 k� �C�#� %�0d  e1�� B ��    �  @��d �K�(gdM� W|(@�@� � ���;�Z3�T0 k� �C�#� %�0d  e1�� B ��    �  @��d �K�(ghM� W|(@�@�� � ���;�Z3�T0 k� �C�#�� %�0d  e1�� B ��    �  @��d �K�(ghM�$W|(@�@| � ���;�Z3�T0 k� �C�#�� %�0d  e1�� B ��    �  @��d �K�(ghM�$W|(@�@| � ���;�Z3�T0 k� �C�#�� %�0d  e1�� B ��    �  @��d �K�(ghL�$W|(@�@| � ���;�Z3�T0 k� �C�#�� %�0d  e1�� B ��    �  @��d �K�(hlL�$W|(@�@| � ���;�Z3�T0 k� �C�#�� %�0d  e1�� B ��    �  @��d �K�(hlL�(W|(@�@|~ � ���;�Z3�T0 k� �C�$� %�0d  e1�� B ��    �  @��d �K�(hlL�(W|(@�@|~ � ���;�Z3�T0 k� �C�$� %�0d  e1�� B ��    �  @��d �K�(hlL�,W|(@�@|~ � ���;�Z3�T0 k� �C�$� %�0d  e1�� B ��    �  @��d �K�(hlL�0W|(@�@|~ � ���;�Z3�T0 k� �C�$� %�0d  e1�� B ��    �  @��d �K�(ilL�0W|(@�@|} � ���;�Z3�T0 k� �C�$� %�0d  e1�� B ��    �  @��d �K�(ilL�4X|(@�@|} � ���;�Z3�T0 k� �C�#4� %�0d  e1�� B ��    �  @��d �K�(ilL�4X|(@�@|} � ���;�Z3�T0 k� �C�#4� %�0d  e1�� B ��    �  @��d �K�(ilL�8Y|(@�@x} � ���;�Z3�T0 k� �C�#4� %�0d  e1�� B ��    �  K��d �K�(jlL�8Y|(@�@x| � ���;�Z3�T0 k� �C�#4� %�0d  e1�� B ��    �  K��d �K�(jlL�<Z|(@�@x| � ���;�Z3�T0 k� �C�#4� %�0d  e1�� B ��    �  K��d �K�(j�lM�<Z|(@�@x| � ���;�Z3�T0 k� �C�#T� %�0d  e1�� B ��    �  K��d �K�(j�lM�<Z|(@�@x| � ���;�Z3�T0 k� �C�#T� %�0d  e1�� B ��    �  K��d �K�(k�hM�@Z|(@�@x| � ���;�Z3�T0 k� �C�#T� %�0d  e1�� B ��    �  K��d �K�(k�hM�@[|(@�@x{ � ���;�Z3�T0 k� �C�#T� %�0d  e1�� B ��    �  K��d �K�(k�hN�@[|(@�@x{ � ���;�Z3�T0 k� �C�#T� %�0d  e1�� B ��    �  K��d �K�(l�hN�@\|(@�@x{ � ���;�Z3�T0 k� �C�#d� %�0d  e1�� B ��    �  K��d �K�(l�hN�@\|(@�@x{ � ���;�Z3�T0 k� �C�#d� %�0d  e1�� B ��    �  K��d �K�(l�hN�@]|(@�@x{ � ���;�Z3�T0 k� �C�#d� %�0d  e1�� B ��    �  K��d �K�$m�dN�@]|(@�@x{ � ���;�Z3�T0 k� �C�#d� %�0d  e1�� B ��    �  K��d �K�$m�dN�@^|(@�@xz � ���;�Z3�T0 k� �C�#d� %�0d  e1�� B ��    �  K��d �K�$m�dO�<^|(@�@xz � ���;�Z3�T0 k� �C�#t� %�0d  e1�� B ��    �  @��2 ���P� O8# o;�!� A�+�@�(2P<  ����#AP� T0 k� �  � %�0d  e1�� Bb  ��/    �   2@��2 ���P� O8# o;�!� A�+�@�(2P<  ����#AP� T0 k� �  � %�0d  e1�� Bb  /�/    �   /@��2 ���P� O8# o;�!� A�+�@�(2P<  ����#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �   +@��2 ���@o� O8# o;�!� A�+�@�(2 <  ����#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �   'CO�2 ���@o� O8#�;�!� A�+�@�(2 <  ����#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �   #CO�2 ���@o� O8#�;�| A�+�@�(2 <  ����#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �    CO�1 ���@o� O8#�;�|  A�+�@�(2 <  ����#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �   CO�1 ���@o� O8#�;�|  A�+�@�(2 <  ����#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �   CO�1��@�� O8#�;�|$ @+�@�(2p< @��P�#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �   CO�1��@��  8#�?�|$ @+�@�(2p< @��P�#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �   CO�0��@��  8#�?�|$ @+�A (1p< @��P�#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �   CO�0��@��  8#�?�|( @+�A (1p< @��P�#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �   CO�/��@��  8#�C�|( @+�A (1p< @��P�#AP� T0 k� �� �� %�0d  e1�� Bb  ��/    �                                                                                                                                                                               � � �  �  �  c A�  �J����   �      6 \���0 ]�(!(  � � Jis  H H	     ���k     JCD��^�    ��            ? Z��          @�     ���   0	%           g<          �����     g<����                   	 Z��          �     ���   0	           ZP�  � �      ���C     ZP���1      ��             *	 Z��          �@
�    ���   8	           W5R   � �	   ��W�     W9_��\j    ����              		 Z��           �  &  ���  8         �ϡO   � �      .�*�    �ϡ��*�K    ����             P  Z��          �p�    ���  P
	
         ���  ��	      B���    ������                             ���               (  ���    P             ��N $ $      V�m�]    �� �m��     n d              
     9         ��     ��B   8

            c~�   	    j�X��     cxq�X��     \��                8         �     ��@   (
 
          ��ss  � �	     ~ �i&    ��ss �a?       w         
     4�        0
`     ��P   8�         ��x3   �
	   � ���    ��x3 ���                     �� d         	 �     ��@   P


	          xg   �	      � ��     xg ��                        d         
 �     ��@   P
B          ��  �	     � ��Z     � ���     ' 4                 ����O         �     ��H   H
	 
                ��      �                                                                           �                               ��        ���          ��                                                                 �                          �  ��        � �ǈ     � �J�      Y                   x                j  �   �   �                              ��        � �          �           "                                                �                         ���������*��m�X � � � ��� � �          
  	     
  3   � �  ���I       �d 0c@ �� 0c� �$ d  �D  d  ��  d` �  d� �D d����X � �� b� E�  a� �d s� �� s� .� `m@ /� n  /�  n  /� n` 
� W� �� �w@ �� x@ 
�< V� 
�� V� 
�\ W  
� W� 
�< W� 
�\ W� �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }` 
�\ W� 
� W� 
�� W����� � 
� W����� � 
�| W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������  ��   ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    B�j l �  B �
� �  �  
�  ��  ��     ��a  �   ����  ��     ��*           ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �O       �� �T ��        � �  ��        �        ��        �        ��        �     ��	       2��        ��                         �w� $  ������                                     �                D��� 	          
  ����%��    �� 2                3 Zarley Zalapski     1:19                                                                        4  4     �C
2� � �
�	ckjX{ krhKkV �[ k^ � �B�^ � B�V �	CP �
CX � C Q �C!P �C#[ �J�D � J�T �J�< �KP � K` �KP � K` � KS � KT �  Kt �  Kh �  KX �  Kr{ *� �b"� �b*� ��"� �� "� �y � �y 
� �r 
� �?#� �? 
� �5%"� �5 &"� �%'� �% 
� �)� � 
� � 
� �',"� �' -"� �.� � 
� �0� � 
� �2� � 
� � 
� � 
� � �6" � � 7!� � �8"" � �9!� � �:!� � �;" �<*$7 �=* O �  *O � * O                                                                                                                                                                                                                         H� R         �    ` 
        �     \ P E ]  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��    ��@�� ��������������������������������������������������������   �4, *� 6 A� ͂�@� @���@���Z����� �����%�                                                                                                                                                                                                                                                                                                                   @@Ҙ                                                                                                                                                                                                                                             A  
  )     �  D�J    	  H                             ������������������������������������������������������                                                                                                                                      �      �      �                �  �          	  
 	 
 	 	 ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ���           )                  (    $    ��  L�J ��   �                             ������������������������������������������������������                                                                     
                                                                �   ��,     1      �        OGM )          	     	 	 ���������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������           x                                                                                                                                                                                                                                     
                                                                        �             


           �   }�    �                  '                           +                     R�               ������������  R�  +������������   	������������    ����������������������������������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" A C 6               	                  � ��/} �c@                                                                                                                                                                                                                                                                                      �Y  "$)F        c      e      k                  m            m                                                                                                                                                                                                                                                                                                                                                                                                         ( =  (=  �  � #��  � #��  EZm �̎�G��d�� �N 5��� ^�����������������������                 } � : ( i
        	 �   &  AG� �   f                    �                                                                                                                                                                                                                                                                                                                                      p B I   $     	                !��                                                                                                                                                                                                                            Y   �� �� ����      �� B 	     ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ������������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     9      0   �                         B     �  �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$     `d ��     `d �$ ^$ �@          �� �         9   ����   ���@ ��  ���@ �$ ^$   �    �� @ 
i   ���8   (   $     c@ �d �� c@ �d �$ g �  ��g  �      �   d   %���� e�����   g��� 	 �     f ^�   `     ��         %      �������2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                               s   D   O   w   w   v   u   f   T   �   �              3@  DDp ��4 ��tp��wpO�tpdfwGfeTwfeWwfUFwdUFweTfp�DDp���p���@�w�p   C   D   O   D   w   u   U   U  F  d  f   f   D   �   �   �DD ���7���uP��e`O�V ffg ffG Ufw UU� FUN dFw ffp DDp ��p ��@ w�p  C4 4D@O�C���O�Dt�GVfeVfdFfdFfdUfffUfffwFff�DDD���� ���                    0   G   W   W   U   E   E   w   �   �   @    fg D� O�� �� w�}�w��}����������M���M���M��������y�                    �   �   �   �   �   �   �   �   ~   w       ���w���w���~���~�DMw�������������y�                        w���w}��wt��wt��w}M�����������   M   M   ~�  p�  p   p   p      �   �   �   �               vd  eVp ffpw�Op���w���G���M�}�                                     v   ub  ub  f   `   P               "  f  U` wfP        p   p   p   p   p   p   p   p                               C4 �y�                              f  vU`vf`D�O������p}�w�  ?�  ?�  ?�  33  3#                                      f  Ug                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  " ! " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "!  " ! " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """ "!    " ""   "   "   "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        ̰ �� ̻ {�����vz� w��  ��  ��  ̘  	�  
� "��,̻�"�� "#3  34  D  
�  �  " "" """ ! ��  ��                               ˹� �ɩ ��� �͋ ��� ��� ��̀��Ȑ���лܹнȝ0ݙ�@43�PCD�@@E�@ E�@ U�� H�  K�  �   ��    �� "�" ���                          �  �   ��  �  ��                �   �   �   "   "   "  !�    ��                              �                        ���� ��� ����                              "  .���"    �     �                         � ���� ��   � � �                                                                                                                                  �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �   �   "   "   "  !�    ��                           ���                         �  ��                    �����                       ��                                 � ���� ��   � � �           � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                         
�� ɪ�̚���ə���̚���ɍ��������̻�̲��"X��
Y���C9�UC33�DC3��  ��  �  ��� "�  ��� ��   �  �    ��  ��  ��  ��  w}  ww  ��  ��� ���������ɋ��˽��˽���� �̰ ̸� ��� �30 333 333 330 TD0 ��� �  ��  ��  ̲/ ����"/ �� � ��     � �  �  ��  �  �   �   �      	  *  ,  +   "   �            �   ������  ��                   �                        ���� ��� ����                               � ��                  �  �˰ ��� �wp ���                                                                                                                                                                               � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �           �     �                                                                                                                                                                                            �  �˰ �̰ �˰ ܻ� �p
���٪����������������� ۼ� �� ��  ��  ��  H�  X� �T �T �U �[  ̻  ��  �  ��   �  "  �"     �   �  �     �   � �  � ��� �ɨ ۚ� ��� �۰ ��  ��  ̘  ��  �C  T@  D   K�  �   "�    ��� ��� ��  ��  /�  /  /    ""�����                                        �� �  �        �  �  ��  �   �                              �   �                      �������  ���    �                    ��� ���� ��                                                                                                                                                                                                       �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �                         �               �  ���ݼ�������ک����   �   �           �   ̰  �˰                                                                                                                                                                                                       �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �      �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                       � ��                  �  �˰ ��� �wp ���                                                                                                                                                                 �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                    "   "       �  �       "  "/�����                     �   ��  �   ��   �       �                                                                                                                                  ̻  ��  rb  wg 
�w ���
���ɛ������̽�̪��̙���̻̽̽���٘"#3 ""DR�U� T� �� 	��  ��  ,� "� "� ""��""�������� �  ��   �   p   z   ��  ��  ��� �̹ �ؚ �ک ��������������32"�D2" UR" EU@ EU@ 4U@ K˰ 
�� ��  �   "   ""  "" ��"/���� �� �     ��  ��  ��  ��  ��  ��  �                             �� ̽   �   �  ��� ��  ��  �   ��        �  ��� ̻� ��� rbp wgz�                    �    ���� �              �  �� ��  �    � ���                                                                                                                                                                                            �gz�������������̼�ˍ��̭��̘ۼ��ۻ��ۼ��˙���4R"#EU"�4UR�TUDN�U � " �"" �"/ �"/�������    �                      �   ��  ̹  ��� ة� ��� ��� �� �"" �"" 3" CR  UP  UT  UT  ET� ��� 
�� ��  �"  "  "   ""�"����� �� � �     ��  ��  �         
   �   �   �   �   �   �   	                        ��  ��  �   �                        �  ��� ̻� ��� rbp wgz�       ����������             ��  �   ��  �                             �  �˰ ��� �wp ���                                                                                                                                                                  ̻  ��  rb  wg 
�w ���
���ɛ������̽�̪��̙���̻̽̽���٘"#3 ""DR�U� T� �� 	��  ��  ,� "� "� ""��""�������� �  ��   �   p   z   ��  ��  ��� �̹ �ؚ �ک ��������������32"�D2" UR" EU@ EU@ 4U@ K˰ 
�� ��  �   "   ""  "" ��"/���� �� �     ��  ��  ��  ��  ��  ��  �                             �� ̽   �   � � �  ��� ��  �    "   "   "  �� ��                   ����������                                ��  ��  ���                   ���                                                                                                                                                                                                �� ��
������ɻ��ܻ� ��� �"�"+�.+� .�� �8 �3 �S DNC E^@E^0������
���"� "  "  " � ���� � ���  �̰ ۼ� �۰ rbp wgp �v� ��������������������̻ڙ˻٪��ݙ˽�̙�+�32" 4"$@"$@ DDP DU@ �� �  "  "  "   "/����� ����                     "   "   �    �   �                          �   �  ��� ��  ��  �   ��        �  ��� ̻� ��� rbp wgz�        �   �  �  �   �               �   �               �� ����� ���  �                   �   �   �   �   �   �                                                                                                                                                �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(XxLL����������D����3333DDDD w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""����������A������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(""""�������I�I������ �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�""""�������I��D���I������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`�D�M�D���M������3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(MD�M�A�����MD�����3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(�""""�����AMAD������ � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(�""""������������������ � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
2� � �
�	ckjX{ krhKkV �[ k^ � �B�^ � B�V �	CP �
CX � C Q �C!P �C#[ �J�D � J�T �J�< �KP � K` �KP � K` � KS � KT �  Kt �  Kh �  KX �  Kr{ *� �b"� �b*� ��"� �� "� �y � �y 
� �r 
� �?#� �? 
� �5%"� �5 &"� �%'� �% 
� �)� � 
� � 
� �',"� �' -"� �.� � 
� �0� � 
� �2� � 
� � 
� � 
� � �6" � � 7!� � �8"" � �9!� � �:!� � �;" �<*$7 �=* O �  *O � * O3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0�������������������������������������������C�G�X�R�K�_��C�G�R�G�V�Y�Q�O� � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� �� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            