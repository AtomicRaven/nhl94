GST@�                                                            \     �                                               
     X   ��J             j�������J���ʲ���������    ����        x9      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"   "D�j��
� " ��
  _                                                                               ����������������������������������      ��    =ob 0Q 4o 1 1  +4   '       �	 
                �	� �7 �V  �	                 nn 	)         :8�����������������������������������������������������������������������������������������������������������������������������b  Qb    14  4c  c   c           	  
        	   
        �G  �   (  (                  nn  )1          88 �����������������������������������������������������������������������������                                      �  9�   @  #   �   �                                                                                'w w  	n)n  )n1n    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������      �L�\I��.Y|0
I�|T����@��9@8]�W3� T0 k� � E�$E? �$1`1	u1�4 � ��?    � %��  �L�\I��.Y|0
I�|U����@��9@8]�W3� T0 k� �0E�4E? �$1`1	u1�4 � ��?    � %��  �P�`I��.Y|0
I�|V����@��9@8]�W3� T0 k� �DE�HE? �$1`1	u1�4 � ��?    � %��  �P�`I��.Y|0
I�|W����@��9@8]�W3� T0 k� �XE�\E? �$1`1	u1�4 � ��?    � %��  �T�`I��.Y|0
I�|W����@��9@8]�W3� T0 k� lE�pE? �$1`1	u1�4 �  ��?    � %��  �X�dI��.Y|0
I�|X����@��9@9]�W3� T0 k� �F��F? �$1`1	u1�4 �  ,�?    � %��  �\�dI��.Y|0
I�|X����?��9@9]�W3� T0 k� �F��F? �$1`1	u1�4 �  ��?    � %��  �`�hI��/Y|0
I�|Y����?��9@9]�W3� T0 k� �F��F? �$1`1	u1�4 �  ��?    � %��  �`�lI��/Y|0
I�|Y����?��9@9]�W3� T0 k� �F��F? �$1`1	u1�4 � ��?    � %��  �d�lI��/Y|0
I�|Z����?��9@9]�W3� T0 k� ��F��F? �$1`1	u1�4 � ��?    � %��  �h�pI��/Y|0
I�|Z����?��9@9]�W3� T0 k� ��F��F? �$1`1	u1�4 � ��?    � %��  �l�tI��/Y|0
I�|Z����?��9@9]�W3� T0 k� ��F��F? �$1`1	u1�4 � ��?    � %��  �p�xI��/Y|0
I�|[����?��9@9]�W3� T0 k� �G�G? �$1`1	u1�4 � ��?    � %��  �t�xI��/Y|0
I�|[����?��9@:]�W3� T0 k� �G�G? �$1`1	u1�4 � ��?    � %��  �x�|I��/Y|0
I�|[����?��9@:]�W3� T0 k� (G�,G? �$1`1	u1�4 � ��?    � %��  �|��I��/Y|0
I�|[����?��9@:]�W3� T0 k� <G�@G? �$1`1	u1�4 � ��?    � %��  ����I��/Y|0
I�|[����?��9@:]�W3� T0 k� PG�TG? �$1`1	u1�4 � ��?    � %��  ����I��.Y|0
I�|[����?��9@;]�W3� T0 k� dG�hG? �$1`1	u1�4 � ��?    � %��  ����I��.Y|0
I�|[����?��9@;]�W3� T0 k� tG�xG? �$1`1	u1�4 � ��?    � %��  ����I��.Y|0
I�|[����?��9@ ;]�W3� T0 k� ��G��G? �$1`1	u1�4 � ��?    � %��  ����I��.Y|0
I�|[����?��9@ <]�W3� T0 k� ��H��H? �$1`1	u1�4 � (�?    � %��  ��͜I��.Y|0
I�|[����?��9@$<]�W3� T0 k� ��G��G? �$1`1	u1�4 � ��?    � %��  �ͤI��.Y|0
I�|[����?��9@$<]�W3� T0 k� ��G��G? �$1`1	u1�4 � ��?    � %��  �ͨI��.Y|0
A�|[����?��9@$<]�W3� T0 k� ��G��G? �$1`1	u1�4 � ��?    � %��  �ͰI��.Y|0
A�|[����?��9@(=]�W3� T0 k� ��F��F? �$1`1	u1�4 � ��?    � %��  �ʹI��-Y|0
A�|[����>��9@(=]�W3� T0 k� 4�F��F? �$1`1	u1�4 � ��?    � %��  �ʹI��-Y|0
A�|[����>��9@(=]�W3� T0 k� 4�F��F? �$1`1	u1�4 � ��?    � %��  �ͼI� -Y|0
A�|[����>��8@,>]�W3� T0 k� 4|F��F? �$1`1	u1�4 � ��?    � %��  ���H� -Y|0
BN|[����>��8@,>]�X3� T0 k� 4xE�|E? �$1`1	u1�4 � ��?   � %��  ���H�-Y|0
BN|[����>��8@,>]�X3� T0 k� 4pE�tE? �$1`1	u1�4 � ��?    � %��  ���H�-Y|0
BN|[����>��8@0?]�X3� T0 k� �lE�pE? �$1`1	u1�4 � ��?    � %��  ���G�-Y|0
BN|[����>��8@0?]�Y3� T0 k� �hD�lD? �$1`1	u1�4 � ��?   � %��  ���G�-Y|0
BN|[����>��8@0?]�Y3� T0 k� �dD�hD? �$1`1	u1�4 � ��?    � %��  ���G�-Y|0
BN|[���� >��8@4?]�Y3� T0 k� �`D�dD? �$1`1	u1�4 �  ��?    � %��  ���G�-Y|0
BN|[���� >��8@4@]�Y3� T0 k� �XC�\C? �$1`1	u1�4 �  ��?    � %��  ���G�,Y|0
BN|[���� >��8@4@]�Z3� T0 k� �TC�XC? �$1`1	u1�4 �  .�?    � %��  ���G�,Y|0
BN|[����$=��8@4@]�Z3� T0 k� �PC�TC? �$1`1	u1�4 �  ��?    � %��  ���H�,Y|0
BN|[����$=��8@8@]�Z3� T0 k� �LC�PC? �$1`1	u1�4 �  ��?    � %��  ���H�,Y|0
@|[����(=��8@8A]�Z3� T0 k� �HB�LB? �$1`1	u1�4 �  ��?    � %��  ���H�,Y|0
@|[����,<��8@8A]�[3� T0 k� �DB�HB? �$1`1	u1�4 �  ��?    � %��  ���H� ,Y|0
@|[����,<��8@<A]�[3� T0 k� �<B�@B? �$1`1	u1�4 �  ��?    � %��  ���I� ,Y|0
@|[����0<��8@<A]�[3� T0 k� �8A�<A? �$1`1	u1�4 �  ��?    � %��   � I�$,Y|0
@|[����0;��8@<B]�[3� T0 k� �4A�8A? �$1`1	u1�4 �  ��?    � %��  !�J�$,Y|0
@|[����4;��8@<B]�\3� T0 k� �0A�4A? �$1`1	u1�4 �  ��?    � %��  -!�J�(,Y|0
@|[����4;��8@@B]�\3� T0 k� �,@�0@? �$1`1	u1�4 �  ��?    � %��  -"�K�,,Y|0
@|[����8:��8@@B]�\3� T0 k� �(@�,@? �$1`1	u1�4 �  ��?    � %��  -#�K�,+Y|0
@|[����8:��8@@C]�\3� T0 k� �$@�(@? �$1`1	u1�4 �  ��?    � %��  - $�L�0+Y|0
@|[����<:��8@@C]�]3� T0 k� �@� @? �$1`1	u1�4 �  ��?    � %��  -(%�L�0+Y|0
@|[����<9��8@DC]�]3� T0 k� �?�?? �$1`1	u1�4 �  ��?    � %��  -0&	> L�4+Y|0
@|[����@9��8@DC]�]3� T0 k� �?�?? �$1`1	u1�4 �  ��?    � %��  -4'	>$M�4+Y|0
@|[����@9��8@DC]�]3� T0 k� �?�?? �$1`1	u1�4 �  ��?    � %��  -<(	>(M�4+Y|0
@|[����D8��8@DD]�]3� T0 k� �>�>? �$1`1	u1�4 �  ��?   � %��  -@)	>(M�8+Y|0
@|[����D8��8@HD]�^3� T0 k� �>�>? �$1`1	u1�4 �  ��?    � %��  -H*	>,M�8+Y|0
@|[����H8��8@HD]�^3� T0 k� �>�>? �$1`1	u1�4 �  ��?    � %��  -P+	N0M�<+Y|0
@|[����H8��8@HD]�^3� T0 k� ��>� >? �$1`1	u1�4 �  ��?    � %��  �T,	N4M�<+Y|0
@|[����L7��8@HD]�^3� T0 k� ��=��=? �$1`1	u1�4 �  ��?    � %��  �T,	N4M�@+Y|0
@|[����L7��9@LE]�^3� T0 k� ��=��=? �$1`1	u1�4 �  ��?    � %��  �X,	N8M�@+Y|0
@|[����P7��9@LE]�_3� T0 k� ��=��=? �$1`1	u1�4 �  ��?    � %��  �\,	N8N�D+Y|0
@|[����P6��:@LE]�_3� T0 k� ��<��<? �$1`1	u1�4 �  ��?    � %��  �\-�<N�D+Y|0
@|[����T6��:@LE]�_3� T0 k� ��<��<? �$1`1	u1�4 �  ��?    � %��  �\-�@N H*Y|0
@|[����T6��<@PF]�_3� T0 k� ��<��<? �$1`1	u1�4 �  ��?    � %��  �`-�DN H*Y|0
@|[����X5��<@PF]�`3� T0 k� ��;��;? �$1`1	u1�4 �  ��?    � %��  �d-�HN L*Y|0
@|[����X5��=@PF]�`3� T0 k� ��;��;? �$1`1	u1�4 �  ��?    � %��  �h.�LO L*Y|0
@|[����\5��>@PF]�`3� T0 k� ��;��;? �$1`1	u1�4 �  ��?    � %��  �l.�PO L*Y|0
@|[����\5��>@PF]�`3� T0 k� ��;��;? �$1`1	u1�4 �  ��?    � %��  �p/�PO P*Y|0
@�\����\4��?@TF]�`3� T0 k� ��:��:? �$1`1	u1�4 �  ��?    � %��  t0�PO P*Y|0
@�\����`4��?@TG]�`3� T0 k� ��:��:? �$1`1	u1�4 �  ��?    � %��  x0�TO T*Y|0
@�\����`4��@@TG]�a3� T0 k� ��:��:? �$1`1	u1�4 �  ��?    � %��  |1�TO T*Y|0
K��\����d4��A@TG]�a3� T0 k� ��9��9? �$1`1	u1�4 �  ��?    � %��  �1XO T*Y|0
K��]����d4��A@TG]�a3� T0 k� ��9��9? �$1`1	u1�4 �  ��?    � %��  �2XO X*Y|0
K��]����d3��B@TG]�a3� T0 k� ��9��9? �$1`1	u1�4 �  ��?    � %��  �3\O X*Y|0
K��]����h3��B@XG]�a3� T0 k� ��9��9? �$1`1	u1�4 �  ��?    � %��  �3\O X*Y|0
K��]����h3��C@XH]�a3� T0 k� ��8��8? �$1`1	u1�4 �  ��?    � %��  �4`O \*Y|0
K��]����h3��D@XH]�b3� T0 k� ��8��8? �$1`1	u1�4 �  ��?    � %��  �4`O \*Y|0
K��^����l3��D@XH]�b3� T0 k� ��8��8? �$1`1	u1�4 �  ��?    � %��  �4`O \*Y|0
K��^����l2��E@XH]�b3� T0 k� ��8��8? �$1`1	u1�4 �  ��?   � %��  �5dO `)Y|0
K��^����l2��F@XH]�b3� T0 k� ��7��7? �$1`1	u1�4 �  ��?    � %��  �5dO `)Y|0
K��^����p2��G@\H]�b3� T0 k� ��7��7? �$1`1	u1�4 �  ��?    � %��  �6dO `)Y|0
K��^����p2��G@\H]�b3� T0 k� ��7��7? �$1`1	u1�4 �  ��?    � %��  �7dO d)Y|0
K��_����p2��H@\I]�b3� T0 k� ��6��6? �$1`1	u1�4 �  ��?    � %��  �8dO d)Y|0
K��_����t1��I@\I]�c3� T0 k� ��6��6? �$1`1	u1�4 �  ��?    � %��  �8dO d)Y|0
K��_����t1��J@\I]�c3� T0 k� ��6��6? �$1`1	u1�4 �  ��?    � %��  �9dO h)Y|0
K��_����t1��J@\I]�c3� T0 k� ��6��6? �$1`1	u1�4 �  ��?    � %��  �:dO h)Y|0
K��_����t1��K@`I]�c3� T0 k� �|5��5? �$1`1	u1�4 �  ��?    � %��  �;dO h)Y|0
K��`����x1��L@`I]�c3� T0 k� �x5�|5? �$1`1	u1�4 �  ��?    � %��  �< ndO h)Y|0
K��`����x1��L@`I]�c3� T0 k� �t5�x5? �$1`1	u1�4 �  ��?    � %��  �< ndO l)Y|0
K��`����x0��M@`I]�c3� T0 k� �p5�t5? �$1`1	u1�4 �  ��?    � %��  �= ndO l)Y|0
K��`����|0��N@`J]�c3� T0 k� �l4�p4? �$1`1	u1�4 �  ��?    � %��  -�> ndO l)Y|0
K��`����|0��N@`J]�d3� T0 k� �d4�h4? �$1`1	u1�4 �  ��?    � %��  -�> ndO l)Y|0
K��`����|0��O@`J]�d3� T0 k� �`4�d4? �$1`1	u1�4 �  ��?    � %��  -�? ndO p)Y|0
K��a����|0��O@`J]�d3� T0 k� �\4�`4? �$1`1	u1�4 �  ��?    � %��  -�@ ndO p)Y|0
K��a�����0��P@dJ]�d3� T0 k� �X3�\3? �$1`1	u1�4 �  ��?    � %��  -�A�dO p)Y|0
K��a�����/��Q@dJ]�d3� T0 k� �T3�X3? �$1`1	u1�4 �  ��?    � %��  ��B�dO p)Y|0
K��a�����/��Q@dJ]�d3� T0 k� �P3�T3? �$1`1	u1�4 �  ��?    � %��  ��C�dO t)Y|0
K��a�����/��R@dJ]�d3� T0 k� �L3�P3? �$1`1	u1�4 �  ��?    � %��  ��D�dO t)Y|0
K��a�����/��R@dK]�d3� T0 k� �H2�L2? �$1`1	u1�4 �  ��?    � %��  ��D�dO t)Y|0
K��b�����/��S@dK]�d3� T0 k� �D2�H2? �$1`1	u1�4 �  ��?    � %��  ��E�dO t)Y|0
K��b�����/��T@dK]�e3� T0 k� �@2�D2? �$1`1	u1�4 �  ��?    � %��  ��F�dO x)Y|0
K��b�����/��T@dK]�e3� T0 k� �<2�@2? �$1`1	u1�4 �  ��?    � %��  � G�dO x)Y|0
K��b�����.��U@hK]�e3� T0 k� �81�<1? �$1`1	u1�4 �  ��?    � %��  �H�dO x)Y|0
K��b�����.��U@hK]�e3� T0 k� �41�81? �$1`1	u1�4 �  ��?    � %��  �I�dO x)Y|0
K��b�����.��V@hK]�e3� T0 k� �01�41? �$1`1	u1�4 �  ��?    � %��  �I�dO |)Y|0
K��b�����.��V@hK]�e3� T0 k� �,1�01? �$1`1	u1�4 �  ��?    � %��  �J�dO |)Y|0
K��c�����.��V@hK]�e3� T0 k� �(0�,0? �$1`1	u1�4 �  ��?    � %��  �K�dO |(Y|0
K��c�����.��V@hK]�f3� T0 k� �$0�(0? �$1`1	u1�4 �  ��?    � %��  �L�dO |(Y|0
K��c�����.��V@hL]�f3� T0 k� � 0�$0? �$1`1	u1�4 �  ��?    � %��  � L�dO |(Y|0
K��c�����.��V@hL]�f3� T0 k� �/� /? �$1`1	u1�4 �  ��?    � %��  �$M�dO �(Y|0
K��c�����-��W@hL]�f3� T0 k� �/�/? �$1`1	u1�4 �  ��?    � %��  �$M�hO �(Y|0
K��c�����-��W@lL]�g3� T0 k� �/�/? �$1`1	u1�4 �  ��?    � %��  �$M�hO �(Y|0
K��c�����-��W@lL]�g3� T0 k� �/�/? �$1`1	u1�4 �  ��?    � %��  �(N�lO �(Y|0
K��c�����-��W@lL]�g3� T0 k� �.�.? �$1`1	u1�4 �  ��?    � %��  �(O�lO �(Y|0
K��d�����-��X@lL]�g3� T0 k� �.�.? �$1`1	u1�4 �  ��?    � %��  �,O�pO �(Y|0
K��d�����-��X@lL]�h3� T0 k� �.�.? �$1`1	u1�4 �  ��?    � %��  �,P�pO �(Y|0
K��d�����-��X@lL]�h3� T0 k� � .�.? �$1`1	u1�4 �  ��?    � %��  �,P�pO �(Y|0
K��d�����-��X@lL]�h3� T0 k� ��.� .? �$1`1	u1�4 �  ��?    � %��  �0Q�tO �(Y|0
K��d�����-��X@lL]�h3� T0 k� ��-��-? �$1`1	u1�4 �  ��?    � %��  �0Q�tO �(Y|0
K��d�����,��Y@lL]�i3� T0 k� ��-��-? �$1`1	u1�4 �  ��?    � %��  �0R�xP �(Y|0
K��d�����,��Y@lM]�i3� T0 k� ��-��-? �$1`1	u1�4 �  ��?    � %��  �4R�xP �(Y|0
K��d�����,��Y@lM]�i3� T0 k� ��-��-? �$1`1	u1�4 �  ��?    � %��  �4S�xP �(Y|0
K��d�����,��Y@pM]�i3� T0 k� ��,��,? �$1`1	u1�4 �  ��?    � %��  �8S�|P �(Y|0
K��e�����,��Y@pM]�i3� T0 k� ��,��,? �$1`1	u1�4 �  ��?    � %��  �8T�|P �(Y|0
K��e�����,��Z@pM]�j3� T0 k� ��,��,? �$1`1	u1�4 �  ��?    � %��  �8T΀P �(Y|0
K��e�����,��Z@pM]�j3� T0 k� ��,��,? �$1`1	u1�4 �  ��?    � %��  �<U΀P �(Y|0
K��e�����,��Z@pM]�j3� T0 k� ��+��+? �$1`1	u1�4 �  ��?    � %��  �<U΀P �(Y|0
K��e�����,��Z@pM]�j3� T0 k� ��+��+? �$1`1	u1�4 �  ��?    � %��  �<V΄P �(a�0
K��e�����,��Z@pM]�j"�� T0 k� ��+��+? �$1`1	u1�4 �  ��?    � %��  �@V΄P �(a�0
K��e�����,��[@pM]�k"�� T0 k� ��+��+? �$1`1	u1�4 �  ��?    � %��  �@W΄P �(a�0
K��e�����+��[@pM]�k"�� T0 k� ��*��*? �$1`1	u1�4 �  ��?    � %��  �@WΈP �(a�0
K��e�����+��[@pM]�k"�� T0 k� ��*��*? �$1`1	u1�4 �  ��?    � %��  �DWΈP �(a�0
K��e�����+��[@pM]�k"�� T0 k� ��*��*? �$1`1	u1�4 �  ��?    � %��  �DXΈP �(a�0
K��e�����+��[@pM]�k"�� T0 k� ��*��*? �$1`1	u1�4 �  ��?    � %��  �DXΌP �(a�0
K��e�����+��[@pN]�l"�� T0 k� ��)��)? �$1`1	u1�4 �  ��?    � %��  �HYΌP �(a�0
@�e�����+��\@tN]�l"�� T0 k� ��)��)? �$1`1	u1�4 �  ��?    � %��  �HYΌP��(a�0
@�e�����+��\@tN]�l"�� T0 k� ��)��)? �$1`1	u1�4 �  ��?    � %��  �HZΐP��(a�0
@�e�����+��\@tN]�l"�� T0 k� ��)��)? �$1`1	u1�4 �  ��?    � %��  �HZΐP��(a�0
@�e�����+��\@tN]�l"�� T0 k� ��(��(? �$1`1	u1�4 �  ��?    � %��  �LZΐP��(Y|0
@�e�����+��\@tN]�l3� T0 k� ��(��(? �$1`1	u1�4 �  ��?    � %��  �L[ΔP��(Y|0
K��e�����+��\@tN]�m3� T0 k� ��(��(? �$1`1	u1�4 �  ��?    � %��  �L[ΔP��(Y|0
K��e�����+��\@tN]�m3� T0 k� ��(��(? �$1`1	u1�4 �  ��?    � %��  �P[ΔP��(Y|0
K��e�����+��]@tN]�m3� T0 k� ��(��(? �$1`1	u1�4 �  ��?    � %��  �P\ΘP��(Y|0
K��e�����*��]@tN]�m3� T0 k� ��'��'? �$1`1	u1�4 �  ��?    � %��  �P\ΘP��(Y|0
K��e�����*��]@tN]�m3� T0 k� ��'��'? �$1`1	u1�4 �  ��?    � %��  �P]ΘP��(Y|0
K��e�����*��]@tN]�m3� T0 k� ��'��'? �$1`1	u1�4 �  ��?    � %��  �T]ΘP��(Y|0
K��e�����*��]@tN]�n3� T0 k� ��'��'? �$1`1	u1�4 �  ��?    � %��  �T]ΜP��(Y|0
K��e�����*��]@tN]�n3� T0 k� ��&��&? �$1`1	u1�4 �  ��?    � %��  �T^ΜP��(Y|0
K��e�����*��]@tN]�n3� T0 k� ��&��&? �$1`1	u1�4 �  ��?    � %��  �T^ΜP��(Y|0
K��e�����*��^@tN]�n3� T0 k� ��&��&? �$1`1	u1�4 �  ��?    � %��  �X^��P��(a�0
K��e�����*��^@xN]�n"s� T0 k� �|&��&? �$1`1	u1�4 �  ��?    � %��  �X_��P��(a�0
K��e�����*��^@xO]�n"s� T0 k� �x%�|%? �$1`1	u1�4 �  ��?    � %��  �X_��P��(a�0
K��e�����*��^@xO]�n"s� T0 k� �t%�x%? �$1`1	u1�4 �  ��?    � %��  �X_��P��(a�0
K��e�����*��^@xO]�n"s� T0 k� �p%�t%? �$1`1	u1�4 �  ��?    � %��  �\_��P��(a�0
K��e�����*��^@xO]�o"s� T0 k� �p%�t%? �$1`1	u1�4 �  ��?    � %��  �\`��P��(a�0
K��e�����*��^@xO]�o"s� T0 k� �l%�p%? �$1`1	u1�4 �  ��?    � %��  �\`��P��(a�0
K��e�����*��^@xO]�o"s� T0 k� �h$�l$? �$1`1	u1�4 �  ��?    � %��  �\a��P��(a�0
K��e�����*��_@xO]�o"s� T0 k� �d$�h$? �$1`1	u1�4 �  ��?    � %��  �`a��P��(a�0
K��e�����*��_@xO]�o"s� T0 k� �`$�d$? �$1`1	u1�4 �  ��?    � %��  �`a��P��(a�0
K��e�����*��_@xO^ o"s� T0 k� �\$�`$? �$1`1	u1�4 �  ��?    � %��  `a��P��(a�0
K��e�����*��_@xO^ o"s� T0 k� �X#�\#? �$1`1	u1�4 �  ��?   � %��  `a��P��(Y|0
K��f�����)��_@xO^ p3� T0 k� �T#�X#? �$1`1	u1�4 �  ��?    � %��  `b n�P��(Y|0
K��f�����)��_@xO^ p3� T0 k� �P#�T#? �$1`1	u1�4 �  ��?    � %��  `b n�P��(Y|0
K��f�����)��_@xO^ p3� T0 k� �L#�P#? �$1`1	u1�4 �  ��?    � %��  db n�P��(Y|0
K��f�����)��_@xO^ p3� T0 k� �H"�L"? �$1`1	u1�4 �  ��?    � %��  �db n�P��(Y|0
K��f�����)��_@xO^ p3� T0 k� �H"�L"? �$1`1	u1�4 �  ��?    � %��  �hc n�P��(Y|0
K��f�����)��_@xO^ p3� T0 k� �D"�H"? �$1`1	u1�4 �  ��?    � %��  �hc n�P��(Y|0
K��f�����)��`@xO^ p3� T0 k� �@"�D"? �$1`1	u1�4 �  ��?    � %��  �hc n�P��(Y|0
K��f�����)��`@xO^ p3� T0 k� �<"�@"? �$1`1	u1�4 �  ��?    � %��  �ld �P��(Y|0
K��f�����)��`@xO^ p3� T0 k� �8!�<!? �$1`1	u1�4 �  ��?    � %��  ~ld �P��(Y|0
K��f�����)��`@|O^ q3� T0 k� �4!�8!? �$1`1	u1�4 �  ��?    � %��  ~ld �P��(Y|0
K��f�����)��`@|O^ q3� T0 k� �0!�4!? �$1`1	u1�4 �  ��?    � %��  ~ld �P��(Y|0
K��f�����)��`@|O^ q3� T0 k� �,!�0!? �$1`1	u1�4 �  ��?    � %��  ~le �P��(Y|0
K��f�����)��`@|O^ q3� T0 k� �(!�,!? �$1`1	u1�4 �  ��?    � %��  ~le �P��(Y|0
K��f�����)��`@|P^ q3� T0 k� �( �, ? �$1`1	u1�4 �  ��?    � %��  ~pe �P��(Y|0
K��f�����)��`@|P^ q3� T0 k� �$ �( ? �$1`1	u1�4 �  ��?    � %��  ~pe �P��(Y|0
K��f�����)��`@|P^ q3� T0 k� �  �$ ? �$1`1	u1�4 �  ��?    � %��  ~pe �P��'Y|0
K��f�����)��a@|P^ q3� T0 k� � �  ? �$1`1	u1�4 �  ��?    � %��  ~pf �P��'Y|0
K��f�����)��a@|P^ q3� T0 k� ��? �$1`1	u1�4 �  ��?    � %��  ~tf �P��'Y|0
K��f�����)��a@|P^q3� T0 k� ��? �$1`1	u1�4 �  ��?    � %��  �tf �P��'Y|0
K��g�����)��a@|P^q3� T0 k� ��? �$1`1	u1�4 �  ��?    � %��  �tf �P��'Y|0
K��g�����)��a@|P^r3� T0 k� ��? �$1`1	u1�4 �  ��?    � %��  �tf �P��'Y|0
K��g�����)��a@|P^r3� T0 k� ��? �$1`1	u1�4 �  ��?    � %��  �xf �P��'Y|0
K��g�����)��a@|P^r3� T0 k� ��? �$1`1	u1�4 �  ��?    � %��  �xg �P��'Y|0
K��g�����)��a@|P^r3� T0 k� ��? �$1`1	u1�4 �  ��?    � %��  �xg �P��'Y|0
K��g�����)��a@|P^r3� T0 k� � �? �$1`1	u1�4 �  ��?    � %��  �xg �P��'Y|0
K��g�����)��a@|P^r3� T0 k� ��� ? �$1`1	u1�4 �  ��?    � %��  �|g �P��'Y|0
K��g�����(��a@|P^r3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  �|g �P��'Y|0
K��g�����(��a@|P^r3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  �|h �P��'Y|0
K��g�����(��a@|P^r3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  �|h �P��'Y|0
K��g�����(��b@|P^r3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  �|h �P��'Y|0
K��g�����(��b@|P^r3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��h �P��'Y|0
K��g�����(��b@|P^r3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��h �P��'Y|0
K��g�����(��b@|P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��h��P��'Y|0
K��g�����(��b@|P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��h��P��'Y|0
K��g�����(��b@|P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��i��P��'Y|0
K��g�����(��b@�P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��i��P �'Y|0
K��g�����(��b@�P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��i��P �'Y|0
@n�g�����(��b@�P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��i��P �'Y|0
@n�g�����(��b@�P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��i��P �'Y|0
@n�g�����(��b@�P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��i��P �'Y|0
@n�g�����(��b@�P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��j��P �'Y|0
@n�g�����(��b@�P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��j��P �'Y|0
E��f�����(��b@�P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��j��P �'Y|0
E��f�����(��b@�P^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��j��P �'Y|0
E��f�����(��c@�Q^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��j��P �'Y|0
E��e�����(��c@�Q^s3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��j��P �'Y|0
E��e�����(��c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��j��P �'Y|0
K��d�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��j��P �'Y|0
K��d�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��d�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��c�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��c�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��c�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��b�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��b�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��b�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��a�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��a�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��l��P��'Y|0
K��a�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ��l��P��'Y|0
K��`�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ~�l��P��'Y|0
K��`�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ~�l��P��'Y|0
K��`�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ~�l��P��'Y|0
K��`�����(� c@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ~�l��P��'Y|0
K��_�����(� d@�Q^t3� T0 k� ����? �$1`1	u1�4 �  ��?    � %��  ~�l��P��'Y|0
K��_�����(� d@�Q^t3� T0 k� �|��? �$1`1	u1�4 �  ��?    � %��  ~�l��P��'Y|0
K��_�����(� d@�Q^u3� T0 k� �x�|? �$1`1	u1�4 �  ��?    � %��  N�l��P��'Y|0
K��_�����(� d@�Q^u3� T0 k� �t�x? �$1`1	u1�4 �  ��?    � %��  N�l��P��'Y|0
K��^�����(� d@�Q^u3� T0 k� �t�x? �$1`1	u1�4 �  ��?    � %��  N�l��P��'Y|0
K��^�����(� d@�Q^u3� T0 k� �p�t? �$1`1	u1�4 �  ��?    � %��  N�l��P��'Y|0
K��^�����(� d@�Q^u3� T0 k� �l�p? �$1`1	u1�4 �  ��?    � %��  N�l��P��'Y|0
K��]�����(� d@�Q^u3� T0 k� �h�l? �$1`1	u1�4 �  ��?    � %��  ��l��P��'Y|0
K��]�����(� d@�Q^u3� T0 k� �d�h? �$1`1	u1�4 �  ��?    � %��  ��l��P��'Y|0
K��]�����(� d@�Q^u3� T0 k� �d�h? �$1`1	u1�4 �  ��?    � %��  ��l��P��'Y|0
K��]�����(�d@�Q^u3� T0 k� �`�d? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��\�����(�d@�Q^u3� T0 k� �\�`? �$1`1	u1�4 �  ��?    � %��  ��k��P��'Y|0
K��\�����(�d@�Q^u3� T0 k� �X�\? �$1`1	u1�4 �  ��?    � %��  n�k��P��'Y|0
K��\�����(�d@�Q^u3� T0 k� �X�\? �$1`1	u1�4 �  ��?    � %��  n�j��P��'Y|0
K��\�����(�d@�Q^u3� T0 k� �T�X? �$1`1	u1�4 �  ��?    � %��  n�j��P��'Y|0
K��\�����(�d@�Q^u3� T0 k� �P�T? �$1`1	u1�4 �  ��?    � %��  n�i��P��'Y|0
K��[�����(�d@�Q^u3� T0 k� �L�P? �$1`1	u1�4 �  ��?    � %��  n�i��P��'Y|0
K� [�����(�d@�Q^u3� T0 k� �H�L? �$1`1	u1�4 �  ��?    � %��  n�h��P��'Y|0
K� [�����(�d@�Q^u3� T0 k� �H�L? �$1`1	u1�4 �  ��?    � %��  n�h��P��'Y|0
K� [�����(�d@�Q^u3� T0 k� �D�H? �$1`1	u1�4 �  ��?    � %��  n�g��P��'Y|0
K� [�����(�d@�Q^u3� T0 k� �@�D? �$1`1	u1�4 �  ��?    � %��  n�g��P��'Y|0
K�Z�����(�d@�Q^u3� T0 k� �<�@? �$1`1	u1�4 �  ��?    � %��  n�f��P��'Y|0
K�Z�����(�d@�Q^u3� T0 k� �<�@? �$1`1	u1�4 �  ��?    � %��  n�f��P��'Y|0
K�Z�����(�d@�Q^u3� T0 k� �8�<? �$1`1	u1�4 �  ��?    � %��  n�e��P��'Y|0
K�Z�����'�d@�Q^u3� T0 k� �4�8? �$1`1	u1�4 �  ��?    � %��  n�e��P��'Y|0
K�Z�����'�d@�Q^v3� T0 k� �0�4? �$1`1	u1�4 �  ��?    � %��  n�e��P��'Y|0
K�Y�����'�e@�R^v3� T0 k� �0�4? �$1`1	u1�4 �  ��?    � %��  n�e��P��'Y|0
K�Y�����'�e@�R^v3� T0 k� �,�0? �$1`1	u1�4 �  ��?    � %��  n�e��P��'Y|0
K�Y�����'�e@�R^v3� T0 k� �(�,? �$1`1	u1�4 �  ��?    � %��  n�d��P��'Y|0
K�Y�����'�e@�R^v3� T0 k� �$�(? �$1`1	u1�4 �  ��?    � %��  n�d��P��'Y|0
K�Y�����'�e@�R^v3� T0 k� �$�(? �$1`1	u1�4 �  ��?    � %��  n�d �P��'Y|0
K�X�����'�e@�R^v3� T0 k� � �$? �$1`1	u1�4 �  ��?    � %��  n�d �P��'Y|0
K�X�����'�e@�R^v3� T0 k� �� ? �$1`1	u1�4 �  ��?    � %��  n�d �P��'Y|0
K�X�����'�e@�R^v3� T0 k� ��? �$1`1	u1�4 �  ��?    � %��  ��d �P��'Y|0
K�X�����'�e@�R^v3� T0 k� ��? �$1`1	u1�4 �  ��?    � %��  ��d �P��'Y|0
K�X�����'�e@�R^v3� T0 k� ��? �$1`1	u1�4 �  ��?    � %��At*^ T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��~��~Q�$1`1	u1�D#�  ��    � -�eAx*^ T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��~��~Q�$1`1	u1�D#�  ��    � -�eAx*^ T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��~��~Q�$1`1	u1�D#�  ��    � -�eAx*^ T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eAx*^ T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA|*^ T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA|)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA|)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA|)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �}��}Q�$1`1	u1�D#�  ��    � -�eA�)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �w}�{}Q�$1`1	u1�D#�  ��    � -�eA�)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �o}�s}Q�$1`1	u1�D#�  ��    � -�eA�)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �k}�o}Q�$1`1	u1�D#�  ��    � -�eA�)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �c}�g}Q�$1`1	u1�D#�  ��    � -�eA�)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �[}�_}Q�$1`1	u1�D#�  ��    � -�eA�)^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �W}�[}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �O}�S}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �K}�O}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �C}�G}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �;}�?}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �7}�;}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �/}�3}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �'}�+}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �#}�'}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �}�}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �}�}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �}�}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �}�}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� �}�}Q�$1`1	u1�D#�  ��    � -�eA�(^T ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� ��}��}Q�$1`1	u1�D#�  ��    � -�eA�'^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� �}��}Q�$1`1	u1�D#�  ��    � -�eA�&^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� �{}�}Q�$1`1	u1�D#�  ��    � -�eA�&^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� �s}�w}Q�$1`1	u1�D#�  ��    � -�eA�&^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� �o}�s}Q�$1`1	u1�D#�  ��    � -�eA�&^U ��  l�Z�,A���\�������(ͼC��,3� T0 k� �g}�k}Q�$1`1	u1�D#�  ��    � -�e  �px \F m c A�p ����x]�FA��^`X"s� T0 k� ��F��F? �$1`1	u1�4 �  ��/   � ��  �px \F m c A�p ����x]�FA��^`X"s� T0 k� ��F��F? �$1`1	u1�4 �  /�/   � ��  �px \F m c A�p ����x]�FA��^`X"s� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  �px�`F m cA�p ����x��FA��^`X"s� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  �px�`F m cA�p ����x��FA��^`X"s� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  �px�`F m cA�p ����w��FA��^`X"s� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  �px�dF m cA�p ����w��FA��^`X"s� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  �px�lF m cA�p ����w�FA��^`X"s� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  =pw�tF Z�D�p���wݼFA��^`X3� T0 k� ��F��F? �$1`1	u1�4 � �/   � ��  =pw�tF Z�D�p���wݼFBN��`X3� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  =lw�tF Z�D�p���v��FBN��`X3� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  =lw�xF Z�D�p���v��FBN��`X3� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  =lv�xF Z�D�p���u��FBN��`W3� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  =hvxF] Z�D�t]���u]�FBN��`W3� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  =hvxF] Z�D�t]���t]�F@�^\W3� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  =huxF] Z�D�t]���t]�F@�^\W3� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  =du|F] Z�D�x]���s]�F@�^\W3� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  Mdu|F] Z�D�x]���s]�F@�^\W3� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  M`t-|F= Z�D�|����r]�F@�^\W3� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  M`t-|F=cD�|����q]�FBN�^\W"�� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  M\s-|F=cD�����p]�FBN�^\W"�� T0 k� ��F��F? �$1`1	u1�4 � ��/   � ��  M\s-|F=cD�����p]�FBN��\W"�� T0 k� � F�F? �$1`1	u1�4 � ��/   � ��  MXr-�F=c D�����o]�FBN��\W"�� T0 k� �F�F? �$1`1	u1�4 � ��/   � ��  MXq-�F=c D�����n]�FBN��\W"�� T0 k� �F�F? �$1`1	u1�4 � ��/   � ��  MTq=�F=c D�����m]�FA���\W"�� T0 k� �F�F? �$1`1	u1�4 � ��/   � ��  MPp=�F=c D�����l]�FA���\W"�� T0 k� �F�F? �$1`1	u1�4 � ��/   � ��  MPo=�F=c D�����k]�FA���\W"�� T0 k� �F�F? �$1`1	u1�4 � ��/   � ��  MLo=�F=c D�����j]�FA���\W"�� T0 k� �F�F? �$1`1	u1�4 � ��/  � ��  ]Hn=�Fmc D�����i]�FA���\W"�� T0 k� � F�$F? �$1`1	u1�4 � ��/   � ��  ]Dm=�Fmc D�����h]�FD>��\W"�� T0 k� �,G�0G? �$1`1	u1�4 � ��*   �  ��  ]Dl=�FmZ� D� ����g]�FD>��\W3� T0 k� �4G�8G? �$1`1	u1�4 � ��*   � !��  ]@k=�FmZ� D��!����f]�FD>��\W3� T0 k� �@F�DF? �$1`1	u1�4 � ��*   � "��  ]<k=�FmZ� D��"����d]�FD>��\W3� T0 k� �HE�LE? �$1`1	u1�4 �  ��*   � #��  ]8j=�F=Z� D��#����c]�FD>��\W3� T0 k� �PE�TE? �$1`1	u1�4 �  ��*   � $��  ]4i=�F=Z� D��$����b]�FD>��\W3� T0 k� �TE�XE? �$1`1	u1�4 �  ��*  � %��  ]0h=�F=Z� D��%����a]�FD>��\W3� T0 k� �HD�LD? �$1`1	u1�4 � �*   � %��  ],g=�F=Z� 	E}�&����_��FE���\W3� T0 k� �@B�DB? �$1`1	u1�4 � ��/   � %��  ](f=�F=Z�$	E}�(���^��FE���\W3� T0 k� �8A�<A? �$1`1	u1�4 � ��/   � %��  ]$e=�FmZ�$	E}�)��
�]��FE���\W3� T0 k� �,@�0@? �$1`1	u1�4 � ��/   � %��  m d=�FmY|$
E}�*��	�[��FE���\W3� T0 k� �$>�(>? �$1`1	u1�4 � ��/   � %��  mc=�FmY|(
E}�+���Z��FE���\W3� T0 k� �=� =? �$1`1	u1�4 � ��/   � %��  mb=�FmY|(
Iݴ,���Y��FF��\W3� T0 k� �<�<? �$1`1	u1�4 � ��/   � %��  ma=�FmY|(
Iݸ-���W��FF��\W3� T0 k� �:�:? �$1`1	u1�4 � ��/   � %��  m`=�FMY|,
Iݸ.	���V��FF��\W3� T0 k� � 9�9? �$1`1	u1�4 � ��/   � %��  m_=�FMY|,
Iݼ/	���V��FF��\W3� T0 k� ��8��8? �$1`1	u1�4 �	 ��/   � %��  m^=�FMY|,
Iݼ0	���V��EF��\W3� T0 k� ��6��6? �$1`1	u1�4 �	 ��/  � %��  m\=�FMY|,
I�1	���U��DF��\W3� T0 k� ��5��5? �$1`1	u1�4 �
 ��/   � %��  m [=�FMY|,
I��2	���T��DF��\W3� T0 k� ��4��4? �$1`1	u1�4 � $�/   � %��  l�Z=�F Y|0
I��3	����T��CE���\W3� T0 k� ��4��4? �$1`1	u1�4 � ��/   � %��  l�Y=�F Y|0
I��3	�� ��S��CE���\W3� T0 k� ��4��4? �$1`1	u1�4 � ��/   � %��  <�X=�F Y|0
I��3	�� ��S��CE���\W3� T0 k� ��4��4? �$1`1	u1�4 � ��/   � %��  <�V=�F Y|0
d��3	�����S��CE���\W3� T0 k� ��4��4? �$1`1	u1�4 � ��/   � %��  <�U=�F Y|0
d��3	�����S��CE���\W3� T0 k� ��5��5? �$1`1	u1�4 �
 ��/   � %��  <�T=�F�Y|0
d��2	�����S��BE���\W3� T0 k� ��5��5? �$1`1	u1�4 �
 ��/   � %��  <�S=�F�Y|0
d��2	�����R��BE���\W3� T0 k� ��5��5? �$1`1	u1�4 �
 ��/   � %��  	��R=�F�Y|0
d��2	�����R��BE���\W3� T0 k� ��5��5? �$1`1	u1�4 �
 ��?   � %��  	��Q=�F�Y|0
d��2	�����R��BE���\W3� T0 k� ��5��5? �$1`1	u1�4 �
 ��?   � %��  	��P=�F�Y|0
d��2	�����R��BE��N\W3� T0 k� ��5��5? �$1`1	u1�4 �	 ��?   � %��  	��O=�F�Y|0
d��2	���}�R��BE��N\W3� T0 k� ��6��6? �$1`1	u1�4 �	 ��?   � %��  	��N=�G�Y|0
d��1���}�Q��BE�� N\W3� T0 k� ��6��6? �$1`1	u1�4 �	 �?    � %��  ��N=�G�Y|0
d��1���}�Q��BE�� N\W3� T0 k� ��6��6? �$1`1	u1�4 � �?    � %��  ��M=�G�Y|0
d��1���}�P��BE��!N\W3� T0 k� ��6��6? �$1`1	u1�4 � ��?    � %��  ��L=�G�Y|0
d��0���}�P��AE��!�\W3� T0 k� ��6��6? �$1`1	u1�4 � ��?    � %��  �K=�G�Y|0
E��0�����O��AE��"�\W3� T0 k� ��7� 7? �$1`1	u1�4 � ��?    � %��  �J=�G�Y|0
E��0�����O��AE��"�\W3� T0 k� ��7� 7? �$1`1	u1�4 � ��?    � %��  \�I=|G�Y|0
E��0�����O��@E��#�\W3� T0 k� � 7�7? �$1`1	u1�4 � ��?    � %��  \�H=|G�Y|0
E��0�����N��@@�#�\W3� T0 k� � 7�7? �$1`1	u1�4 � ��?   � %��  \�G=|G�Y|0
E��0�����N��@@�$�\W3� T0 k� �7�7? �$1`1	u1�4 � ��?    � %��  \�G=|G� Y|0
BM�0�����N��@@�$�\W3� T0 k� �8�8? �$1`1	u1�4 � ��?    � %��  \�F=|G� Y|0
BM�0�����M��@@�$�\W3� T0 k�  9�9? �$1`1	u1�4 � ��U    � %��  \�E=xG�$Y|0
BM�0�����M��@@�%�\W3� T0 k� �:��:? �$1`1	u1�4 � ��U    � %��  \�D=xG�(Y|0
BM�0�����L��@@�%�\W3� T0 k� �;��;? �$1`1	u1�4 � ��U    � %��  \�C=xG�,Y|0
BM�0�����L��@@�&�\W3� T0 k� �;��;? �$1`1	u1�4 � ��U    � %��  \�C=xG�,Y|0
F�0�����L��@@�&�\W3� T0 k� �;��;? �$1`1	u1�4 � ��U    � %��  \�B=xG�0Y|0
F�0�����K��?@�&�XW3� T0 k� � ;�;? �$1`1	u1�4 � ��U    � %��  \�A=xG�4Y|0
F�0�����K��?@�'�XW3� T0 k� � ;�;? �$1`1	u1�4 �  ��U   � %��  \�@=tG�8Y|0
F�0�����K��?@�'�XW3� T0 k� �<�<? �$1`1	u1�4 �  ,�U    � %��  l�@=tG�<Y|0
F�1�����J��?@�(�TW3� T0 k� �<�<? �$1`1	u1�4 �  ��U    � %��  l�?=tG�@Y|0
E��1�����J��?@�(�TW3� T0 k� �<� <? �$1`1	u1�4 � �U    � %��  l�>=tG�DY|0
E��1�����J��?@�(�TW3� T0 k� ,<�0<? �$1`1	u1�4 � ��_    � %��  l�>=tG�HY|0
E��1�����I��?@�)�PW3� T0 k� @<�D<? �$1`1	u1�4 � ��_    � %��  l�==tG�LY|0
E��1�����I��?@�)�LW3� T0 k� T<�X<? �$1`1	u1�4 � ��_    � %��  l�<=tG�LY|0
E��1�����I��>@�*�LW3� T0 k� h<�l<? �$1`1	u1�4 � ��_    � %��  l�<=pG�PY|0
FM�1�����I��>@�*�HW3� T0 k� |<��<? �$1`1	u1�4 � ��_    � %��  l�;=pG�TY|0
FM�1�����H��>@�*�HW3� T0 k� ��=��=? �$1`1	u1�4 � ��_    � %��  l�:=pH�\Y|0
FM�2�����H��>@�+�DW3� T0 k� ��=��=? �$1`1	u1�4 � ��_    � %��  l�:=pH�`Y|0
FM�2�����H��>@�+�@W3� T0 k� ��=��=? �$1`1	u1�4 � ��_    � %��  l�9=pH�dY|0
FM�2�����G��>@�+�@W3� T0 k� ��=��=? �$1`1	u1�4 � ��_    � %��  l|9=pH�hY|0
F]�2�����G��>@�,^<W3� T0 k� ��=��=? �$1`1	u1�4 �	 ��?    � %��  l|8=pHlY|0
F]�2�����G��>@�,^<W3� T0 k� ��=��=? �$1`1	u1�4 �	 ��?    � %��  lx7=lHpY|0
F]�2�����G��=@�,^8W3� T0 k� � =�=? �$1`1	u1�4 �
 ��?    � %��  lx7=lHtY|0
F^ 2�����F��=@�-^4W3� T0 k� �>�>? �$1`1	u1�4 � ��?    � %��  lt6=lHxY|0
F^ 2�����F��=@�-^4W3� T0 k� �(>�,>? �$1`1	u1�4 � ��?    � %��  lt6=lH�Y|0
Fn2�����F��=@�-^0W3� T0 k� �<>�@>? �$1`1	u1�4 � ��?    � %��  lp5=lH�Y|0
Fn3�����F��=@�-^0W3� T0 k� �L>�P>? �$1`1	u1�4 � ��?    � %��  lp5=lH�Y|0
Fn3�����E��=@�.^,W3� T0 k� �`>�d>? �$1`1	u1�4 � ��?    � %��  ll4=lH�Y|0
Fn3�����E��=@�.^,W3� T0 k� �t>�x>? �$1`1	u1�4 � ��?    � %��  ll4=lH� Y|0
Fn3�����E��=@�.^(W3� T0 k� ߈>��>? �$1`1	u1�4 � ��?    � %��  lh3=hH� Y|0
Fn3���� E��=@�/^(W3� T0 k� ߘ?��?? �$1`1	u1�4 � ��?    � %��  lh3=hH��!Y|0
Fn3���� D��<@�/^$W3� T0 k� �?��?? �$1`1	u1�4 � ��?    � %��  lh2=hH��"Y|0
Fn3���� D��<@�/^$W3� T0 k� ��?��?? �$1`1	u1�4 � ��?    � %��  ld2=hH��"Y|0
Fn3���� D��<@�/^ W3� T0 k� ��?��?? �$1`1	u1�4 � ��?    � %��  ld1=hH��#Y|0
Fn3���� D��<@�0^ W3� T0 k� ��?��?? �$1`1	u1�4 � ��?    � %��  l`1=hH��#Y|0
Fn4����D��<@�0^W3� T0 k� ��?��?? �$1`1	u1�4 � ��?    � %��  l`0=hH��$Y|0
Fn4����C��<@�0^W3� T0 k� �?�?? �$1`1	u1�4 � ��?    � %��  l\0=hH��$Y|0
Fn4����C��<@�0^W3� T0 k� � ?�$?? �$1`1	u1�4 � ��?    � %��  l\/=hH��%Y|0
Fn 4����C��<@�1^W3� T0 k� �4@�8@? �$1`1	u1�4 � ��?    � %��  l\/=hH��%Y|0
Fn 4����C��<@�1^W3� T0 k� �H@�L@? �$1`1	u1�4 � ��?    � %��  lX.=dH��&Y|0
Fn 4����C��<@�1^W3� T0 k� �X@�\@? �$1`1	u1�4 � ��?    � %��  lX.=dH��&Y|0
Fn$4����C��<@�1^W3� T0 k�  l@�p@? �$1`1	u1�4 � ��?    � %��  lX.=dH��'Y|0
Fn$4����C��;@�2^W3� T0 k�  �@��@? �$1`1	u1�4 � ��?    � %��  lT-=dH��'Y|0
E�(4����C��;@�2^W3� T0 k�  �@��@? �$1`1	u1�4 � ��?    � %��  lT-=dH��(Y|0
E�(4����C��;@�2^W3� T0 k�  �@��@? �$1`1	u1�4 � ��?    � %��  lP,=dH��(Y|0
E�,4����C��;@�2^W3� T0 k�  �A��A? �$1`1	u1�4 � ��?    � %��  lP,=dH��)Y|0
E�05����C��;@�3^W3� T0 k� ��A��A? �$1`1	u1�4 � ��?    � %��  lP,=dH�)Y|0
E�05����C��;@�3^W3� T0 k� ��A��A? �$1`1	u1�4 � ��?    � %��  lL+=dH )Y|0
E�45����B��;@ 3^W3� T0 k� ��A��A? �$1`1	u1�4 � ��?    � %��  lL+=dH )Y|0
E~86����B��;@ 3^W3� T0 k� �A�A? �$1`1	u1�4 � ��?    � %��  \L*=dH )Y|0
E~<7����B��;@ 3^W3� T0 k� �A�A? �$1`1	u1�4 � ��?    � %��  \H*=`H )Y|0
E~@7����B��;@ 4^W3� T0 k� ,A�0A? �$1`1	u1�4 � ��?    � %��  \H*=`H )Y|0
E~@8����B��;@ 4^ W3� T0 k� @B�DB? �$1`1	u1�4 � ��?    � %��  \H)=`I )Y|0
E~D9����B��;@4^ W3� T0 k� TB�XB? �$1`1	u1�4 � ��?   � %��  \D)=`I *Y|0
D�H:����B��;@4^ W3� T0 k� dB�hB? �$1`1	u1�4 � ��?    � %��  \D)=`I  *Y|0
D�L;����B��;@4]�W3� T0 k� xB�|B? �$1`1	u1�4 � ��?    � %��  �D(=`I $*Y|0
D�P<����B��:@5]�W3� T0 k� ��B��B? �$1`1	u1�4 � ��?    � %��  �D(M`I ,*Y|0
D�P=����B��:@5]�W3� T0 k� ��B��B? �$1`1	u1�4 � ��?    � %��  �@'M`I 0*Y|0
D�T>����A��:@5]�W3� T0 k� ��B��B? �$1`1	u1�4 � ��?    � %��  �@'M`I 4+Y|0
D�X?����A��:@5]�W3� T0 k� ��B��B? �$1`1	u1�4 � ��?    � %��  �@&M`I 8+Y|0
D�\@����A��:@5]�W3� T0 k� ��C��C? �$1`1	u1�4 � ��?    � %��  @&M`I�<+Y|0
D�\A����A��:@5]�W3� T0 k� ��C��C? �$1`1	u1�4 � ��?    � %��  <%M`I�@+Y|0
D�`C����A��:@6]�W3� T0 k� � C�C? �$1`1	u1�4 � ��?    � %��  <$M`I�D+Y|0
D�dD����A��:@6]�W3� T0 k� �C�C? �$1`1	u1�4 � ��?    � %��  <$M`I�H,Y|0
D�hE����A��:@6]�W3� T0 k� �$C�(C? �$1`1	u1�4 � ��?    � %��  <#M\I�P,Y|0
D�hG����A��:@6]�W3� T0 k� �8C�<C? �$1`1	u1�4 � ��?   � %��  �<"\I�T,Y|0
D�lH����A��:@6]�W3� T0 k� �LC�PC? �$1`1	u1�4 � ��?    � %��  �<"\I�X,Y|0
D�lJ����A��:@6]�W3� T0 k� �`D�dD? �$1`1	u1�4 � ��?    � %��  �<!\I�`,Y|0
D�pK����A��:@7]�W3� T0 k� �tD�xD? �$1`1	u1�4 �
 ��?    � %��  �@ \I�d,Y|0
D�tL����@��:@7]�W3� T0 k� ҄D��D? �$1`1	u1�4 �
 ��?    � %��  �@ \I�h-Y|0
I�tM����@��:@7]�W3� T0 k� ҘD��D? �$1`1	u1�4 �	 ��?    � %��  �@\I�p-Y|0
I�xO����@��:@7]�W3� T0 k� �D��D? �$1`1	u1�4 � ��?    � %��  �@\I�t-Y|0
I�xP����@��:@7]�W3� T0 k� ��D��D? �$1`1	u1�4 � ��?    � %��  �D\I�x-Y|0
I�xQ����@��:@7]�W3� T0 k� ��D��D? �$1`1	u1�4 � ��?    � %��  �D\I��-Y|0
I�|R����@��:@8]�W3� T0 k� ��E��E? �$1`1	u1�4 � ��?    � %��  �H�\I��-Y|0
I�|S����@��9@8]�W3� T0 k� ��E��E? �$1`1	u1�4 � ��?    � %��  �H�\I��-Y|0
I�|T����@��9@8]�W3� T0 k� �E�E? �$1`1	u1�4 � ��?    � %��                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��b  ]�,b,b  ����        �  �    ��  �           	    ��      	 ���           `       ���   (
	          d̻          �����     d̻����                      5	 Z��          ְ     ���  H
          P޳         ����     P޳����                    $	 Z��           �     ���   8�

          '�<   � �
      ��eG     '�<��^=       j   	            Z��           �P�    ���   P	B 
          
gm ��	      .�     
gm�                            ����               P  ���    8		 1 	             X(�  � �	   B��g     XQ��ؔ    ���                4 Z���         � �    ���  (	          �ͻ         V�s�;    �ͻ�s�;                        �         
      ��@   8	          '��         j��>~     '����7R    �� l              
   �         �     ��@   	@          eK�         ~���     eC����m     u d               �� �         `     ��@    		�           R"6        ����     R���~�     5 =                ��         	  #p     ��@   P            vU�          ���]�     vM���X�     { F                 �          
 �       ��H   H


           �S ��     � �3q      �S �3q                             ���7              Q  ��@    0)                ��      �                                                                           �                               ��        ���          ��                                                                 �                          5  ��        � Exv     ap F5t    �d�� "              x                j  �   �   �                              ��        � F          G                                                               �                           ����������s�������� ��� E F    
      	       
      �� P1�w       �d �^@ �d _@ �d  b  ��  _� ��  i` �D  h� �� i  �� 0i@ �  i� �D i����X � �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0� ���� � 
�� V  
�| V  
�\ W� 
�| W� 
�| W����� � 
�� W� 
�| W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �������� %�� _  ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"   "D�j�
�� " �
� �  �  
�  1    ��     ��x  �    '    ��     ���       v��  ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �?B      �� � �  ���        � � �  ���        �        ��        �        ��        � 
    ��	     @�����        ��                         I:  �� ��                                    �                ����	            1�w���%��   %�� . F�f $           �TOR 47%) mehlik     0:00                                                                        1  1     �cV � c^ � �c~7 c�/ �c�I c�Q �B�: � B�2 �	C$ �
cj � � cr � �KB2 �KE* � KH1 �KI* �KK' �k�$ �C � �C  � pC$	 �"� � � "� �"� � �*�"�A "�S	�A	
�P*:{9 )�{9 )�{9 )�{) !*K{9 )�{)  *G{9  *A{ � %*P{ � &*F{'*:{) (*G{9  *A{9  *B{9  *B{9  *B{9  *B{3 .*O{C /*K{S )�{51*{] *
{53*{] *
{ � 5*As% 6*Ps= *<sU8*
oU9*6w]  *LOQ;*6wY  *LO=  *F|S *
lD  *DL                                                                                                                                                                                                                         x� P `       �    @ 
        �     ` P E a  ��        
            �������������������������������������� ���������	�
��������                                                                                          ��    ��~�z� ��������������������������������������������������������   �4, :  ��@�@���                                                                                                                                                                                                                                                                                                                                                        � $@aA,�d���)                                                                                                                                                                                                                           �    %    ��  L�J                                   �������������������������������������������������������                                                                                                                                     �    �?                         � ; z           	 	 ���������������������������������������� � � ����������  � ������  �������������� �������� ������ ����� ����������� ������������� ������ ���� ��� �� ��� ������ ������������� �� ����������������������������������������������������������� ����                                 �  
  (    ��	  E�J      �  	                           ������������������������������������������������������                                                                                                                          	                  �    �          �    �w           �     
  
 	     ������������ �� ����� ��������   ��� � ������� ������ ����� �������� ����� ������� ����� ����� ������������� �� ������� �����������  �������������������� ��������� �������������� �� �������� � �������� ������������� ������� �            �                                                                                                                                                                                                                                                                                                    
         �             


           �   }�         wwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwww , J >                                 � t��Z �\                                                                                                                                                                                                                                                                                   	n)n  )n1n        k      a                  m            k                                                                                                                                                                                                                                                                                                                                                                                                                �  � �  � (��  � ��  � ��  � ��  � Z��  ����������������������������������������������u          :   y � :����         �   & AG� �   �   
           	aj�                                                                                                                                                                                                                                                                                                                                   p I H   �      ��        "         !��                                                                                                                                                                                                                        Y   �� �~ ��      �� Z    
���������������������������������������� � � ����������  � ������  �������������� �������� ������ ����� ����������� ������������� ������ ���� ��� �� ��� ������ ������������� �� ����������������������������������������������������������� ���� ������������ �� ����� ��������   ��� � ������� ������ ����� �������� ����� ������� ����� ����� ������������� �� ������� �����������  �������������������� ��������� �������������� �� �������� � �������� ������������� ������� �     �     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    .      6                             4     �  �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$ ^h  ��     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@       �      �     ��    `d �  `b���������� �  � �Q  ��Q          ��   E���� � ��� �� � ��� �$ ^$           �N X�� �) 9        X J��     �    9"  ��  yf  y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  ""   "! " ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                   " ""   "" "!  "" "  """ !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                            " ""   "" !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r` "�"�����   �� �          ����   �       �                                   �    ���  ��                    ��  ��  ���   �       �                        �   ��  ���  � �    �      ��  �   �    �          �         �                                                                                             �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w             ���                         �  ��                    �����                         �     �                                                                                                                                                                                     �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   ��  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �   �   �                .                      ��� ���� ��"  "/�����                            �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .            �  ������� ��                        ���                � ���� ��   � � �                                                                                                                                         �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �   �" �!  �  �� �   �                �  �� Ș ��  ��  �                �   �                               � ����ݼ� ����                                                                                                                                                                               � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �                                                                                                                                                                                                       �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �   �   "   "   "  !�    ��                                    ��  ��  �   �                          �   �   ��� ������ �   �      �       �                        �   ��  ���  � �    �               � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ���� ��� ����                                     	����                                                �   ���                            �   �                                                                                                  �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        T   S   C   3   30  30  ;�  ��  ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ���                   ���                                      ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                     �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   ��  ��  ��  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                                          �   �  �      � �������������               �  �     �   �  �  �                                                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                 ���� ���  ��    �"   "  !�    ��                                 �   �                      �������  ���    �                      �    �                    ��                                                                                                                                                                                                    �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""������������������""""������������������������""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""���������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��������������D�����3333DDDDI����D��DI����3333DDDDADAIA����D������3333DDDD��������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqcV � c^ � �c~7 c�/ �c�I c�Q �B�: � B�2 �	C$ �
cj � � cr � �KB2 �KE* � KH1 �KI* �KK' �k�$ �C � �C  � pC$	 �"� � � "� �"� � �*�"�A "�S	�A	
�P*:{9 )�{9 )�{9 )�{) !*K{9 )�{)  *G{9  *A{ � %*P{ � &*F{'*:{) (*G{9  *A{9  *B{9  *B{9  *B{9  *B{3 .*O{C /*K{S )�{51*{] *
{53*{] *
{ � 5*As% 6*Ps= *<sU8*
oU9*6w]  *LOQ;*6wY  *LO=  *F|S *
lD  *DL3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������$���.�U�[�M��1�O�R�S�U�[�X� � � � � � � � �=��;�������������������������������������������.�G�R�K��2�G�]�K�X�I�N�[�Q� � � � � � �,�>�0�������������������������������������������;�O�I�N�G�X�J��<�S�K�N�R�O�Q� � � � � �,�>�0�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������=��;� ���������������������������������������=��;�	�
�������������������� � � � � � �����������������������������������������%��������������������,�>�0� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                