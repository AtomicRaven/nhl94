GST@�                                                            \     �                                               �   �                        ���������	 ʰ��������������z���        �h      #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    B�j B����
��
�"    B�jl �   B ��
  �                                                                               ����������������������������������       ��    =b? 0Q0 45 118  4             	 

    
               ��� �4 �  ��                 nn 	)
         8:�����������������������������������������������������������������������������������������������������������������������������o  b  o   1  +    '           �                  	  7  V  	                  �  !          := �����������������������������������������������������������������������������                                $`     <  ��   @  #   �   �                                                                                '    	n)n
  !�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    Ld�L��s��������A[�0 _� �˹O��Z3�T0 k� �,&�0&�1�"qe1�t B ��/    ����8Ld �L��w�������A[�0 _� �˺O��Z3�T0 k� �`'�d'�1�"qe1�t B ��/    ����8Ld 
�L��w�������A[�0 c� �˺O��Z3�T0 k� �|(��(�1�"qe1�t B ��/    ����8Lg�
�L��{�������A[�/ c� �ϺO��Z3�T0 k� ��(��(�1�"qe1�t B ��/    ����8Lk�
�L��{�������A[�/ c� �ϺO��Z3�T0 k� ��)��)�1�"qe1�t B ��/    ����8Lk�
�L��{�������A[�/ c� �ϺO��Z3�T0 k� ��)��)�1�"qe1�t B ��/    ����8Lk�
�L���������A[�/ c� �ϺO��Z3�T0 k� ��*��*�1�"qe1�t B ��/    ����8Lk�
�L���������A[�/ c� �ϺO��Z3�T0 k� � *�*�1�"qe1�t B ��/    ����8Lo�
�L���������A[�/ c� �ϺO��Z3�T0 k� �+� +�1�"qe1�t B ��/    ����8Lo�
�L���������A[�/ c� �ӺO��Z3�T0 k� �4+�8+�1�"qe1�t B ��/    ����8Lo�
�L�̃�������A[�/ c� �ӺO��Z3�T0 k� �P,�T,�1�"qe1�t B ��/    ����8Lo�
�L�̃�������A[�/ c� �ӺO��Z3�T0 k� �l,�p,�1�"qe1�t B ��/    ����8Lo�
�L�̃�������A[�/ c� �ӺO��Z3�T0 k� ��-��-�1�"qe1�t B ��/    ����8Lo�
�L�̇�������A[�. c� �ӻO��Z3�T0 k� ��-��-�1�"qe1�t B (�/    ����8Ls�
�L�̇�������A[�. c� �ӻO��Z3�T0 k� Ę.��.�1�"qe1�t B ��/    ����8Ls�
�L�̇�������A[�. c� �׻O��Z3�T0 k� Ĕ.��.�1�"qe1�t B ��/    ����8Ls�
�@̇�������A[�. c� �׻O��Z3�T0 k� Č/��/�1�"qe1�t B ��/    ����8Ls�
�@ ̋�������A[�. g� �׻O��Z3�T0 k� Ą/��/�1�"qe1�t B ��/    ����8Ls�
�@ ̋�=�����A[�. g� �׻O��Z3�T0 k� Ā0��0�1�"qe1�t B ��/    ����8Lw�
�@ ̋�=�����A[�. g� �׻O��Z3�T0 k� �x0�|0�1�"qe1�t B ��/    ����8Lw�
�@ ̋�=�����A[�. g� �׻O��Z3�T0 k� �p1�t1�1�"qe1�t B ��/    ����8Lw�
�@ ̏�=�����A[�. g� �׻O��Z3�T0 k� �l1�p1�1�"qe1�t B ��/    ����8Lw�
�@ ̏�<������A[�. g� �ۻO��Z3�T0 k� �d2�h2�1�"qe1�t B ��/    ����8Lw�
�@$̏�<������A[�. g� �ۻO��Z3�T0 k� �\2�`2�1�"qe1�t B ��/    ����8Lw�
�@$̏�<������A[�. g� �ۻO��Z3�T0 k� �X3�\3�1�"qe1�t B ��/    ����8L{�
�@$̓�<������A[�. g� �ۻO��Z3�T0 k� �P3�T3�1�"qe1�t B ��/    ����8L{�
�@$̓�<������A[�- g� �ۻO��Z3�T0 k� �H4�L4�1�"qe1�t B ��/    ����8L{�
�@$̓�<������A[�- g� �ۻO��Z3�T0 k� �D4�H4�1�"qe1�t B ��/    ����8L{�
�@$̓�<������A[�- g� �ۼO��Z3�T0 k� �<5�@5�1�"qe1�t B ��/   ����8K�{�
�@$̓��������A[�- g� �߼O��Z3�T0 k� �45�85�1�"qe1�t B ��/    ����8K�{�
�@(̗��������A[�- g� �߼O��Z3�T0 k� �06�46�1�"qe1�t B ��/    ����8K�{�
�@(̗��������A[�- g� �߼O��Z3�T0 k� �(6�,6�1�"qe1�t B ��/    ����8K��
�@(̗��������A[�- g� �߼O��Z3�T0 k� � 7�$7�1�"qe1�t B
 ��/    ����8K��
�@(̗��������A[�- g� �߼O��Z3�T0 k� �7� 7�1�"qe1�t B	 ��/    ����8K��
�@(̗��������A[�- g� �߼O��Z3�T0 k� �8�8�1�"qe1�t B ��/    ����8C��
�@(̛��������A[�- g� �߼O��Z3�T0 k� 8�8�1�"qe1�t B ��/    ����8C��
�@(̛��������A[�- k� �߼O��Z3�T0 k� 9�9�1�"qe1�t B ��/    ����8C��
�@,����������A[�- k� �߼O��Z3�T0 k�  9�9�1�"qe1�t B ��/    ����8C��
�@,����������A[�- k� ��O��Z3�T0 k� �:��:�1�"qe1�t B ��/    ����8C��
�@,����������A[�- k� ��O��Z3�T0 k� �:��:�1�"qe1�t B ��/    ����8C��
�@,������"����A[�- k� ��O��Z3�T0 k� ��;��;�1�"qe1�t B ��/    ����8C��
�@,������"����A[�- k� ��O��Z3�T0 k� ��;��;�1�"qe1�t B ��/    ����8C��
�@,������"����A[�- k� ��O��Z3�T0 k� ��;��;�1�"qe1�t B ��/    ����8C�{�
�@,������"����A[�, k� ��O��Z3�T0 k� ��<��<�1�"qe1�t B  ��/    ����8C�{�
�@,������"����A[�, k� ��O��Z3�T0 k� ��<��<�1�"qe1�t B  ,�/    ����8C�{�
�@0������"����A[�, k� ��O��Z3�T0 k� �=��=�1�"qe1�t B  ��/    ����8C�w���@0������"����A[�, k� ��O��Z3�T0 k� �=��=�1�"qe1�t B  ��/    ����8C�w���@0������"����A[�, k� ��O��Z3�T0 k� �>��>�1�"qe1�t B ��/    ����8C�w���@0���L��"����A[�, k� ��O��Z3�T0 k� �>��>�1�"qe1�t B ��/    ����8C�s���@0���L��"����A[�, k� ��O��Z3�T0 k� �?��?�1�"qe1�t B ��/    ����8C�s���@0���L��"����A[�, k� ��O��Z3�T0 k� ��?��?�1�"qe1�t B ��/    ����8C�o���@0���L������A[�, k� ��O��Z3�T0 k� ��@��@�1�"qe1�t B ��/   ����8C�o���@0���L������A[�, k� ��O��Z3�T0 k� ��@��@�1�"qe1�t B ��/    ����8C�k���@0���L������A[�, k� ��O��Z3�T0 k� ��A��A�1�"qe1�t B ��/    ����8C�k���@4���L������A[�, k� ��O��Z3�T0 k� ��A��A�1�"qe1�t B ��/    ����8C�g���@4���L������A[�, k� ��O��Z3�T0 k� ÈB��B�1�"qe1�t B ��/    ����8C�g���@4���L������A[�, k� ��O��Z3�T0 k� ÄB��B�1�"qe1�t B ��/    ����8C�c���@4���L������A[�, k� ��O��Z3�T0 k� �|C��C�1�"qe1�t B ��/    ����8C�_���@4���L������A[�, k� ��O��Z3�T0 k� �tC�xC�1�"qe1�t B ��/    ����8C�_���@4���L������A[�, k� ��O��Z3�T0 k� �pD�tD�1�"qe1�t B ��/    ����8C�[���@4̯� ������A[�, k� ��O��Z3�T0 k� �hD�lD�1�"qe1�t B ��/    ����8C�W���@4̳� ������A[�, o� ��O��Z3�T0 k� �`E�dE�1�"qe1�t B ��/   ����8C�S���@4̳� ��"����A[�, o� ��O��Z3�T0 k� �\E�`E�1�"qe1�t B ��/    ����8C�S���@4̳� ��"����A[�, o� ��O��Z3�T0 k� �TF�XF�1�"qe1�t B ��/    ����8C�O���@4̳� ��"����A[�, o� ��O��Z3�T0 k� �LF�PF�1�"qe1�t B ��/    ����8C�K���@8̷� ��"����A[�, o� ��O��Z3�T0 k� �HG�LG�1�"qe1�t B ��/    ����8C�G���@8̷� ��"����A[�, o� ��O��Z3�T0 k� �@G�DG�1�"qe1�t B ��/    ����8C�C���@8̷� ��"����A[�, o� ��O��Z3�T0 k� �<H�@H�1�"qe1�t B ��/    ����8C�?���@8̷� ��"����A[�+ o� ��O��Z3�T0 k� �4H�8H�1�"qe1�t B ��/    ����8C�;���@8̷� ��"����A[�+ o� ��O��Z3�T0 k� �,I�0I�1�"qe1�t B ��/    ����8C�7���@8̻� ��"����A[�+ o� ��O��Z3�T0 k� �(I�,I�1�"qe1�t B ��/    ����8C�3���@8̻����"����A[�+ o� ��O��Z3�T0 k� � J�$J�1�"qe1�t B ��/    ����8C�/���@8̻����"����A[�+ o� ��O��Z3�T0 k� �J�J�1�"qe1�t B ��/    ����8C�+���@8̻��������A[�+ o� ��O��Z3�T0 k� �J�J�1�"qe1�t B ��/    ����8E�'���@8̻��������A[�+ o� ��O��Z3�T0 k� �K�K�1�"qe1�t B ��/    ����8E�#���@8̻��������A[�+ o� ��O��Z3�T0 k� K�K�1�"qe1�t B ��/    ����8E����@8̿��������A[�+ o� ��O��Z3�T0 k�  L�L�1�"qe1�t B ��/    ����8E����L�<̿��������A[�+ o� ��O��Z3�T0 k� �L��L�1�"qe1�t B ��/    ����8E����L�<̿��������A[�+ o� ��O��Z3�T0 k� �M��M�1�"qe1�t B ��/    ����8E����L�<̿��������A[�+ o� ��O��Z3�T0 k� �M��M�1�"qe1�t B ��/    ����8E����L�<̿��������A[�+ o� ��O��Z3�T0 k� ��N��N�1�"qe1�t B ��/    ����8E����L�<̿��������A[�+ o� ��O��Z3�T0 k� ��N��N�1�"qe1�t B  ��/    ����8E����L�<�×�������A[�+ o� ��O��Z3�T0 k� ��O��O�1�"qe1�t B  ��/    ����8E����L�<�×�������A[�+ o� ��O��Z3�T0 k� ��O��O�1�"qe1�t B  .�/    ����8E����L�<�×�������A[�+ o� ��O��Z3�T0 k� ��P��P�1�"qe1�t B  ��/    ����8E�����L�<�×�������A[�+ o� ��O��Z3�T0 k� �P��P�1�"qe1�t B  ��/    ����8E�����L�<�×�������A[�+ o� ��O��Z3�T0 k� �Q��Q�1�"qe1�t B  ��/    ����8E�����L�<�×�������A[�+ o� ��O��Z3�T0 k� �Q��Q�1�"qe1�t B  ��/    ����8E�����L�<�Ǘ�������A[�+ o� ��O��Z3�T0 k� �R��R�1�"qe1�t B  ��/    ����8E�����L�<�Ǘ�������A[�+ o� ��O��Z3�T0 k� �R��R�1�"qe1�t B  ��/    ����8E�����L�<�Ǘ�������A[�+ o� ��O��Z3�T0 k� ��S��S�1�"qe1�t B ��/    ����8E�����L�<�Ǘ�������A[�+ o� ��O��Z3�T0 k� ��S��S�1�"qe1�t B ��/    ����8E�����L�@�ǘ�������A[�+ o� ��O��Z3�T0 k� ��T��T�1�"qe1�t B ��/    ����8E�����L�@�ǘ�������A[�+ o� ��O��Z3�T0 k� ��T��T�1�"qe1�t B ��/    ����8E�����L�@�ǘ�������A[�+ o� ��O��Z3�T0 k� ��U��U�1�"qe1�t B ��/    ����8C�_�K�C��	��s��7����C��u^���P��Z3�T0 k� ������1�"qe1�t B  ��(    ����CC�_�C�C��	ܬ�{��7����C��u^��� P��Z3�T0 k� �����1�"qe1�t B  ��(    ����BC�|^�;�C��	ܬ���7����C��v^����P��Z3�T0 k� �����1�"qe1�t B  ��(    ����AC�|^�/�C��	ܬ����7����C��v]�����P��Z3�T0 k� �׺�ۺ�1�"qe1�t B  ��(    ����@C�x^��C���	ܬ����7��{�C��w]���P��Z3�T0 k� �Ǹ�˸�1�"qe1�t B  ��(    ����?C�t^��C���	�����7��s�C��x]���P��b��T0 k� ����÷�1�"qe1�t B  ��(    ����>C�p^��C���	�
����7��k�C��x]۰��P��b��T0 k� �������1�"qe1�t B  ��(    ����=C�p^��C���	�
����3��_�C��yMϯ��P��b��T0 k� �������1�"qe1�t B  ��(    ����<C�l^���C���	�	����3��W�C��yMǮ��P��b��T0 k� �������1�"qe1�t B  ��(    ����;C�h^��C���	�	����3��O�C��yM����P��b��T0 k� �������1�"qe1�t B  ��(    ����:C�d^�C���	ܬ	ͯ��3��G�EN�zM����P��b��T0 k� �������1�"qe1�t B  ��(    ����9C�\^ߧC���	ܬͷ��3��7�EN�zM����P{�b��T0 k� �������1�"qe1�t B  �(    ����8C�X^רOM��	ܬͻ��/�	~/�ENxzM���@w�b��T0 k� �������1�"qe1�t B  ��(    ����8C�T^ϨOM��	ܬͿ��/�	~'�ENpzM��w�@o�b��T0 k� �������1�"qe1�t B  ��(    ����8C�P^ǩOM��	��Ù�/�	~�ENdzM��s�@k�b��T0 k� �������1�"qe1�t B  ��(    ����8DL^��OM{�	��Ǚ�/�	~�C�\zM��k�@g�Z3�T0 k� �������1�"qe1�t B  ��(    ����8DD^��OMg�	��˗�/�	~�C�LzM��[��[�Z3�T0 k� �{����1�"qe1�t B  ��(    ����8D@^��OM_�	��ϗ�/�	��C�DzM��S��W�Z3�T0 k� �s��w��1�"qe1�t B  ��(    ����8D8^��OMW�	ܬ�Ӗ�/�	���C�8z=��K��O�Z3�T0 k� �s��w��1�"qe1�t B  ��(    ����8D4^��OMK�	ܬ�Ӗ�/�	���E�0z=��C��K�Z3�T0 k� �s��w��1�"qe1�t B  ��(    ����8D0^��OMC�	ܬ�ו�/�	��E�(z=��;��C�Z3�T0 k� �s��w��1�"qe1�t B  ��(    ����8D(^��OM;�	ܬ�ە�/�	��E� z={�3��?�Z3�T0 k� �o��s��1�"qe1�t B  ��(    ����8D$^{�OM3�	ܬ�۔�/�	}�E�z=s�+��7�Z3�T0 k� �g��k��1�"qe1�t B  ��(    ����8D^s�OM'�L��ߔ�/�	}�E�z=k�#��3�Z3�T0 k� �_��c��1�"qe1�t B  ��(    ����8D^g�OM�L��ߔ�+�	}ߪE�z=g���+�Z3�T0 k� �[��_��1�"qe1�t B  ��(    ����8D^_�OM�L��ߓ�+�	}۪E��z=_���'�bs�T0 k� �W��[��1�"qe1�t B  ��(    ����8D]W�OM�L����+�	}תE��z=W����bs�T0 k� �O��S��1�"qe1�t B  ��(    ����8D]O�OM�L����+�	�ӪC��z=S����bs�T0 k� �G��K��1�"qe1�t B  ��(    ����8D ]G�OL��L����+�	�ϪC��z=K�����bs�T0 k� �C��G��1�"qe1�t B  ��(    ����8D�]�?�OL��L����+�	�˪C��z-C�����bs�T0 k� �?��C��1�"qe1�t B  ��(    ����8D�]�7�OL�L����+�	�ǪC��z-?������bs�T0 k� �;��?��1�"qe1�t B  ��(    ����8D�]�/�OL�L����+�	�êC��z-7������bs�T0 k� �;��?��1�"qe1�t B  ��(    ����8D�]�'�OLߡL����+�	}��C�z-3�������bs�T0 k� �;��?��1�"qe1�t B  ��(    ����8D�]��OLנL����+�	}��C�z-/�������bs�T0 k� �7��;��1�"qe1�t B  ��(    ����8D�]	��OL˞L����+�	}��C�z }#������bs�T0 k� �3��7��1�"qe1�t B  ��(    ����8C��]	��OLÞ�����+�	}��C�z }������Z3�T0 k� �3��7��1�"qe1�t B  ��(    ����8C��]	���C��������+����C�z }������Z3�T0 k� �3��7��1�"qe1�t B  ��(    ����8C�]	���C��������+����C�z }������Z3�T0 k� �3��7��1�"qe1�t B  ��(    ����8C�]	��C��������+����C��z }������Z3�T0 k� �/��3��1�"qe1�t B  ��(    ����8C�]	��C��������+����C�xz }������Z3�T0 k� �+��/��1�"qe1�t B  ��(    ����8C�]	��C���L��ۖ�+����C�lz }������Z3�T0 k� �+��/��1�"qe1�t B  ��(    ����8C��]	�۴E̗�L��ח�+����C�dz }������Z3�T0 k� �'��+��1�"qe1�t B  ��(    ����8C��]	�״Ȅ�L��ә�+����C�\z �������Z3�T0 k� �'��+��1�"qe1�t B  ��(    ����8C��]	�״E��L��Ǜ�+����EMLz ���k����Z3�T0 k� ���#��1�"qe1�t B  ��(    ����8C�x]MӴE�w�ܰ�Ý�+�	}��EM@y ����c����Z3�T0 k� ���#��1�"qe1�t B  ��(    ����8C�p]M˴I|s�ܰ����+�	}��EM8y ����[����Z3�T0 k� �����1�"qe1�t B  ��(    ����8C�h]MǵI|k�ܰ����+�	}�EM0y ����S����Z3�T0 k� �����1�"qe1�t B  ��(    ����8C�`]MõI|g�ܴ����+�	}{�EM(y ����K����Z3�T0 k� �����1�"qe1�t B  ��(    ����8C�X]M��I|_�ܴ����+�	}w�C� x ����C���Z3�T0 k� �����1�"qe1�t B  ��(    ����8C�P]M��I|[�|�����+�	}s�C�x ����;��{�Z3�T0 k� �����1�"qe1�t B  ��(    ����8C�H]M��ELS�|�����+�	�o�C�x ����3��s�Z3�T0 k� �����1�"qe1�t B  ��(    ����8C�4]M��ELG�|� ����+�	�g�C��w ���#��c�Z3�T0 k� �����1�"qe1�t B  ��(    ����8C�,]M��ELC�|��M���+�	�c�EL�v �����[�Z3�T0 k� �����1�"qe1�t B  ��(    ����8C�$]M��EL?�|��M���+�	�_�EL�v �����S�Z3�T0 k� �����1�"qe1�t B  ��(    ����8C�]=��EL;�|��M���+�	}[�EL�u �����O�Z3�T0 k� �����1�"qe1�t B  ��(    ����8C�]=��E<3�|��M���+�	}W�EL�u ��� ���G�Z3�T0 k� �����1�"qe1�t B  ��(    ����8D ]=��E<+�|��M���+�	}O�EL�t ��� ��O7�Z3�T0 k� �����1�"qe1�t B  ��(    ����8D�]=�E<'���M���+�	}K�EL�s ��� ��O/�Z3�T0 k� �����1�"qe1�t B  ��8    ����8D�]={�E<#���M���+��G�EL�s ��� ��O'�Z3�T0 k� �����1�"qe1�t B  ��8    ����8D�]=s�E<���M���+��?�EL�r ��� ��O�Z3�T0 k� �����1�"qe1�t B  ��8    ����8D�]=o�E<���M���+��;�E<�r,����O�Z3�T0 k� �����1�"qe1�t B  ��8    ����8D�]=c�E<�|��M���+��3�E<�p,����O�Z3�T0 k� �����1�"qe1�t B  ��8    ����8D�]=_�E<�|��M���+��+�E<�o-���O�Z3�T0 k� �����1�"qe1�t B  ��8    ����8D�]�[�E<�|��M��+��'�E<�n-���N��Z3�T0 k� �����1�"qe1�t B  ��8    ����8D�]�W�E<�|��M��+��#�E<|n-���N��Z3�T0 k� �����1�"qe1�t B  ��8    ����8D�]�O�E;��|��M{��+���E<tm-���>��Z3�T0 k� �����1�"qe1�t B  ��8    ����8D�]�G�E;��|��Mw��+���E<dk-���>��Z3�T0 k� ���#��1�"qe1�t B  ��8    ����8D�]�C�E+��|��Ms��+���E<\i-���>��Z3�T0 k� �#��'��1�"qe1�t B  ��8    ����8D�]�?�E+�|��Ms��+���E<Th-�{�>��Z3�T0 k� �#��'��1�"qe1�t B  ��8    ����8D�]�?�E+�|��Mo��+����E<Lg-��s�>��Z3�T0 k� �'��+��1�"qe1�t B  �8    ����8Dt]�;�E+�|��Mk�|/���E,@d��c�>��Z3�T0 k� �#��'��1�"qe1�t B ��?    ����8Dl]�;�E+�|��Mg�|/���E,8c��[�>��Z3�T0 k� ���#��1�"qe1�t B ��?    ����8Dd]=;�E+����Mg�|/���E,4b��S�>��Z3�T0 k� �����1�"qe1�t B ��?    ����8D\]=;�E����Mc�|/��߻E,,`��K�N��Z3�T0 k� �����1�"qe1�t B ��?    ����8C�H]=?�E�����_�|/��ӽE, ^�'��7�N��Z3�T0 k� �����1�"qe1�t B ��?    ����8C�@\=C�E�����[�|/��˾E,\�+��/�N��Z3�T0 k� �����1�"qe1�t B ��?    ����8C�8\=C�E�����[�|/��ǿE,[�/��'�N� Z3�T0 k� �����1�"qe1�t B ��?    ����8C�0\=C�@�����W�|/����E,Y�7���N�Z3�T0 k� �����1�"qe1�t B ��?    ����8C�(\=G�@�����S�|/����E,W�;���N|Z3�T0 k� �����1�"qe1�t B ��    ����8C�\=K�@�����O�|/����E,T�G���NpZ3�T0 k� ������1�"qe1�t B	 ��    ����8C�\-K�@�����K�|/����E, S�K����NlZ3�T0 k� ������1�"qe1�t B	 ��    ����8C�\-O�BK�����G�|/����E�Q�O����Nd	Z3�T0 k� �������1�"qe1�t B
 ��    ����8C� \-O�BK�����C�|/����E�O�W����N`
Z3�T0 k� �������1�"qe1�t B
 ��    ����8C��\-S�BK�����C��/�̋�E�N�[����^\Z3�T0 k� �������1�"qe1�t B ��    ����8C��\-S�BK�����?��/�̇�E�L�c����^TZ3�T0 k� �������1�"qe1�t B ��    ����8C��\-W�BK�����;��/���E�K�g����^PZ3�T0 k� �������1�"qe1�t B ��    ����8C��\-[�D������3��/��s�E�H�w����^DZ3�T0 k� �������1�"qe1�t B ��    ����8C��\-_�D������/��/�	|k�E�F�{����>@Z3�T0 k� �������1�"qe1�t B ��    ����8C��\-c�D������+��/�	|g�E�E�����><Z3�T0 k� �������1�"qe1�t B ��    ����8C��\�g�D������'��/�	|_�E�D�����>4Z3�T0 k� ������1�"qe1�t B ��    ����8C��\�k�D���ܿ��#��/�	|[�E�B�����>0Z3�T0 k� ������1�"qe1�t B ��    ����8C��\�o�D���ܿ����/�	|S�E�A�� ��>,Z3�T0 k� ������1�"qe1�t B ��O    ����8C��\�s�D���ܻ����/�	�K�E��>����>$Z3�T0 k� ������1�"qe1�t B ��O    ����8C��\-w�D���ܻ����/�	�G�E��=���>Z3�T0 k� �������1�"qe1�t B ��O    ����8D�\-{�D��ܻ����/�	�?�E��<��w�> Z3�T0 k� �������1�"qe1�t B ��O    ����8D�\-�D��ܻ�M��/�	�;�E��;��
o�>"Z3�T0 k� �������1�"qe1�t B ��O    ����8Dx\-��D��ܻ�M��+�	�7�E��:��g�.#Z3�T0 k� �������1�"qe1�t B ��O    ����8Dh\-��D��ܷ�L���+�	|/�D��8��W�.'Z3�T0 k� �������1�"qe1�t B ��O    ����8D`\-��D��ܷ�L���+�	|+�D��7��O�.)Z3�T0 k� ������1�"qe1�t B ��O    ����8DX\-��D��ܷ�L���+�	|+�D��6��G�. *Z3�T0 k� ������1�"qe1�t B ��O    ����8DL\-��D��ܷ�L���+�	|'�D��6��;�-�,Z3�T0 k� ������1�"qe1�t B ��O    ����8DD\��D��ܷ�L���+�	|#�D��5��3�-�.Z3�T0 k� ������1�"qe1�t B ��O    ����8D<\��D�#�ܷ�<���+�	��D��4��+�-�0Z3�T0 k� ������1�"qe1�t B ��O    ����8D,\� D�+�ܷ�<���+�	��D��3���-�3Z3�T0 k� �������1�"qe1�t B ��O    ����8I�$\�D�/�ܷ�<���'�	��D��3�� �-�5Z3�T0 k� �������1�"qe1�t B ��O    ����8I�\�D�3�ܷ�<���'�	��D� 2��"�-�7Z3�T0 k� �������1�"qe1�t B ��O    ����8I�\�D�7�ܷ�<���'�L�D�2��%	��-�9Z3�T0 k� �������1�"qe1�t B ��O    ����8I�\�D�C�ܷ�<���'�L�D�1��)	����<Z3�T0 k� ̟�����1�"qe1�t B ��O    ����8I� \�
E�G�ܷ�<���'�L�D�1��+	����>Z3�T0 k� ̛�����1�"qe1�t B ��O    ����8I��\�E�K�ܷ�<���'�L�D�1��-	����@Z3�T0 k� ̗�����1�"qe1�t B ��O    ����8I��\�E�S�ܷ�<���#�<�D�1	}�/	����AZ3�T0 k� ̓�����1�"qe1�t B ��O    ����8I��\�E�W�ܷ�<���#�<�D�1	}�2	����CZ3�T0 k� ̓�����1�"qe1�t B ��O    ����8I��\��E�c�L��<���#�<�D�1	~ 6	����FZ3�T0 k� ܋�����1�"qe1�t B
 ��O    ����8I��\��Ig�L��,���#�<�D� 1	~ 8	����HZ3�T0 k� ܋�����1�"qe1�t B
 ��O    ����8I��\��Io�L��,���#�;��D�$1	~9	����JZ3�T0 k� ܇�����1�"qe1�t B	 ��O    ����8I��\�Is�L��,���#���D�(1	�;	����KZ3�T0 k� ܃�����1�"qe1�t B	 ��O    ����8I��\�Iw�L��,���#���D�,2	�=	����MZ3�T0 k� ������1�"qe1�t B ��O    ����8I��\�Iw� ��,������D�82	�=	�����MZ3�T0 k� �{����1�"qe1�t B ��O    ����8I��\� I,w� ��,������D�<2	�>	�����NZ3�T0 k� �w��{��1�"qe1�t B ��O    ����8I��]�(I,w� ��,����;��D�@3�@����OZ3�T0 k� �s��w��1�"qe1�t B ��O    ����8I��]�0I,w� ��,����;��E�D3�@����PZ3�T0 k� �s��w��1�"qe1�t B ��O    ����8I��]�<I,{����,���;��E�P4�B����RZ3�T0 k� �k��o��1�"qe1�t B ��O    ����8I��]�DI{����,���;��E�T5�D����SZ3�T0 k� �g��k��1�"qe1�t B ��O    ����8I��]~LI{����,x ��;��E�\5�E�w���TZ3�T0 k� �g��k��1�"qe1�t B ��O    ����8I��]~TI{����x��;��E�`6�F�o���UZ3�T0 k� �c��g��1�"qe1�t B ��O    ����8I��]~dI{����t��+��E�l7�F�c���WZ3�T0 k� [��_��1�"qe1�t B  ,�O    ����8I��]~h@l{����t��+��E�p8�G�[���XZ3�T0 k� [��_��1�"qe1�t B  ��O    ����8I��]~p@l����t	��+��E�x9�H�S���YZ3�T0 k� W��[��1�"qe1�t B  ��O    ����8I��]~x @l�����t
��+��E��:� H�O���ZZ3�T0 k� S��W��1�"qe1�t B ��O    ����8I��]~| @l�����t��+��E|�:� I�G���[Z3�T0 k� O��S��1�"qe1�t B ��O    ����8I��]~� @l�����p�����E|�<� K�;���\Z3�T0 k� �K��O��1�"qe1�t B ��O    ����8I��]~� @�������t�����E|�=��K�3���]Z3�T0 k� �G��K��1�"qe1�t B ��O    ����8I�|]~� @�������t�����E|�>=�L�+���^Z3�T0 k� �C��G��1�"qe1�t B ��O    ����8I�|]n� @�������t�����E|�@=�L�'���^Z3�T0 k� �C��G��1�"qe1�t B ��O    ����8I�|]n�@�������t�����E|�A=�M����_Z3�T0 k� �?��C��1�"qe1�t B ��O    ����8I�x]n�@���L���t��+��E|�B=�M����_Z3�T0 k� ;��?��1�"qe1�t B ��O    ����8I�t]n�E���M��x��+��E|�E=�N����`Z3�T0 k� 7��;��1�"qe1�t B ��O    ����8I�t]>�E���M��x��+��E|�F=�N����aZ3�T0 k� 3��7��1�"qe1�t B ��O    ����8I�t]>�E���M��|��+��E|�G=�O���aZ3�T0 k� /��3��1�"qe1�t B ��O    ����8I�t]>�E���M��|����E|�I=�O����aZ3�T0 k� �+��/��1�"qe1�t B ��O    ����8I�p]>�E���M��� ���El�J=�O����bZ3�T0 k� �+��/��1�"qe1�t B ��O    ����8I�p]>�Ė�M���!���El�L=�O����bZ3�T0 k� �'��+��1�"qe1�t B ��O    ����8I�p]>�Ė�M���#���El�M=�O����bZ3�T0 k� �#��'��1�"qe1�t B ��O    ����8I�p]>�Ẽ�M��%����El�QM�O���bZ3�T0 k� ���#��1�"qe1�t B ��O    ����8I�p]>�Ẽ�M��'����El�RM�O߾� bZ3�T0 k� �����1�"qe1�t B ��O    ����8I�p]N�E܃�]#��(����El�TM�Oۼ�bZ3�T0 k� �����1�"qe1�t B ��O    ����8I�p]N�E��]'��)����El�VM�N׻�bZ3�T0 k� �����1�"qe1�t B ��O    ����8I�p]N�E��]'��*����El�WM�N׹�bZ3�T0 k� �����1�"qe1�t B ��O    ����8I�p]N�E��]+�	�,���#�El�Y��NӸ�bZ3�T0 k� �����1�"qe1�t B ��O    ����8I�p]N�E�{�]/�	�-���'�El�[��N�Ϸ�bZ3�T0 k� �����1�"qe1�t B ��O    ����8A]p]N�E�w�]/�	�.���/�E\�\�M�˵�bZ3�T0 k� �����1�"qe1�t B ��O    ����8A]p]N�C�s�]7�	�0��7�E\�`�L�ǳ�bZ3�T0 k� �����1�"qe1�t B  ��O    ����8A]p]N�C�o�]7�	�1��?�E\�a�L�Ǳ~aZ3�T0 k� ������1�"qe1�t B  ��O    ����8A]p]N�C�o��;�	,�2��C�E\�c�K�ð~ aZ3�T0 k� ������1�"qe1�t B  ��O    ����8A]p]N�C�k��?�	,�3��G�E\�e��K�ï~$aZ3�T0 k� �������1�"qe1�t B  .�O    ����8Ap]^�C�g��?�	,�4��O�E\�f��J�í~$`Z3�T0 k� �������1�"qe1�t B  ��O    ����8Ap]^�E\c��C�	,�4��W�E\�h��I�ì~(`Z3�T0 k� ������1�"qe1�t B  ��O    ����8Ap]^�E\_��C�	,�5��[�E\�i��I����,_Z3�T0 k� ������1�"qe1�t B  ��O    ����8Ap]^�E\[��G� l�6��c�E\�k��H����0_Z3�T0 k� �����1�"qe1�t B  ��O    ����8Ap]^�E\W��K� l�7��g�E\�l��G����4^Z3�T0 k� �����1�"qe1�t B  ��O    ����8Ap]^�E\S��K� l�7��o�E\�n��F����4^Z3�T0 k� �����1�"qe1�t B  ��O    ����8Ap]^�
ELO��O� l�8���w�EL�o��E�æ�8]Z3�T0 k� �����1�"qe1�t B  ��O    ����8Ap]^�ELC��S���:�����EL�r�|C�ä�<\Z3�T0 k� �ߡ���1�"qe1�t B  ��O 
   ����8Ap]^�EL?��S���;�����EL�s�xB�ã�@[Z3�T0 k� �۠�ߠ�1�"qe1�t B  ��O 
   ����8Ap]^�EL;��W���<�����EL�t�tA�â�DZZ3�T0 k� �۟�ߟ�1�"qe1�t B  ��O 
   ����8Ap]n�E�7��W���=�����C��u�p?�Ǡ�DYZ3�T0 k� �ן�۟�1�"qe1�t B  ��O 
   ����8A]p]n�E�/��W���>�����C��v�l>�ǟ�HXZ3�T0 k� �Ӟ�מ�1�"qe1�t B  ��O 
   ����8A]p]n�E�+��X��?�����C��w�h=�˞�LXZ3�T0 k� �Ӟ�מ�1�"qe1�t B  ��O 
   ����8A]p]n� E�'��X��@�����C��x�d<�˝�LWZ3�T0 k� �ϝ�ӝ�1�"qe1�t B  ��O 
   ����8A]p]n��E���X��A�����C��y�`:�Ϝ�PVZ3�T0 k� �˜�Ϝ�1�"qe1�t B  ��O 
   ����8A]l]n��E���X��B�����C��z�\9�ӛ�TUZ3�T0 k� �ǜ�˜�1�"qe1�t B  ��O 
   ����8C�l]n��E���X
��D��|��C��{�T6�י�XSZ3�T0 k� �Ú�ǚ�1�"qe1�t B  ��O 
   ����8C�l]n��E���X��E��|��EL�|�P4�ۘ�\QZ3�T0 k� ����Ú�1�"qe1�t B  ��O 
   ����8C�h]n��E����X��G��|��EL�|�L2�ߗ�\PZ3�T0 k� ����Ù�1�"qe1�t B  ��O 
   ����8C�h]n��E[���X��H��|��EL�}�H1���`OZ3�T0 k� �������1�"qe1�t B  ��O 
   ����8C�d]n��E[��X��I��|��EL�}�D/���`NZ3�T0 k� ����Ø�1�"qe1�t B  ��" 
   ����8C�`]n��E[��X��L��|��EL�~�<+���dKZ3�T0 k� �������1�"qe1�t B  ��" 
   ����8C�\]n��E[ߢ�X��M��|��EL�~�<*���hJZ3�T0 k� �������1�"qe1�t B  ��" 
   ����8C�\]���E[ס�T��N��}�EL��<*����lIZ3�T0 k� �������1�"qe1�t B  ��" 
   ����8C�X]���E[ϡ�X��P��}�EL��4)����lHZ3�T0 k� �������1�"qe1�t B  ��" 
   ����8C�T]���E[Ǡ�X��Q��}�EL��0)����pFZ3�T0 k� �������1�"qe1�t B  *�" 
   ����8C�P]���E[���X��S��}#�C���$(��xDZ3�T0 k� 럖����1�"qe1�t B  *�" 
   ����8C�L]���E[���X��U��m'�C���'��xBZ3�T0 k� 뛖����1�"qe1�t B  *�" 
   ����8C�L]���E[���X��V��m+�C���'��|AZ3�T0 k� 뗖����1�"qe1�t B  *�" 
   ����8C�H]���E[���X��W��m3�C���&���?Z3�T0 k� 듖����1�"qe1�t B  .�" 	   ����8C�H]���E[���X��X��m7�C���%���>Z3�T0 k� 돖����1�"qe1�t B  ��" 	   ����8C�D]���EK���X��[��mC�C���$�'�ތ;Z3�T0 k� 닕����1�"qe1�t B  ��" 	   ����8D@]���EK���Xܼ\��mG�C����#�/�ސ:Z3�T0 k� ۇ�����1�"qe1�t B  ��" 	   ����8D@]���EK���Xܼ]��mK�C����"�3�ޔ8Z3�T0 k� ۇ�����1�"qe1�t B  ��" 	   ����8D@]���EK���Xܸ^��mO�C��~��!�;�ޘ7Z3�T0 k� ۇ�����1�"qe1�t B  ��" 	   ����8D<]���EK��=X�_��mS�C��~�� �C�ޘ5bs�T0 k� ۇ�����1�"qe1�t B  ��" 	   ����8D<]���EK��=T�`��mS�C��}���G�ޠ4bs�T0 k� ۇ�����1�"qe1�t B  ��" 	   ����8D<]���EK��=T�a��mW�C�x}���O�ޤ2bs�T0 k� �������1�"qe1�t B ��" 	   ����8D<]���E;��=T�b��][�C�t}��S�ި1bs�T0 k� �������1�"qe1�t B  ��" 	   ����8D<]���E;��=P�d"��]_�C�h|��_�ް.bs�T0 k� �������1�"qe1�t B  ��" 	   ����8D<]���E;��=P�e"��]c�C�`{��g�޴,bs�T0 k� �������1�"qe1�t B  ��" 	   ����8D<]���E;��=L�f"��]c�C�\z��o�޸*bs�T0 k� �������1�"qe1�t B  ��" 	   ����8D<]��E;��=L�f"���g�E�Tz��s��)bs�T0 k� �������1�"qe1�t B  ��" 	   ����8D<]��E;��=H�g"���g�E�Ly��{���'bs�T0 k� �������1�"qe1�t B  ��" 	   ����8D<]��E+��=D��h"���k�E�Hx������%bs�T0 k� �������1�"qe1�t B  ��" 	   ����8D<]��E+��=D��h"���k�E�@w������$Z3�T0 k� �������1�"qe1�t B  ��" 	   ����8D<]��E+��M@��i"���o�E�8w������"Z3�T0 k� �������1�"qe1�t B  ��" 	   ����8A�<]��E+��M@��i"���o�E�4v������!Z3�T0 k� �������1�"qe1�t B  ��" 	   ����8A�<]��E+��M<��j"���o�E�,u������Z3�T0 k� �������1�"qe1�t B  ��"    ����8A�<]��@��M8��j���s�E�$t�������Z3�T0 k� �������1�"qe1�t B  ��"    ����8A�<]��@��M4��j���s�E�s�������Z3�T0 k� �ˣ�ϣ�1�"qe1�t B  ��"    ����8A�<]��@��M4��j���s�E�s��	�����Z3�T0 k� �Ӧ�צ�1�"qe1�t B  ��"    ����8A�<]��@��M,�|k���w�C�q���Ä��Z3�T0 k� �ߩ���1�"qe1�t B  ��"    ����8A�<]��E��M(�xk���{�C� p���˄	��Z3�T0 k� �׫�۫�1�"qe1�t B  ��"    ����8A�<]���E��M$�xk���{�C��p���Ӆ	��Z3�T0 k� �Ϭ�Ӭ�1�"qe1�t B  ��"    ����8A�<]���E��M$�tk���{�C��o���ۅ	� b��T0 k� �ϭ�ӭ�1�"qe1�t B  ��"    ����8A�<]���E��] �pk����C��n����	�b��T0 k� �ˮ�Ϯ�1�"qe1�t B  ��"    ����8BM<]���E��]�pj����I��n�� ��	�b��T0 k� �˰�ϰ�1�"qe1�t B  ��"    ����8BM<]���E���]�lj����I��m�����	�b��T0 k� �ϴ�Ӵ�1�"qe1�t B  ��"    ����8BM<]���E���]�hj"�����I��m������
b��T0 k� �ӷ�׷�1�"qe1�t B  ��"    ����8BM<]���E���]�hj"�����I��m�����
b��T0 k� �ӻ�׻�1�"qe1�t B  ��"    ����8BM<]���E���]�di"��]��I��l�����
b��T0 k� �׽�۽�1�"qe1�t B  ��"    ����8B�<]���E�ǯ] �`i"��]��I��l�����
	b��T0 k� �ߺ���1�"qe1�t B  ��"    ����8B�<]���E�˯\��\h"��]��I��k�����	�b��T0 k� �����1�"qe1�t B  ��"    ����8B�@]���E�ϰ\��Xh"��]��I��k����'�	� b��T0 k� �����1�"qe1�t B  �"    ����8B�@]	��E�Ӱ���Xg"��M��I��k ���/�	�$Z3�T0 k� �����1�"qe1�t B  �"    ����8B�@]	��E�ױ���Tg"��M��I��j ���3�	�$Z3�T0 k� �����1�"qe1�t B  ��"    ����8E�D]	��E�۱���Tf"��M��I��i ���;�	�(Z3�T0 k� ������1�"qe1�t B  ��"    ����8E�D]	��E�߲��
�Pe"��M��I��h �� �C�,Z3�T0 k� �������1�"qe1�t B  ��"    ����8E�H]	��E����	�Ld��M��I��g �� �O�0Z3�T0 k� �����1�"qe1�t B  ��"    ����8E�L]	.��E�����Hc�����I��f �� �W�4 Z3�T0 k� �����1�"qe1�t B  ��"    ����8E�P]	.��E�����Hb����I��e �� �[�7�Z3�T0 k� �����1�"qe1�t B  ��"    ����8E�P\	.��E������Da����I��d �� �c�;�Z3�T0 k� �����1�"qe1�t B  ��"    ����8E�T\	.��E������D`����I��d �� �k�O;�Z3�T0 k� �����1�"qe1�t B  ��"    ����8E�X\	.��E�����@`���{�I��c �� �o�O?�Z3�T0 k� �����1�"qe1�t B  ��"    ����8E�X\	��E�����@_���{�I��b �� �w�O?�Z3�T0 k� ���#��1�"qe1�t B  ��"    ����8E�\[	��B\����<^���w�A[�a �� �{�OC�Z3�T0 k� �'��+��1�"qe1�t B  ��"    ����8E�`[	��B\��� �<\���s�A[�` �� ���OG�Z3�T0 k� �+��/��1�"qe1�t B  ��"   ����8E�dZ	��B\�����8[���s�A[�` �� ���OG�Z3�T0 k� �/��3��1�"qe1�t B  ��"    ����8E�dZ	��B\�����8Z���o�A[�_ �� ���OK�Z3�T0 k� �7��;��1�"qe1�t B  ��"    ����8E�hY	.��B\#�����4Y���o�A[�^ �� ���OK�Z3�T0 k� �;��?��1�"qe1�t B  ��"    ����8E�hY	.��B\+�����4X���k�A[�] �� ���OO�Z3�T0 k� �C��G��1�"qe1�t B  ��"    ����8E�lX	.��B\/�����0W���g�A[�\ �� ���OO�Z3�T0 k� �G��K��1�"qe1�t B  ��"    ����8E�pW	.��B\7�����0V���c�A[�\ �� ���OS�Z3�T0 k� �O��S��1�"qe1�t B  ��"    ����8CMpW	.��B\;�����0T���c�A[�[ �� ���OS�Z3�T0 k� �S��W��1�"qe1�t B  ��"    ����8CMtV���B\C�����,S���_�A[�Z �� ���OW�Z3�T0 k� �[��_��1�"qe1�t B  ��"    ����8CMxU���B\G�����,R���[�A[�Y �� ���OW�Z3�T0 k� �_��c��1�"qe1�t B  ��"    ����8CMxT���B\O�����(P���W�A[�X �� ���O[�Z3�T0 k� �g��k��1�"qe1�t B  ��"    ����8CM|S���BlS�����(O���S�A[�X �� ���O[�Z3�T0 k� �o��s��1�"qe1�t B  ��"    ����8CM|R���Bl[�����$N���O�A[�W �� �ÜO_�Z3�T0 k� �s��w��1�"qe1�t B  ��"    ����8CM�QΧ�Blc�����$L���K�A[�V � �ǜO_�Z3�T0 k� �{����1�"qe1�t B  ��"    ����8CM�PΧ�Blg�����$K���G�A[�U � �˝Oc�Z3�T0 k� ������1�"qe1�t B  ��"    ����8CM�OΧ�Blo����� I��MC�A[�U � �ϝOc�Z3�T0 k� �������1�"qe1�t B  ��"    ����8CM�NΧ�Blw����� H��M;�A[�T � �מOc�Z3�T0 k� �������1�"qe1�t B  ��"    ����8CM�MΣ�Bl{����F��M3�A[�S � �۟Og�Z3�T0 k� �������1�"qe1�t B  ��"    ����8CM�Lޣ�Bl���{��E��M'�A[�S � �ߟOg�Z3�T0 k� �������1�"qe1�t B  ��"    ����8C]�Kޣ�Bl���w��C��M�A[�R � ��Ok�Z3�T0 k� �������1�"qe1�t B  ��"    ����8C]�Jޟ�Bl���s��A����A[�Q � ��Ok�Z3�T0 k� �������1�"qe1�t B  ��"    ����8C]�Hޟ�Bl��s�@����A[�Q � ��Oo�Z3�T0 k� �������1�"qe1�t B  ��"    ����8C]�Gޛ�B|��o�>����A[�P � ��Oo�Z3�T0 k� �������1�"qe1�t B  ��"    ����8C]�Fޛ�B|��k�<�����A[�O � ��Oo�Z3�T0 k� �������1�"qe1�t B  ��"   ����8C]�Dޗ�B|��k�;�����A[�O � ���Os�Z3�T0 k� �������1�"qe1�t B  ��"    ����8C]�Cޓ�B|��g�9����A[�N � ���Os�Z3�T0 k� �������1�"qe1�t B  ��"    ����8C]�Aޏ�B|��c�7����A[�N � ���Os�Z3�T0 k� �������1�"qe1�t B  ��"    ����8C]�@B|��c�6����A[�M � ��Ow�Z3�T0 k� �������1�"qe1�t B  ��"    ����8C]�>B|��c�4���۵A[�L � ��Ow�Z3�T0 k� �������1�"qe1�t B  ��"    ����8C]�=B|��_�2���ӷA[�L � ��O{�Z3�T0 k� �������1�"qe1�t B  ��"   ����8Cm�;B|��_�1���˸A[�K � ��O{�Z3�T0 k� �������1�"qe1�t B  ��"    ����8Cm�:��B|���_��/���ǹA[�K � ��O{�Z3�T0 k� �������1�"qe1�t B  ��"   ����8Cm�8�{�B|���[��-�����A[�J � ��O�Z3�T0 k� ������1�"qe1�t B  ��"    ����8Cm�7�w�B����[��,�����A[�J � ��O�Z3�T0 k� �����1�"qe1�t B  ��"    ����8Cm�5�s�B����[��*�����A[�I � ��O�Z3�T0 k� �����1�"qe1�t B  ��"    ����8Kݨ3�o�B����[��(�����A[�I #� ��O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8Kݬ2�g�B���[��&�����A[�H #� �#�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8Kݬ0�c�B��[��%�����A[�H #� �'�O��Z3�T0 k� �#��'��1�"qe1�t B  ��"    ����8Kݬ/�_�B��[��#�����A[�G '� �+�O��Z3�T0 k� �'��+��1�"qe1�t B  ��"    ����8Kݰ.�[�B��W��!��̛�A[�G '� �/�O��Z3�T0 k� �/��3��1�"qe1�t B  ��"    ����8Kݰ,�S�B��W����̛�A[�F '� �/�O��Z3�T0 k� �7��;��1�"qe1�t B  ��"    ����8Kݴ+�O�B�#�S����̗�A[�F '� �3�O��Z3�T0 k� �?��C��1�"qe1�t B  ��"    ����8Kݴ)�G�B�'�S�� ��̓�A[�E +� �7�O��Z3�T0 k� �C��G��1�"qe1�t B  ��"    ����8Kݴ(�C�B�/�S�� ��̏�A[�E +� �;�O��Z3�T0 k� �K��O��1�"qe1�t B  ��"    ����8Kݸ'�;�B]7�S��$��̋�A[�D +� �;�O��Z3�T0 k� �S��W��1�"qe1�t B  ��"    ����8Kݸ%�7�B]?��O��$��̋�A[�D /� �?�O��Z3�T0 k� �[��_��1�"qe1�t B  ��"    ����8Kݸ$�/�B]C��O��(��̇�A[�D /� �C�O��Z3�T0 k� �_��c��1�"qe1�t B  ��"    ����8K�#�+�B]K��O��(��̃�A[�C /� �G�O��Z3�T0 k� �g��k��1�"qe1�t B  ��"    ����8K�!�#�B]S��O��,����A[�C /� �G�O��Z3�T0 k� �l�p�1�"qe1�t B  ��"    ����8K� ��FM[��O��,����A[�B 3� �K�O��Z3�T0 k� �x �| �1�"qe1�t B  ��"    ����8K���FM_��O��0���{�A[�B 3� �O�O��Z3�T0 k� �� �� �1�"qe1�t B  ��"    ����8K���FMg��O��4���w�A[�A 3� �O�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K���FMk��K��4	���w�A[�A 3� �S�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K����FMs��K��8���s�A[�A 7� �W�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K����F={��K��<���o�A[�@ 7� �W�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K���F=��K��<���o�A[�@ 7� �[�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K���F=���K��@���k�A[�@ 7� �_�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K���F=���K��D ���g�A[�? 7� �_�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��۝F=� �G��K����g�A[�? ;� �c�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��םF-��G�|K����c�A[�? ;� �c�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��ϝF-��G�|O����c�A[�> ;� �g�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��ǞF-��G�|S����_�A[�> ;� �g�O��Z3�T0 k� ��	��	�1�"qe1�t B  ��"    ����8K��ÞF-��G�|W����[�A[�> ?� �k�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K����F-��G�|[����[�A[�= ?� �o�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K����F��G�|[����W�A[�= ?� �o�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��-��F��G�|_���W�A[�= ?� �s�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��-��F��C�|c���S�A[�< ?� �s�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��-��F��C�\c���S�A[�< ?� �w�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��-��F��C�\g���O�A[�< C� �w�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��-��F-��C�\k���O�A[�; C� �{�O��Z3�T0 k� �����1�"qe1�t B  ��"   ����8K��-��F-��C�\k���K�A[�; C� �{�O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��-��F-��C�\o���K�A[�; C� ��O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��-��F-��C�\s���G�A[�: C� ��O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��-��F-��C�\w���C�A[�: G� ���O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��{�F=��C�\{���?�A[�: G� ���O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��w�F=��?�\���;�A[�: G� ���O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K��s�F=��?�\����7�A[�9 G� ���O��Z3�T0 k� �����1�"qe1�t B   �"    ����8K� k�F=��C�\����7�A[�9 G� ���O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K�g�F=��C�\����3�A[�9 G� ���O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K�c�FM��C�\����/�A[�9 K� ���O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K�_�FM��C�\����+�A[�8 K� ���O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K�[�FM��C�l����+�A[�8 K� ���O��Z3�T0 k� �����1�"qe1�t B  ��"    ����8K�S�FM��C�l����'�A[�8 K� ���O��Z3�T0 k� ���1�"qe1�t B �"    ����8K��O�FM��C�l����#�A[�8 K� ���O��Z3�T0 k� �,�0�1�"qe1�t B ��/    ����8K��K�F]��G�l�����A[�7 K� ���O��Z3�T0 k� �H�L�1�"qe1�t B ��/    ����8K��G�F]��G�l�����A[�7 K� ���O��Z3�T0 k� �d�h�1�"qe1�t B ��/    ����8K��C�F]��G�l�����A[�7 O� ���O��Z3�T0 k� �|���1�"qe1�t B ��/    ����8K��?�F]��G�l�����A[�7 O� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8K� �;�F]�	�G�l�����A[�6 O� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8K�$�7�Fm�	�G�l�����A[�6 O� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8K�$�3�Fm�	�G�l�����A[�6 O� ���O��Z3�T0 k� �����1�"qe1�t B	 ��/    ����8K�(�/�Fm�	�K�l�����A[�6 O� ���O��Z3�T0 k� ���1�"qe1�t B
 ��/    ����8K�,�+�Fm�	�K�l�����A[�6 O� ���O��Z3�T0 k� �� �1�"qe1�t B ��/    ����8K�,�+�Fm�	�K�l�����A[�5 S� ���O��Z3�T0 k� �8�<�1�"qe1�t B ��/    ����8CN0�'�Fm�	�K�l�����A[�5 S� ���O��Z3�T0 k� �T�X�1�"qe1�t B ��/    ����8CN0�#�Fm�	�K�l�����A[�5 S� ���O��Z3�T0 k� �l�p�1�"qe1�t B ��/    ����8CN4�#�Fm�	�K�l�����A[�5 S� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8CN8��Fm�
�K�l������A[�5 S� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8CN8��Fm�
�K�l������A[�4 S� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8E�<��Fm�
�O�l������A[�4 S� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8E�<��Fm�
�O�l������A[�4 S� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8E�@��Fm�
�O�l������A[�4 W� ���O��Z3�T0 k� ���1�"qe1�t B ��/    ����8E�@��Fm�
�O�l������A[�4 W� ���O��Z3�T0 k� �(�,�1�"qe1�t B ��/    ����8E�D��Fm�
�O�l������A[�4 W� ���O��Z3�T0 k� �D�H�1�"qe1�t B ��/    ����8E�D��Fm�
�O�l������A[�3 W� ���O��Z3�T0 k� �\�`�1�"qe1�t B ��/    ����8E�D��Fm�
�O�l������A[�3 W� ���O��Z3�T0 k� �x�|�1�"qe1�t B ��/    ����8E�H��Fm��O�l������A[�3 W� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8E�H��Fm��O�l߿����A[�3 W� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8E�H��Fm��S�l߾����A[�3 W� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8K�L
��@��S�l�����A[�3 W� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8K�L
��@��S�l�����A[�2 [� ���O��Z3�T0 k� ��� �1�"qe1�t B ��/    ����8K�L	�@��W�l�����A[�2 [� ���O��Z3�T0 k� ���1�"qe1�t B ��/    ����8K�P	�@��W�l�����A[�2 [� ���O��Z3�T0 k� �0�4�1�"qe1�t B ��/    ����8K�P�@��W�l�����A[�2 [� ���O��Z3�T0 k� �L�P�1�"qe1�t B ��/    ����8K�P�@ �[�l�����A[�2 [� ���O��Z3�T0 k� �h�l�1�"qe1�t B ��/    ����8K�T�@ �[�l�����A[�2 [� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8K�T=�@ �_�l�����A[�2 [� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8K�T=�@ �_�l�����A[�1 [� ���O��Z3�T0 k� �����1�"qe1�t B ��/    ����8K�T=�@�c�l�����A[�1 [� ���O��Z3�T0 k� �� �� �1�"qe1�t B ��/    ����8K�X=�@�c�l������A[�1 [� ���O��Z3�T0 k� �� �� �1�"qe1�t B ��/    ����8LX=�L��c�l������A[�1 [� ���O��Z3�T0 k� �!�!�1�"qe1�t B ��/    ����8LXm�L��g�l������A[�1 _� �øO��Z3�T0 k� � !�$!�1�"qe1�t B ��/    ����8LXm�L��g�\������A[�1 _� �ùO��Z3�T0 k� �<"�@"�1�"qe1�t B ��/    ����8L\m�L��k�\������A[�1 _� �ùO��Z3�T0 k� �X"�\"�1�"qe1�t B ��/    ����8L\m�L��k�\������A[�1 _� �ùO��Z3�T0 k� �p#�t#�1�"qe1�t B ��/    ����8L\m�L��k�\������A[�0 _� �ǹO��Z3�T0 k� ��#��#�1�"qe1�t B ��/    ����8L\�L��o�\������A[�0 _� �ǹO��Z3�T0 k� ��$��$�1�"qe1�t B ��/    ����8L`�L��o�\������A[�0 _� �ǹO��Z3�T0 k� ��$��$�1�"qe1�t B ��/    ����8L`�L��o��������A[�0 _� �ǹO��Z3�T0 k� ��%��%�1�"qe1�t B ��/    ����8L`�L��s��������A[�0 _� �ǹO��Z3�T0 k� ��%��%�1�"qe1�t B ��/    ����8L`�L��s��������A[�0 _� �˹O��Z3�T0 k� �&�&�1�"qe1�t B ��/    ����8                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��#� ]�!! � ����  Y Y     ��u:G    ��;��v{�    ���D   
             ���8            ���     ���  @
          ����   � �
     ��BE    �����BE                       _	���8           p�    ���   0	


 
          ��  � � 	    �� �     ����     X �               p ���8�         �P�     ���   8	          ��?b   � �
	   �1�I    ��'%�1��    m                ���8          +P�    ���   @

(         ��B�   � �
     .�?F�    ��B��?F�                       	���8           ؠ�    ���   H

 

         ��]�  ��      B� �Y    ��]�� �Y                            ���8             �  ���    8

 '            ���6    
	   V��
�    �����]    ���^              
 a �         ֐     ��H   0	
           +_         j��?�     +c���?�    ��                  ; �         �     ��@   (
          ��,�         ~�[��    ��1��[�    �� _               �� �          �  �  ��@   8�         ����   [      � <]p    ���� <P}     l �              	 �� j         	 �     ��@   (
          ��ǃ  $ �    ����    �������    �� a                             
 �     ��@   P

B          ����
	      � �     �� �                              ���e                ��@    8		 1                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          U  ��        � ���  T�& �X� <,��u                 x                 j     �   �                          U    ��       � �       T   �           "                                                  �                         �u�B���1�?� �����[ <�� ��� � �   	         
     
      I�� I��       B� �[� �d  a� �� 0g  D� \� �$  b ���< ����J ����X � �d @_  �� 0_� �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ���� ����� ����� ����� � 
�< V� 
� W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����8������ �  ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j B���
��
��"    B�j l �  B �
� �  �  
�      ��     ��s  �        ��     ���      ��    ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �/      ��t �  ���        �# �  ���        �        ��        �        ��        �    \�     6�� �        ��                         �$ ( 	�� �                                    �                 ����             �s���%��  ���8 2               11 Owen Nolan gilny    3:56                                                                        3  3      �)kj_I kr_%cV �=c^	�$�; CBCC �	C � � 
C" � � C# � �C$ � � C& � � C' � �C. � �C4 � �C8 � �B� � �B� � �B� � �c~ � �J� zKE jKK �"�@ � "�R �"�< �*�KH"� �H "�8� �8 
� p!* | �"!� | �#"8 � � $"E � � %"G � �&* | � '"P �(" � )"F �*!� |0+"6 |8 ,"D �P -"C �X ."G �X  "K �P 0"C �X 1"G �X  "K �X  "K �X 4"K �X  "K �X  "K �X  "K �X 8"H �X  "G �X  "G �X ;"K �X  "K �X ="K �X  "K �X  "K �                                                                                                                                                                                                                         �� R         �     @ 
             R P E h  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    � `�� ��������������������������������������������������������   �4, @� * R�� ~� �@.@C��@���G�                                                                                                                                                                                                                                                                                                                                � {@�@��                                                                                                                                                                                                                                     ~  
  2     �  9<�J      �                             ������������������������������������������������������                                                                                                                                        �  � �                      ��                     ����������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� �������������������            �                  �     (    ��   L�J      [�  	                           ������������������������������������������������������                                                                                                                               	     �    _�              �          F @ �             	 	 �������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ����            b                                                                                                                                                                                                                                                           
                              	                   �             


           �   }�                 '�                                              'u  N�                     ������������  R���������������������������������    ��������������������  '}  's����  +�����������������ww�ww333wwwwwwww�ww�ww�ww�ww333wwww 0 I =                                 � �`� �\                                                                                                                                                                                                                                                                                    	n)n
  !�                                      c            m                                                                                                                                                                                                                                                                                                                                                                                                             � ��  � P��  � 2��  � #��  EZm_  �N U��8������������������������������������                      � p           �   & AG� �  �   
              �                                                                                                                                                                                                                                                                                                                                      p G I   �     p                !��                                                                                                                                                                                                                            Y   �� �~ ���      �� ^      ����������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� ��������������������������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ����             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    B   !   2      T                       f     �   �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��     *�X  �  '] >     �f ��     �f �$ ^$ �@      ����� ��   �����    ����� ��   ����� �$ ^$       �  *�                  �������� 
� � ��� �� � ��� �$  � �  �� �  �      �  ��   f�����������J   g��� 	  �     f ^�         �����      f      ��$^�������J���J���� ��      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                          �  �_ <� ���\~~����    UUU�333����~~~~����~~~~����    _�� 3�p �<� �?� �3��|��p��<�                                          �                           �   S  <  <  �  ��  S�<~~~�����~~~����~~~~����~~~~����~~~~����~~~~����~~~~����~~|����3~|3�����~|�<���<~~|;�����~~�3���    �   p  �   �   ��  �p  <�                         _  33?   S�  S�  S�  S�  S�  S�  S�  S3~~~~����~~~~����~~~~��������3333~|5 ��P ~�P ��P ~�P ��P ��P 33P <~| S�� S�~ S�� S�~ S�� S�� S33<~ �����~ �<� |?�~������<~33<�335 33? _      ~~~~����~~~~����  UU                   �        UUUU                            UUP          �                   UUU                            UUU�                            ~~~~                           wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����   �   �   �   ����                                     	�  		  	 � 	 	 	   	   	   	   	  ��                  ��   	   	   	   	   	   	 	 	 � 		  	�                 �   	    �   	    �   	    �   	   	   �  	   �  	   �  	   �                                      
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  "!  " ! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  "!  " ! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  "!    " ""  !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                              
      �  �  ��  �� �� �� 	�� D� EH EZ  DZ 4J 34Z3EH�T��ʄ
����ܩ���� ""�""�""�"/� �� �  ��� ̽� ��� �w� ��� ��� ��� ˻���ܚ��ة��ی����˻ݼˍ�ۻ���Ѕ" �" R�  B      ��  ��  �     �            � �� �   �       �  ��  �  ��  �            �� �̽���ݪ۽w�}�֪�vv���p���          �  ��  �  �  ��  �                    �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                                                                                                                                                                ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .      �   �   �   D   E�  U�  UO                         "  "  "                                                                                                                                                                   �   �   �   ,  ,  ,   *   �  �  �  �  �  �  �  �  �� �� 
B+ 
B" C"  D3  ��  ̘ �� �� +  �"/�"/��� ��  ��  ��    ��  ̽  ��  ��  w}� wz� ��� ��� ��� ��� ̼� ̼� ��� ��� �ۀ ͉� ��@ #4E 34U 3EU 4EU EP D�  ̀ ��� �� �+" �""��"/���� �     �   �  �  �  �   �   �  �                     �   �                       �� �� ��               �  �  �     �   �  �  �                                            � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                  "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��                       "  "  "           �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                        "  .���"    �     �                                                                                                                                                                                                      �� �����ݼڜ��ک��ک��z�	��� 
�� 
�� 	�� ̘ ɪ  ��  �  �� �� ������������ ���  � � � �� �� ������ ��                      �   ��  ��  �̰ ��� ��˰�̻��̻���������ˉ�U��EP�ET �I� ٕ  �D� �L� ��� ��" ����/�"�"�""�����                         /�� �                                         �  ��  �� ��  �� ���                              �������  �                     �  �   �  �  ��  �  ��  �                                                                                                                                                                                                                  �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �     �   �  �  �                   ���� �                                        �  �  �  �   �               �  �� ��  �    � ���                                                                                                                                                                                             	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                � ��                    ���� �                                           �   ���                            �   �                                                                                                    �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �              "      �           �  �   �   ��  �            ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ���                                                                                                                                                                                                               
  �  ̈ �� ,�  ""   "                       �������݅]̻�U�˅U3�U\�BU\�3 "��",�"��"��� ��  �             ݽ���۹����" ��" ��"��".�  �"  �/� .���" � ��              �   .   �   � � �� �� ��                    ��  ��  ���            � ˹ Y�����
�ڛ��٩ �� �̽���ݪ۽w�}�֪�vv���p��� ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ���   ���� �                                           �   ���                            �   �                                                                                                                1    1   "    �   �   �� �����  �    �   �   ,   "   "                   ���ۼ����� 9��C��UTDD�D33��0��  "��
/� � �, �"  �"   �   ˻ڛ��Ȱ��  ��  ��  TJ  EJ  DT  4E  �P  ��  �   /   ��  ��� �                                     � 	�� �� �˙	���
������                Ͱ  ˻  ˻  ۻ  ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                                                                      � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                          �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��                  �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""������������������������""""������ADAIA�A""""�������I�A�A�A""""�����DD�I""""�������DAADAI""""������IDA��""""��������DD��I�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD������������������������3333DDDD�A�AM�M�DM��M334CDDDD�A�AM�M�DDM����3333DDDDDM����DD�����3333DDDDMAM��D�DDM�����3333DDDDDD����M��DM�����3333DDDD������������DD������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(����������������� � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(����������������� 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5���������������� x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x���������������� w w x y�������H���������������������������������H������yxww����������������  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(���������������� , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,���������������� +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+���������������� 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5���������������� =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=����������������     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( ���������������� � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � ����������������� � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � ����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq)kj_I kr_%cV �=c^
�$�; CBCC �	C � � 
C" � � C# � �C$ � � C& � � C' � �C. � �C4 � �C8 � �B� � �B� � �B� � �c~ � �J� zKE jKK �"�@ � "�R �"�< �*�KH"� �H "�8� �8 
� p!* | �"!� | �#"8 � � $"E � � %"G � �&* | � '"P �(" � )"F �*!� |0+"6 |8 ,"D �P -"C �X ."G �X  "K �P 0"C �X 1"G �X  "K �X  "K �X 4"K �X  "K �X  "K �X  "K �X 8"H �X  "G �X  "G �X ;"K �X  "K �X ="K �X  "K �X  "K �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������7�G�Z�Y��<�[�T�J�O�T� � � � � � � � � �:�>�/����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0��������������������������������������������]�K�T��8�U�R�G�T� � � � � � � � � � �:�>�/�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������:�>�/� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�A�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                