GST@�                                                           �o�                                                       ���     �               ����e J���ʲ���������� �������        :i     #    ����                                d8<n    �  ?     �b����  �
fD�
�L���"����D"� j   " B   J  jF�"    "�j* ,  �����
�"     �j@ �    ��
  -                                                                               ����������������������������������      ��    oo b go  4  +c  c  'c       ��       	  
    	G 7� V( 	(                 �n 1         8:8�����������������������������������������������������������������������������������������������������������������������������=?  00  45  18                         
     
                ��  �4  �  ��                  EY            : �����������������������������������������������������������������������������                                �          �   @  &   �   �                                                                                 '      �1n  EY    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��[FK��D���=TO}o���E���lǥA���_������T0 k� �o��s�U8D"!%�0d   ��    ����@��[F[��D���=TL}{���E���lӢA���c������T0 k� ������U8D"!%�0d   ��    ����B��[F[��D���=TJ}���E���lסA���c������T0 k� ������U8D"!%�0d   ��    ����D��[F[��D���MTI}����E���l۟A]��g������T0 k� ,�����U8D"!%�0d   ��    ����F��[F[��D���MTG}����E|��l۝A]��g������T0 k� ,�����U8D"!%�0d   ��    ����H��[F[��D���MTE}����E|��lߜA]��k������T0 k� ,�����U8D"!%�0d  	 ��    ����J��[Fk��D���MTC}����E|��l�A]��k������T0 k� ,�����U8D"!%�0d  	 ��    ����L��[Fk��D���MTB}����E|��l�A]��o������T0 k� ,�����U8D"!%�0d  
 ��    ����N��[Fk��D���MP>m����E|��l�A��s������T0 k� ������U8D"!%�0d  
 ��    ����Q��[Fk��D���MP=m����E|��\�A��w����#�T0 k� ����U8D"!%�0d  
 ��    ����T��[Fk��D���MP;m����El��\�A��{�Ο�#�T0 k� ����U8D"!%�0d   ��    ����W�[Fk��D���ML9m����El��\�A���Ο�#�T0 k� �#��'�U8D"!%�0d   ��    ����Z�[Fk��D���ML7m���#�El��\�A����Ο�#�T0 k� �/��3�U8D"!%�0d   ��    ����]�[Fk��D���]L5m��|#�El��\�CM����Ο�#�T0 k� �?��C�U8D"!%�0d   ��    ����`�[Fk��D���]H3m��|'�El��\�CM����Ο�#�T0 k� �K��O�U8D"!%�0d   ��    ����c�[Fk��D��]D0m��|'�El��\��CM���� n��#�T0 k� -g��k�U8D"!%�0d   ��    ����f [Fk��D��]D.m��|+�D<��\��CM�Η� n��#�T0 k� -s��w�U8D"!%�0d   ��    ����i[Fk��D��]@,m��|+�D<��\��CM�Λ� n��#�T0 k� -�����U8D"!%�0d   ��    ����l[Fk��D��]@*m��|+�D<��\��CM�Σ� n��#�T0 k� -�����U8D"!%�0d   ��    ����o[Fk��D��]<(]��|+�D<��\��CM�Χ� n����T0 k� -�����U8D"!%�0d   ��    ����r�[Fk��D�'�]<&]��|+�D<��\��CM�Ϋ� �����T0 k� =�����U8D"!%�0d   ��    ����u�$[Fk��D�+�]8$]��|/�D<�����CM�γ� �����T0 k� =�����U8D"!%�0d   ��    ����x�,[Fk��D�/�]4"]��|/�D<�����EͰη� �����T0 k� =�����U8D"!%�0d   ��    ����{�<ZFk��D�;�m0���|/�D<�����EͰ��� �����T0 k� =�����U8D"!%�0d   ��    �����@ZB���D�C�m,���|/�D<�����Eͬ��� �����T0 k� ������U8D"!%�0d   ��    ������HZB���D�G�m(���|/�D<�����Eͬ	������T0 k� �����U8D"!%�0d  
 ��    ������PYB���D�K�m$���|/�D<����Eͬ	������T0 k� ����U8D"!%�0d  
 ��    ������XYB���D�S�m$���|/�DL����Eͬ	������T0 k� ����U8D"!%�0d  
 ��    ������`YB���D�W�m ���|/�DL����Eͨ	������T0 k� �'��+�U8D"!%�0d  
 ��    ������hXE���D�[�m���|/�DL����Eͨ	����#�T0 k� �7��;�U8D"!%�0d  	 ��    ������pXE���D�c�m���|/�DL���Eͨ	�� ���#�T0 k� �C��G�U8D"!%�0d  	 ��    �����~xWE���D�g�m���|/�DL����C��	.�� ���#�T0 k� �O��S�U8D"!%�0d   ��    �����~�WE��D�k�m���|/�El����C��	.�� ���#�T0 k� �_��c�U8D"!%�0d   ��    �����~�VE��D�w�m	���|/�El����C��	.�� ���#�T0 k� N{���U8D"!%�0d   ��    �����~�UD��D��m�ӿ|/�El����C��	.�� n��#�T0 k� N�����U8D"!%�0d   ��    �����~�TD��D���]�Ͼ|/�El����E=���� n��#�T0 k� N�����U8D"!%�0d   ��    �����~�SD��D���] �Ͻ|/�El����E=��� n��#�T0 k� N�����U8D"!%�0d   ��    �����~�SD��D���\��ϼ|/�El����E=��� n��#�T0 k� N�����U8D"!%�0d   ��    �������RD��D���\���˺|/�E\����E=��� n��#�T0 k� .�����U8D"!%�0d   ��    �������QD��D���\���˹|/�E\����E=��������T0 k� .�����U8D"!%�0d   ��    �������PD��D���\���Ǹ|/�E\����E=�
�������T0 k� .�����U8D"!%�0d   ��    �������ND�#�D���\��ö|/�E\���#�E=��������T0 k� .�����U8D"!%�0d   ��/    �������ME�'�E���\����|/�I����'�CM��#������T0 k� ?���U8D"!%�0d   ��/    �������KE�+�E���\����|/�I����+�CM��+������T0 k� ?���U8D"!%�0d    ��/    �������JE�3�E���\����|/�I����/�CM��/������T0 k� ?��#�U8D"!%�0d    ��)    �������IE�7�E���\����|/�I����3�CM��3������T0 k� ?#��'�U8D"!%�0d    ,�)    �������GE�?�F��L��}��|/�I����;�E=���?������T0 k� �/��3�U8D"!%�0d    ��)    �������EE�C�F��L��}��|/�I����C�E=��/C������T0 k� �;��?�U8D"!%�0d   ��)    �������DE�K�F��L��}��|/�I����G�E=��/K������T0 k� �G��K�U8D"!%�0d   ��)    ������BE�O�F��L��}��|/�I����K�E=��/O������T0 k� �O��S�U8D"!%�0d   ��)    ������AE�S�F��L��}��|/�I����O�E=��/S������T0 k� �[��_�U8D"!%�0d   ��)    ������@B�[�F��L�����|/�I����S�E=��/[������T0 k� �c��g�U8D"!%�0d   ��)    ������>B�_�F��L�����|/�I����W�E-��/_������T0 k� �g��k�U8D"!%�0d   ��)    �����	�<B�_�F��L�����|/�I����c�E-�� k������T0 k� �{���U8D"!%�0d   ��)    �����	�$:B�_�F��L�����|/�I����g�E-�� s������T0 k� ������U8D"!%�0d   ��)    �����	�(9B�_�F �L�����|/�I����o�E-�� w������T0 k� ������U8D"!%�0d   ��)    �����	�,8B�_�F �<����|/�I����s�E-�� ������T0 k� ������U8D"!%�0d   ��)    �����	�07B�_�F �<����|/�I����w�E-�� �������T0 k� ������U8D"!%�0d   ��)    �����	�46B�_�E��<����|/�I�����E-�� �������T0 k� /�����U8D"!%�0d   ��)    �����	�85B�_�E��<����|/�I������E-�� �������T0 k� /�����U8D"!%�0d   ��)    �����	�<4B�_�E�'�<����|/�I������E-�� �������T0 k� /�����U8D"!%�0d   ��)    �����	�@4B�_�E�/�<��
��|/�A������E-�� �������T0 k� /�����U8D"!%�0d   ��)    �����	�@3B�_�E�7�<��
��|/�A�����E-�� �������T0 k� /�����U8D"!%�0d   �)    ������D2B�_�B�;�<��
�|/�A��-��E�� �������T0 k� ������U8D"!%�0d   �)    ������H1B�_�B�C�<��
{�|/�A��-��E�� ������T0 k� ������U8D"!%�0d   ��)    ������L0B�_�B�S�<��
s�|/�A��-��E��������T0 k� ������U8D"!%�0d   ��)    ������P/@_�B�[�<��
o�|/�A��-��E��������T0 k� ������U8D"!%�0d   ��)    ������T.@_�B�_�<��
k�|/�A��-��E��������T0 k� ������U8D"!%�0d   ��)    ������X.@_�B�g�<��
k�|/�A�{�-��E��������T0 k� ������U8D"!%�0d   ��)   ������X-@c�B�o�<��
g�|/�A�{�-ǠE��������T0 k� /�����U8D"!%�0d    ��)    ������\,@c�B�w� ���
c�|/�BL{�-ˡB������#���T0 k� /�����U8D"!%�0d    ��)    ������`,@c�B�� ��
_�|/�BL{�-ӢB������+���T0 k� /�����U8D"!%�0d    ��)    ������`+@c�B��� ��
[�|/�BL{�-ۣB�������/���T0 k� /� �� U8D"!%�0d    /�)    ������d*@c�B��� ��
W�|/�BL{�ߥB�������7���T0 k� /���U8D"!%�0d    ��)    ������h*@c�B��� ��
S�|/�BL{��B�������?���T0 k� ����U8D"!%�0d    ��)    ������h)@g�B��� ��
S�|/�B�{��B�������C���T0 k� ����U8D"!%�0d    ��)    ������l(@g�B��� ��
O�|/�B�{��B�������K���T0 k� ����U8D"!%�0d    ��)    ������l(@g�E��� ��
K�|/�B����B�������S���T0 k� ����U8D"!%�0d    ��)    ������p'@g�E��� ��
G�|/�B���B������[���T0 k� ����U8D"!%�0d    ��)    ������t'@g�E��� �{�
C�|/�B���B������_���T0 k� ����U8D"!%�0d    ��)    ������t&@g�E��� �{�
C�|/�B���B������g���T0 k� ����U8D"!%�0d    ��)    ������x%@g�E��� �{�
?�|/�B����B������o���T0 k� ��� U8D"!%�0d    ��)    ������x%@g�E��� �{�
;�|/�B�����B�����w���T0 k� � �U8D"!%�0d    ��)    ������|$@k�E��� �w�
7�|/�B����'�B�ÿ�����T0 k� � �U8D"!%�0d    ��)    �������$@k�E��� �w�
7�|/�B����/�B�Ǿ������T0 k� �
�
U8D"!%�0d    ��)    �������#@k�E��� �w�
3�|, B����3�B�˽�����T0 k� ��� U8D"!%�0d    ��)    �������#@k�I�� �w�
/�|, B����;�B�ϼ#�����T0 k� ����U8D"!%�0d    ��)    �������"@k�I�� �w�
/�|, B���C�B�׺ ����T0 k� ����U8D"!%�0d    ��)    �������"@k�I�� �s�
+�|, B���K�B�۹$����T0 k� ����U8D"!%�0d    ��)    �������!@k�I�� �s�
'�|, B���S�B�߸(����T0 k� ����U8D"!%�0d    ��)    �������!@k�I� �s�
'�|, B���[�B���(����T0 k� ����U8D"!%�0d    ��)    ������� @o�E�� �s�
#�|,B���_�B���,_����T0 k� � �U8D"!%�0d    ��)    ������� @o�E�� �s�
#�|,B���g�B���,	_����T0 k� ��U8D"!%�0d    ��)    �������@o�E�� �o�
�|,B���o�B����,
_����T0 k� ��U8D"!%�0d    ��)   �������@o�E�� �o�
�|,B���w�B����0_����T0 k� ��U8D"!%�0d    ��)    �������@o�E�#� �o�
�|,B����B���0_����T0 k� ��U8D"!%�0d    ��)    �������@o�E�+� �o�
�|,B̯����B���0_����T0 k� ��U8D"!%�0d    ��)    �������@o�E�/� �o�
�|,B̷����B���4_����T0 k� ��U8D"!%�0d    ��)    �������@o�E�7� �k�
�|,B̻����B���4_����T0 k� ��U8D"!%�0d    ��)    �������@o�E�;� �k�
�|,B̿����B���4_����T0 k� ��U8D"!%�0d    ��)    �������@o�E�C� �k�
�|,B������B�#��4_����T0 k� ��U8D"!%�0d    ��	    �������@s�@aG� �k�
�|,B���~��B�+��4_����T0 k� ��U8D"!%�0d    ��	    �������@s�@aK� �k�
�|,B���~��B�/��4_����T0 k� ��U8D"!%�0d    ��	    �������@s�@aS� �k�
�|,B���~��B�7�@4_����T0 k� �!�!U8D"!%�0d    ��	    �������@s�@aW� �g�
�|,B���~��B�?�@4_����T0 k� �%�%U8D"!%�0d    ��	    �������@s�@a[� �g�
�|,B���~��B�G�@0o����T0 k� �)�)U8D"!%�0d    ��	    �������@s�@a_� �g�
�|,B���~��B�O�@0 `���T0 k� �,�,U8D"!%�0d    ��	    �������@s�@ag� �g�
��|,B���~��B�S�@0"`���T0 k� �.�.U8D"!%�0d    ��	    �������@s�@ak� �g�
��|,B���~��B�[��0#`���T0 k� �.�.U8D"!%�0d    ��	    �������@s�@ao� �g�
��|,B���~��K�c��,%`���T0 k� �.�.U8D"!%�0d    ��	    �������@s�@as� �g�
��|,B������K�g��,&`���T0 k� � /�/U8D"!%�0d    ��	    �������@s�@a{� �c�
��|,B�����K�o��,(`���T0 k� � /�/U8D"!%�0d    ��	    �������@w�@a|  �c�
��|,B�����K�s��()`���T0 k� ��0� 0U8D"!%�0d    ��	    �������@w�@a�  �c�
��|,B�����K�{��(+`#���T0 k� ��1��1U8D"!%�0d    ��	    �������@w�@a�  �c�
�|,B����K���(,`'���T0 k� ��3��3U8D"!%�0d    ��	    �������@w�@a�  �c�
�|,B����K����(.`+���T0 k� ��4��4U8D"!%�0d    ��	    �������@w�@a�  �c�
�|,B�#���K����$/`/���T0 k� ��6��6U8D"!%�0d    ��	    �������@w�@a� �c�
�|,B�+���K����$1`3���T0 k� ��7��7U8D"!%�0d    ��	    �������@w�@a� �_�
�|,B�3���K����$2`7���T0 k� ��9��9U8D"!%�0d    ��	    �������@w�@a� �_�
�|,B�;�#�K����$3`;���T0 k� ��:��:U8D"!%�0d    ��	    �������@w�@a� �_�
�|,B�C�'�K����$5`?���T0 k� ��;��;U8D"!%�0d    ��	    �������@w�@a� �_�
�|,B�G�+�K���� 6`C���T0 k� ��=��=U8D"!%�0d    ��	    �������@w�@a� �_�
�|,B�O�3�K���� 7`G���T0 k� ��>��>U8D"!%�0d    ��	    �������@w�@a� �_�
�|,B�W�7�K���� 8`K���T0 k� ��?��?U8D"!%�0d    ��	    �������@w�@a� �_�
�|,B�_�;�K���� :`O���T0 k� ��@��@U8D"!%�0d    ��	    �������@{�@a� �_�
�|,B�g�C�K����;`S���T0 k� ��B��BU8D"!%�0d    ��	    �������@{�@a� �[�
ߣ|,B�o�G�K�×�<`W���T0 k� ��C��CU8D"!%�0d    ��	    �������@{�@a� �[�
ߣ|,B�w�K�K�ǖ�=`[���T0 k� ��D��DU8D"!%�0d    ��	    �������@{�@a� �[�
ߣ|,B���S�K�ϖ�>`[���T0 k� ��E��EU8D"!%�0d    ��	    �������@{�@a� �[�
ۣ|,B����W�K�ӕ�@`_���T0 k� ��F��FU8D"!%�0d    ��	    �������@{�@a� �[�
ۣ|,B����[�K�ה�A`c���T0 k� ��G��GU8D"!%�0d    ��	    �������@{�@a� �[�
ۣ|,B����c�K�۔�B`g���T0 k� ��I��IU8D"!%�0d    ��	    �������@{�@a� �[�
ף|,B����g�K�ߓ�C`k���T0 k� ��J��JU8D"!%�0d    ��	    �������@{�@a� �[�
ף|,B����k�K���D`o���T0 k� ��K��KU8D"!%�0d    ��	    �������@{�@a� �[�
ף|,B����s�K���E`o���T0 k� ��K��KU8D"!%�0d    ��	    �������@{�@a� �[�
ӣ|,B����w�K���F`s���T0 k� ��L��LU8D"!%�0d    ��	    �������@{�@a� �W�
ӣ|,B�����K���G`w���T0 k� ��M��MU8D"!%�0d    ��	    �������@{�@a� �W�
ӣ|,B���߃�K����H`{���T0 k� ��N��NU8D"!%�0d    ��	    �������@{�@a� �W�
ӣ|,B������K����I`{���T0 k� ��J��JU8D"!%�0d    �	    �������@{�@a� �W�
ϣ|,B������K����J`���T0 k� ��G��GU8D"!%�0d   ��    �������@{�@a� �W�
ϣ|,B������K���K`����T0 k� ��C��CU8D"!%�0d   ��    �������@�@a� �W�
ϣ|,B������K���L`����T0 k� ��?��?U8D"!%�0d   ��    �������@�@a� �W�
ˢ|,B������K���M`����T0 k� �p;�t;U8D"!%�0d   ��    �������@�@a� �W�
ˢ|,B������K���N`����T0 k� �\8�`8U8D"!%�0d   ��    �������@�@a� �W�
ˢ|,B������K���O`����T0 k� �H4�L4U8D"!%�0d   ��    �������@�@a� �W�
ˢ|,B�����K���P`����T0 k� �00�40U8D"!%�0d   ��    �������@�@a� �W�
Ǣ|,E�����K���PP����T0 k� �-� -U8D"!%�0d   ��    �������@�@a� �W�
Ǣ|,E����K���QP����T0 k� �)�)U8D"!%�0d   ��    �������@�@a� �S�
Ǣ|,E����K�#��RP����T0 k� ��%��%U8D"!%�0d   ��    �������@�@a� �S�
Ǣ|,E�'���K�#��SP����T0 k� ��!��!U8D"!%�0d   ��    �������@�@b  �S�
â|,E�/���K�'��TP����T0 k� ����U8D"!%�0d   ��    �������@�@b  �S�
â|,E�7���K�+��UP����T0 k� ����U8D"!%�0d   ��    �������@�@b �S�
â!�,E�C���K�/��Up����T0 k� ����U8D"!%�0d   ��    �������@�@b �S�
â!�,E�K���K�3��Vp����T0 k� ����U8D"!%�0d   ��    �������@�@b �S�
��!�,E�S���K�7��Wp����T0 k� �p�tU8D"!%�0d   ��    �������@�@b �S�
��!�,E�[���K�;��Xp����T0 k� �\�`U8D"!%�0d  	 ��    �������@�@b �S�
��!�,E�c���K�;��Xp����T0 k� �H�LU8D"!%�0d  	 ��    �������@�@b �S�
��!�,E�k���K�?��Y`����T0 k� �0�4U8D"!%�0d  	 ��    �������@�@b �S�
��!�,E�s�o��K�C��Z`����T0 k� � �  U8D"!%�0d  	 ��    �������@�@b �S�
��!�,E�{�`�K�G��[`����T0 k� ����U8D"!%�0d  
 ��    �������@�@b �S�
��!�,E���`�K�G��[`����T0 k� ������U8D"!%�0d  
 ��    �������@��@b �S�
��!�,E���`�K�K��\`����T0 k� ������U8D"!%�0d  
 ��   �������@��@b �S�
��!�,E���`�K�O��]`����T0 k� ������U8D"!%�0d  
 ��    �������@��@b �O�
��|,E���`�K�S��]`����T0 k� ������U8D"!%�0d  
 ��    �������@��@b  �O�
��|,K���`�K�S��^P����T0 k� ������U8D"!%�0d  
 ��    �������@��@b  �O�
��|,K���`�K�W�P_P����T0 k� ������U8D"!%�0d  
 ��    �������@��@b$ �O�
��|,K���`�B�[�P_P����T0 k� �s��w�U8D"!%�0d  
 ��    �������@��@b$ �O�
��|,K���`#�B�[�P`P����T0 k� �_��c�U8D"!%�0d  
 ��   �������@��@b( �O�
��|,K���`'�B�_�PaP����T0 k� �G��K�U8D"!%�0d  
 ��    �������@��@b( �O�
��|,	K���`'�B�c�PaP����T0 k� �3��7�U8D"!%�0d  
 ��    �������
@��@b( �O�
��|,	K���`+�B�g�PbP����T0 k� ���#�U8D"!%�0d  
 ��    �������
@��@b, �O�
��|,	K���`/�Ek�PbP����T0 k� ����U8D"!%�0d  
 ��    �������
@��@b, �O�
��|,	K���P/�Eo�Pc����T0 k� ������U8D"!%�0d  
 ��    �������
@��@b0 �O�
��|,	K���P3�Es�P d����T0 k� ������U8D"!%�0d  	 ��    �������
@��@b0 �O�
��!�,	K���P3�Ew�P d����T0 k� ������U8D"!%�0d  	 ��    �������
@��@b4 �O�
��!�,	K���P3�E{�P e����T0 k� ������U8D"!%�0d  	 ��    �������
@��@b4 �O�
��!�,	K���P7�E�P e����T0 k� ������U8D"!%�0d  	 ��    �������
@��@b8 �O�
��!�,	K���P7�E��P f����T0 k� ������U8D"!%�0d   ��    �������	@��@b8 �O�
��!�,	K���7�E���P f����T0 k� �s��w�U8D"!%�0d   ��    �������	@��@b8 �O�
��!�,	K���7�E���P g����T0 k� �_��c�U8D"!%�0d   ��    �������	@��@b< �O�
��!�,	K���7�E���P g����T0 k� �G��K�U8D"!%�0d   ��    �������	@��@b< �O�
��!�,	K���7�E���P h����T0 k� �3��7�U8D"!%�0d   ��    �������	@��@b@ �O�
��!�,	K���7�E��� h����T0 k� ���#�U8D"!%�0d   ��    �������	@��@b@ �O�
��!�,	K���7�E��� i����T0 k� ����U8D"!%�0d   ��    �������	@��@b@ �K�
��!�,	K�'��3�E����i����T0 k� �����U8D"!%�0d   ��    �������	@��@bD �K�
��|,	K�+��3�E����j����T0 k� �ߜ��U8D"!%�0d   ��   �������	@��@bD �K�
��|,	K�3��3�E����j����T0 k� �ǘ�˘U8D"!%�0d   ��    �������@��@bD �K�
��|,	K�7��/�E����k����T0 k� ������U8D"!%�0d   ��    �������@��@bH �K�
��|,	K�;��/�E���k ����T0 k� ������U8D"!%�0d   (�    �������@��@bH �K�
��|,
K�C��/�EÆ�l ����T0 k� 럒���U8D"!%�0d   ��    �������@��@bH �K�
��|,
K�G��+�EǇ�l ����T0 k� 룔���U8D"!%�0d   ��    �������@��@bL �K�
��|,
K�K��'�Eˈ�m ����T0 k� 맕���U8D"!%�0d   ��    �������@��@bL �K�
��|,
K�O��'�EӉ/�m ����T0 k� 뫗���U8D"!%�0d   ��    �������@��@bL �K�
��|,
K�W��#�E׉/�m ����T0 k� 믘���U8D"!%�0d   ��    �������@��@bP �K�
��|,
K�[���Eۊ/�n ����T0 k� ۳����U8D"!%�0d    ��    �������@��@bP �K�
��|,
K�_���Eߋ/�n ����T0 k� ۳����U8D"!%�0d    ��    �������@��@bP �K�
��|,
K�c���E�/�o ����T0 k� ۷����U8D"!%�0d    -�    �������@��@bT �K�
��|,
K�g���L_�/�o ����T0 k� ۻ����U8D"!%�0d    ��    �������@��@bT �K�
��|,
K�o�P�L_�/�o ����T0 k� ۿ��àU8D"!%�0d    ��    �������@��@bT �K�
��|,
K�s�P�L_�/�p ����T0 k� �á�ǡU8D"!%�0d    ��    �������@��@bX �K�
��|,
K�w�P�L_�/�p ����T0 k� �ǣ�ˣU8D"!%�0d   ��    �������@��@bX �K�
��|,
K�{�P�L_��q ����T0 k� �Ǥ�ˤU8D"!%�0d   ��    �������@��@bX �K�
��|,
K��P�L_��q ����T0 k� �˦�ϦU8D"!%�0d   ��    �������@��@b\ �K�
��|,
Kσ�P�L_��q ����T0 k� �ϧ�ӧU8D"!%�0d   ��    �������@��@b\ �K�
��|,
Kχ�@�L_��r ����T0 k� ө�שU8D"!%�0d   ��    �������@��@b\ �K�
��|,
Kϋ�@�L_���r ����T0 k� ת�۪U8D"!%�0d   ��    �������@��@b\	 �K�
��|,
KϏ�O��L_���r ����T0 k� ۬�߬U8D"!%�0d   ��    �������@��@b`	 �K�
��|,
Kϗ�O��L_���s ����T0 k� ߯��U8D"!%�0d   ��    �������@��@b`	 �K�
��|,
Kϛ����L_���s ����T0 k� ���U8D"!%�0d   ��    �������@��@b`	 �K�
��|,
Kϟ���L_��_�t ���T0 k� ���U8D"!%�0d   ��    �������@��@bd	 �K�
��|,
Kϣ���Lo��_�t ���T0 k� ���U8D"!%�0d   ��    �������@��@bd	 �K�
��|,
Kϧ���Lo��_�t ���T0 k� ���U8D"!%�0d   ��    �������@��@bd	 �K�
��|,
Kϫ���Lo��_�u ���T0 k� ���U8D"!%�0d   ��    �������@��@bd	 �K�
��|,
Kϯ��Lo��_�u {���T0 k� �����U8D"!%�0d   ��    �������@��@bh	 �K�
��|,
Kϳ�ߡLo��_�u {���T0 k� ������U8D"!%�0d   ��    �������@��@bh	 �K�
��|,
KϷ�ۡL`�_�v {���T0 k� ������U8D"!%�0d    ��    �������@��@bh	 �K�
��|,KϷ�עL`�_�v {���T0 k� �����U8D"!%�0d    ��    �������@��@bh	 �K�
��|,Kϻ�ӢL`�_�v {���T0 k� ����U8D"!%�0d    ��    �������@��@bl	 �G�
��|,K���ӢL`�_�v w���T0 k� ����U8D"!%�0d    ��    �������@��@bl	 �G�
��|,K���ϣL`�_�w w���T0 k� ����U8D"!%�0d    /�    �������@��@bl	 �G�
��|,K���ˣL`�_�w w���T0 k� ����U8D"!%�0d    ��    ������ @��@bl	 �G�
��|,K�˿ǣL`�_�w w���T0 k� ����U8D"!%�0d    ��    ������ @��@bl	 �G�
��|,K�˿äL`�_�w w���T0 k� ����U8D"!%�0d    ��    ������ @��@bp	 �G�
��|,K�ϿäL`�_�x w���T0 k� ����U8D"!%�0d    ��    ������ @��@bp	 �G�
��|,B�ӿ��L`�_�x s���T0 k� ����U8D"!%�0d    ��    ������ @��@bp	 �G�
��|,B�׿��L`�_�x s���T0 k� ����U8D"!%�0d    ��    ������ @��@bp	 �G�
��|,B�ۿ/��L`�_�y s���T0 k� ���#�U8D"!%�0d    ��    ������ @��@bp	 �G�
��|,B�ۿ/��L`�_�y s���T0 k� �#��'�U8D"!%�0d    ��    ������ @��@bt	 �G�
��|,B�߾/��L`�_�ys���T0 k� �'��+�U8D"!%�0d    ��   ������ @��@bt
 �G�
��|,B��/��L`�_�ys���T0 k� �'��+�U8D"!%�0d    ��    ������ @��@bt
 �G�
��|,E��/��L`�_�zo���T0 k� �+��/�U8D"!%�0d    ��    ������ @��@bt
 �G�
��|,E��/��L`�_�zo���T0 k� �/��3�U8D"!%�0d    ��   ������ @��@bt
 �G�
��|,E��/��L`�_�zo���T0 k� �3��7�U8D"!%�0d    ��    ������ @��@bx
 �G�
��|,E��/��L`�_�zo���T0 k� �7��;�U8D"!%�0d    $�    ������ @��@bx
 �G�
��|,E���/��L`�_�z�o���T0 k� �3��7�U8D"!%�0d    ��    ������ @��@bx
 �G�
��|,E���/��L`�_�{�k���T0 k� �3��7�U8D"!%�0d    ��    ������ @��@bx
 �G�
��|,E���/��L`�_�{�k���T0 k� �3��7�U8D"!%�0d    ��    ������@��@bx
 �G�
��|,E��/��L`�_�{�k���T0 k� �3��7�U8D"!%�0d    ��    ������@��@bx
 �G�
��|,E��/��L`�_�{�g���T0 k� �/��3�U8D"!%�0d    ��    ������@��@b|
 �G�
��|,E��/��L`�_�|�g���T0 k� �/��3�U8D"!%�0d    ��    ������@��@b|
 �G�
��|,E��/��L`�_�|�c���T0 k� �/��3�U8D"!%�0d    ��    ������@��@b|
 �G�
��|,E��/��L`�_�|�c���T0 k� �/��3�U8D"!%�0d    ��    ������@��@b|
 �G�
��|,E��/��L`�_�|�_���T0 k� �+��/�U8D"!%�0d    ��    ������@��@b|
 �G�
��|,E��/��L`�_�|�_���T0 k� �+��/�U8D"!%�0d    ��    ������@��@b|
 �G�
��|,E�#�/��L`�_�}�[���T0 k� �+��/�U8D"!%�0d    ��    ������@��@b|
 �G�
��|,E�#�/��L`�_�}�[���T0 k� �'��+�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E�#�/��L`�_�}�[���T0 k� �'��+�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E�#�/��L`�_�}�W���T0 k� �'��+�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E�#�/��L`�_�}�W���T0 k� �'��+�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/�L`�_�}�W���T0 k� �#��'�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/�L`�_�~�W���T0 k� �#��'�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/{�LP�_�~W���T0 k� �#��'�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/{�LP�_�~S���T0 k� �#��'�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/w�LP�_�~S���T0 k� ���#�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/w�LP�_�~S���T0 k� ���#�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/s�LP�_�~S���T0 k� ���#�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/s�LP�_�S���T0 k� ���#�U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/o�A��_�O���T0 k� ����U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/o�A��_�O���T0 k� ����U8D"!%�0d    ��    ������@��@b�
 �G�
��|,E��/k�A��_�O���T0 k� ����U8D"!%�0d    ��    ������@��@b�
 �G�
��|,C��/k�A��_�O���T0 k� ����U8D"!%�0d    ��    ������@��@b�
 �G�
��|,C��/g�A�#�_�O���T0 k� ����U8D"!%�0d    ��    ������@��@b�
 �G�
��|,C��/g�A�#�_�� O���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C��/g�A�#�_� K���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C��/c�A�#�_� K���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C��/c�A�#�_� K���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C���/_�A�#�_� K���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C���_�A�#�_�~ K���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C���_�D0�_�~ K���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C��[�D0�_�~ K���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C��[�D0�_�~ G���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C��[�D0�_�} G���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C��W�D0�_�} G���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C�ߦ�W�D0�_�} G���T0 k� ����U8D"!%�0d    ��   ������@��@b� �G�
��|,C�ۦ�S�D0�_�} G���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C�צ�S�D0�_�} G�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,C�ӥ�O�D0�_�| G�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,Lϥ�O�D0�_�| G�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,Lˤ�K�D0�_�| C�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,LǤ�G�D0�_�| C�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,Lã�G�D@�_�| C�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,L���C�D@�_�{ C�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,L���?�D@�_�{ C�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,L���;�D@�_�{ C�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,L���7�D@�_�{ C�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,L���3�D@�_�{ C�##�T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,L���/�D@�_�z C���T0 k� ����U8D"!%�0d    ��    ������@��@b� �G�
��|,L���+�DO��_�z ?���T0 k� �����U8D"!%�0d    ��    ������@��@b� �G�
��|,L/���'�DO��_�z ?���T0 k� �����U8D"!%�0d    ��    ������@��@b� �G�
��|,L/���#�DO��_�z ?���T0 k� �����U8D"!%�0d    ��    ������@��@b� �G�
��|,L/����DO��_�z ?���T0 k� �����U8D"!%�0d    ��    ������@��@b� �G�
��|,L/����E_�_�z ?���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/����E_�_�y ?���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/����E_�_�y ?���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/����E_�_�y ?���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/����E_�_�y ?���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/����E_ߒ_�y ?���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/�����E_ۓ_�y ;�#�T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/�����E_ד_�y ;�#�T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/���E_Ӕ_�x ;�#�T0 k� ������U8D"!%�0d    ��   ������@��@b� �G�
��|,L/{���E_˔_�x ;�#�T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/w���C�Ǖ_�x ;�#�T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/w���C�Ö_�x ;�#�T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/s��߭Cￖ_�x;�#�T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/o��۬Cﻗ_�x;�#�T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/k��׫C﷗_�x;�#�T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/k��ӫI���_�w;�#�T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/g��ϪI���_�w;�#�T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/c�˩I���_�w;���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/c�ǨI���_�w�7���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/_�çI���_�w�7���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/_���I���_�w�7���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/[���I���_�w�7���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/W���I���_�w�3���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/W���I���_�w�3���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/S���I���_�v�3���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/S���I���_�v�/���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/O����I���_�v�+���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/K����I���_�v�+���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/K����I���_�v�'���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/G����I���_�v�'���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/G����I���_�v�#���T0 k� ������U8D"!%�0d    ��   ������@��@b� �G�
��|,L/C����I���_�v����T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/C����I���_�v����T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/?����I���_�v����T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/?����I���_�u����T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/;����I���_�u����T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/;����I����u����T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/7����I����uP���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L7����I����uP���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L3����I����u_����T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L3����A_���u_����T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/����A_���u_����T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L/����A_���u_���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,L+����A_���u_���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,C�+����A_���u_���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,C�'����L���uO���T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,C�'����L��/�tOۏ��T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,C�#����L��/�tO׎��T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,C�����L��/�tOϏ��T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,E���ÎL��/�tOˏ��T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,E���ÍL��/�tOǏ��T0 k� ������U8D"!%�0d    ��    ������@��@b� �G�
��|,E���ǍL��/�tO����T0 k� �Ͽ�ӿU8D"!%�0d    ��    ������@��@b� �G�
��|,E���ˍL��/�tO����T0 k� �Ͽ�ӿU8D"!%�0d    ��    ������@��@b� �G�
��|,E���όL��/�tO����T0 k� �Ͽ�ӿU8D"!%�0d    ��    ������@��@b� �G�
��|,E���ӌL��/�tO����T0 k� �Ͽ�ӿU8D"!%�0d    ��    ������@��@b� �G�
��|,E���ӌL/���tO����T0 k� �Ͽ�ӿU8D"!%�0d    ��    ������@��@b� �G�
��|,E���׋L/���tO����T0 k� �˿�ϿU8D"!%�0d    ��    �����,\C�'�E]L3k��L� �Dg�� JI�D
�_��xZ��T0 k� ��8��8U8D"!%�0d    ��    � 4�8,XC�#�E]@6k��L� �E]_��GI�D�_��xZ��T0 k� ��5��5U8D"!%�0d    ��    � 4�8,TC��E]<7{��L� �E][��EI�D�_��xZ��T0 k� ��3��3U8D"!%�0d    ��    � 4�8,PC��E]<7{��L� �E]W��EI�D�_��xZ��T0 k� ��2��2U8D"!%�0d    �    � 4�8,LC��E]87{��L��E]K��CI�D�_��xZ��T0 k� ��1��1U8D"!%�0d    ��    � 4�8,L C��E]87{��L��E]G��CI�D�_��xZ��T0 k� ��1��1U8D"!%�0d    ��    � 4�8,H!C��E]47{��L��E]?�� BFD�_��xZ��T0 k� ��/��/U8D"!%�0d    ��    � 4�8,H"C��E]47{��<��E];���AFD�_��xY��T0 k� ��-��-U8D"!%�0d    ��    � 4�8,H$E>�E]07{��<��EM3���AFD�_��xY��T0 k� ��+��+U8D"!%�0d    ��    � 4�8D&E=��E]07{�<��EM'���?FH�_��xY��T0 k� ��)��)U8D"!%�0d    ��    � 4�8D'E=��E]07;�<��EM#���>FH�_��xX��T0 k� ��(��(U8D"!%�0d    ��    � 4�8D(E=��E],7;��x�EM���=FH �_��xX��T0 k� ��'��'U8D"!%�0d    ��    � 4�8D)E=��E],7;�
�t�EM���<FL!�_��xW��T0 k� ��&��&U8D"!%�0d    ��    � 4�8D+E=��E],7;��l�EM���:FL%�_��xV��T0 k� ��#��#U8D"!%�0d    ��    � 4�8D,E=��A,7;��h�EM���9FP&�[��xU��T0 k� ��"��"U8D"!%�0d    ��    � 4�8D-E=��A,7;�L`�EL����8FP(�[��xT��T0 k� ��!��!U8D"!%�0d    ��    � 4�8D.CM��A(7;�L\�EL����6FP)�[��xT��T0 k� �� �� U8D"!%�0d    ��    � 4�8H0CM��A(6;�LT	�EL����4E�P)�[��xR��T0 k� ����U8D"!%�0d    ��    � 4�8�L1CM��EM$6;�LL
�EL����2E�T*�[��xQ��T0 k� ����U8D"!%�0d    ��    � 4�8�T2CM��EM$6;�LH
�E<���1E�X+�[��xP��T0 k� ����U8D"!%�0d    ��    � 4�8�\3E�׾EM 6+�<H
�E<���0E�X,�[��xO��T0 k� ����U8D"!%�0d    ��    � 4�8�l4E�ϻEM5+�$<H
�E<���-E�`.	�[��xM��T0 k� ����U8D"!%�0d    ��    � 4�8�l4E�˹E=5+�&<H
�E<���+E�`/	�[��xL��T0 k� ����U8D"!%�0d    ��    � 4�8p5E�ǷE=5+�(<D�CL��\�)E�d0	�[��xK��T0 k� ����U8D"!%�0d    ��    � 4�8t6E�õE=4+�*<D�CL��\�(E�h1	�[��xI��T0 k� ����U8D"!%�0d    ��    � 4�8|8Eͻ�E=3+�.<D�CL��\�$E�p3	�[��xG��T0 k� ����U8D"!%�0d    ��G    � 4�8�9Eͷ�B�3+�0<@�CL��\�"E�t4	�[��xE��T0 k� ����U8D"!%�0d    ��G    � 4�8�:Eͳ�B�2+�3<@�CL��\�!E�x5	�[��xD��T0 k� ����U8D"!%�0d    ��G    � 4�8�:Eͯ�B�1+�5,@�CL��\�E�|6	�[��xC��T0 k� ����U8D"!%�0d    ��G    � 4�8�<Eͣ�B�0+�9,<|CL���E��8	�[��x@��T0 k� ��	��	U8D"!%�0d    ��G    � 4�8�=E͟�B�0+�;,<|CL��E��8	�[��x>��T0 k� ����U8D"!%�0d    ��G    � 4�8�>E͛�B�/+�=,<|CL{��E��9	�[��x<��T0 k� ����U8D"!%�0d    ��G    � 4�8�>E͓�B�.+�?,@|CLw��E��:	�[��x;��T0 k� ����U8D"!%�0d    ��G    � 4�8�?E͏�B�-+�B@| C\o��E��:	�[��x9��T0 k� ����U8D"!%�0d    ��G 	   � 4�8�AE̓�B�,+�F@| C\g��E��;	�[��x6��T0 k� ������U8D"!%�0d    ��G 	   � 4�8�BE��B�+�HD|C\_���E��<	�[��x4��T0 k� ������U8D"!%�0d    ��G 	   � 4�8�BE�w�C*�JD|C\[���E��<	�[��x2��T0 k� ������U8D"!%�0d    ��G 	   � 4�8�CE�s�C)�LD|C\W���E��=	�[��x0��T0 k� ������U8D"!%�0d    ��G 	   � 4�8�DE�o�C(�NH|E�O���E��=	�[��x.��T0 k� ������U8D"!%�0d    ��G 	   � 3�8�EE�_�C'�RL|E�G���E��=	�[��x+��T0 k� ������U8D"!%�0d    ��G 	   � 2�8�FE�[�C&�TL|E�?�	�E��>	�[��x)��T0 k� ������U8D"!%�0d    ��G 	   � 1�8�FE�S�C%�VP|E�;�	�E��>	�[��x'��T0 k� ������U8D"!%�0d    ��G 	   � 0�8�GE�O�C$�XP|E�3�	�E��>	�[��x%��T0 k� ������U8D"!%�0d    ��G 	   � /�8�HE�G�C#�ZT|E�/�	�E��>	�[��x#��T0 k� ������U8D"!%�0d    ��G 	   � .�8�HE�?�C!��\T|E�'�	� E��>	�[��x!��T0 k� ������U8D"!%�0d    ��G 
   � -�8��JE�3�C ��_X|E��	��E��=	�[��x��T0 k� ������U8D"!%�0d    ��G 
   � ,�8��JE�+�C ��a,\|
C��	��E��=	�[�	�x��T0 k� ������U8D"!%�0d    ��G 
   � +�8��KE�'�C$��c,\|	C��	��E��=	�[�	�x��T0 k� ������U8D"!%�0d    ��G 
   � *�8��LE��C$�e,`|C��	��E��<	�[�	�x��T0 k� ������U8D"!%�0d    ��G 
   � )�8��ME��C(�h,d|C�����E��<	�[�	�x��T0 k� ������U8D"!%�0d    ��G 
   � (�8��ME��C,�j,d| E;�����E��;	�[�	�x��T0 k� ������U8D"!%�0d    ��G 
   � '�8��NE���C0�l,d| E;�����C��;	�[�	�x��T0 k� ������U8D"!%�0d    ��G 
   � &�8��OE���C0�m,h|  E;�����C��:	�[�	�x��T0 k� ������U8D"!%�0d    ��G 
   � %�8� OE��C4�o,h|'�E;�����C� :	�[�	�x��T0 k� ������U8D"!%�0d    ��G 
   � $�8�PE��E-8�rl�'�E;����C�9N[�	�x��T0 k� ������U8D"!%�0d    ��G 
   � #�8�QE�ۆE-<�sl�'�E;����E�8N[�	�x��T0 k� ������U8D"!%�0d    ��G 
   � "�8�RE�ӆE-@� up�+�E;����E�8N[�	�x
��T0 k� ������U8D"!%�0d   �G 
   �  �8	=RE�ˇE-D�vp�+�E;����E�7N[�	�x	��T0 k� �����U8D"!%�0d   ��O 
   � �8	=$SE���E-L�y�t�+�E+��ܓ�E�6N[�	�x��T0 k� �_��c�U8D"!%�0d   ��O 
   � �8	=(SE���E-L
�z�x�+�E+��ܓ�E�5 [�	�x��T0 k� �O��S�U8D"!%�0d   ��O 
   � �8	=,TE���E-P� |�x�+�E+��ܓ�E�4 [�	�x��T0 k� �;��?�U8D"!%�0d   ��O 
   � �8	M,TD���E-T�$}�|�'�E+��ܓ�E�3 [�	�x��T0 k� �+��/�U8D"!%�0d   ��O    � �8	M0TD���E-X�,~�|*'�E+��ܓ�E�2 [�	�x��T0 k� ����U8D"!%�0d  	 $�O    � �8	M8UD���E`�8���*'�E+��̏�E�1 [�	�x��T0 k� <���U8D"!%�0d  	 ��O    � �8	M<UD���Ed�@�|�*'�E+��̏�E�0 n[�	�x��T0 k� <���U8D"!%�0d  	 ��O    � �8	=<UE���El �H�|�*'�E+��̏�C�/ n[�	�x��T0 k� <���U8D"!%�0d  	 ��O    � �8	=@UE�{�Es��P�|�*'�E+��̏�C�/ n[�	�x ��T0 k� <���U8D"!%�0d  	 ��O    � �8	=DUE�w�Ew�|X�|�*'�E+��̏�C�. n[�	�{���T0 k� <���U8D"!%�0d   ��O    � �8	=DUE�o�E{�|`�|�*#�E+��̏�C�- n[�	�{���T0 k� ����U8D"!%�0d   ��O    � �8	=HUE�g�E�|h��*#�E��̏�C�- �[�	�{���T0 k� ����U8D"!%�0d   ��O    � �8	MLUE�[�E��|x�*#�E��̏�C�+ �[�	�{���T0 k� ����U8D"!%�0d   ��O    � �8	MLUFW�E��|��*#�E��̏�C�+ �[�	�{���T0 k� ����U8D"!%�0d   ��O    � �8	MPUFO�B���|��*#�E��̏�C�* �[�	�{���T0 k� ����U8D"!%�0d   ��O    � �8	MPUFK�B�����~�*#�E��̏�C�)N[�	�{���T0 k� ����U8D"!%�0d   ��O    � �8	MPUFC�B�����~�*#�E��̏�C�)N[�	�{���T0 k� ����U8D"!%�0d   ��O    � �8�TUF?�B�����}�*�E��̋�C�(N[�	�{���T0 k� ����U8D"!%�0d   ��O    � 
�8�TUE|;�B�����}ܨ*�E��̋�C�(N[�	�{���T0 k� ����U8D"!%�0d   ��O    � 	�8�TVE|3�E����|ܬ*�E��̋�C� 'N[�	�{���T0 k� L���U8D"!%�0d   ��O    � �8�XVE|+�E����{ܴ*�E��̋�C��&N[�	�{���T0 k� L���U8D"!%�0d   ��O    � �8�\VE|#�E����{ܸ*�E��܋�C��%N[�	�{���T0 k� L���U8D"!%�0d   ��O    � �8�\VE|�E����zܼ*�E���܋�C��%N[�	�{���T0 k� L���U8D"!%�0d   ��O    � �8�`WI��E����y��*�E���܋�C��$^[�	�{���T0 k� ,���U8D"!%�0d   ��O    � �8�`WI��E����x��*�E���܏�C��#^[�	�{���T0 k� ,���U8D"!%�0d   ��O    � �8�dWI��E����w��*�E���܏�C��#^[�	�{���T0 k� ,���U8D"!%�0d   ��O    � �8�hXI��E�����v��*�E�����C��"^[�	�{���T0 k� ,���U8D"!%�0d    ��O    � �8�lYI��E�����u��*�D˿���D�!^[�N{���T0 k� ����U8D"!%�0d    ,�O    �  �8pYI��E�����t�*�D�Ǘ��D�!^[�N{���T0 k� ����U8D"!%�0d    ��O    ����8pYI���E�����r�*�D�Ϙ��D� ^[�N{���T0 k� ����U8D"!%�0d    ��O    ����8tZI���E����q�*�D�ט��D� ^[�N{���T0 k� ����U8D"!%�0d    ��O    ����8tZI���E��� p�*�D�ߙ	���D� ^[�N{���T0 k� ����U8D"!%�0d   ��O    ����8xZI���E���o�*�D��	���D�^[� {���T0 k� ����U8D"!%�0d   ��O    ����8xZF�E���n�*�D��	���D�n[� {���T0 k� ����U8D"!%�0d   ��O    ����8|[F�E���m���D���	���D�n[� {���T0 k� ,���U8D"!%�0d   ��O    ����8|[F�E�'��k���D���	���D�n[� {���T0 k� ,���U8D"!%�0d   ��O    ����8�[F��E�7�} i��D�����D�n[� n{���T0 k� ,���U8D"!%�0d   ��O    ����8�[F��E~;�}$g�
��D�����D�n[� n{���T0 k� ,���U8D"!%�0d   ��    ����8�[F��E~C�}(f�	��D�����D�n[� n{���T0 k� ����U8D"!%�0d   ��    ����8�[F��E~G�},d���D�'����D� �[� n{���T0 k� ����U8D"!%�0d   ��    ����8�[F��E~O�}4c���D�/����D� �[� n{���T0 k� ����U8D"!%�0d   ��    ����8�[F��E~[�}<`�(��D�;�|��D� �[� {���T0 k� ����U8D"!%�0d   ��    ����8�[F��D�c�}@^�,��D�C�|��D� �[� {���T0 k� ����U8D"!%�0d   ��    ����8�[E���D�g�mD]�4��D�K�|��D� n[� {���T0 k� ����U8D"!%�0d   ��    ����8 �[E���D�o�mD]�8��D�O�|��D� n[� ���T0 k� ����U8D"!%�0d   ��    ����8 �[E���D�s�mH[�@ ��D�W�|��D� n[� ���T0 k� ,���U8D"!%�0d   ��    ����8 �[E���D��mLX�K���D�c�|��D� n[������T0 k� ,���U8D"!%�0d   �    ����9 �[FK��D���=LW�S���D�k�|��D� [������T0 k� ,+��/�U8D"!%�0d   ��    ����:��[FK��D���=PU�W���D�s�|��D� [������T0 k� ,7��;�U8D"!%�0d   ��    ����;��[FK��D���=PT}_���D�w�|��D� [������T0 k� �G��K�U8D"!%�0d   ��    ����<��[FK��D���=PR}c���E��lèD� _������T0 k� �S��W�U8D"!%�0d   ��    ����=��[FK��D���=PQ}k���E���lçA�� _������T0 k� �c��g�U8D"!%�0d   ��    ����>                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \���� ]�((  � �          � �w     � �{       <           
   � 8�         ��     ���   (         ��(_   *	      ��"�    ��(_�"�           	               ���          �`     ���   8�           +         ��     *M ��7      �                  .          �      ���   	@
          ����    U       �\�    �����\�                      �$          !      ���   H$
         ��ƿ   � �       .�#x    ��ƿ�#U      ��   
           ���$           & 
`     ���   H
!          �|  ��	      B���     �|���                             ���k              L  ���      0            ��H ^ ^	    V��*[    ��B����    ��:            8����         l��      ��@ 0
%          ��܆  / /     j��5�    ��c����    ��d              #����         p�     ��@   0
          ��i � �
	   ~��eM    �������y    n��            	����         ��  &  ��`  8
           tK�  � �	   ����     t[����    �              Q ����         	 ��    ��h  8         ��k�  T T    ���W    ��|2��S    ����              ����         
 � b     ��@  P	          + ��
	      � �ޝ     + �ޝ                           ��@        ��    �  ��@    P                   ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��"�  ��        �����  ���M4��5  �����                   x                j  �   �	   �                         ��    ��        ���      ��  ��           "                                                �                          �" ���#����������� �������         	  
      
   � 
  lY ܻ�C       �� �o� �� p� � p� �$ q  �D q  �d q@ �$ �r@ �$ s@ �D  s` ބ s� �� s� $d n ��� ���� ����  ����. ����< ����J ����X � 
�\ W  
�< W� 
�� W� 
�\ W� � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }`���� � � }`���� � 
�| V  
�\ V� 
�� V� 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����������� -  ������  
�fD
��L���"����D" � j  "  B   J jF�"    "�j * , ����
��"     �j @�    �
� �  �  
�  I��  ��     �   �        ��     �        t��  ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �      �� �  ���        �t �  ��        �        ��        �        ��        � 	 	  �     /������        ��                         ��  0 � ���                                     �                ����            ������%��  ������                 8 Geoff Sanderson     0:01                                                                        6  4     � �
�b �cj � � cp � �
kV � �k_ �  ka � kb � �k~ � � 	k� � � 
k� � � k� � � k� � � k� � �c� � � c� � � c� � �c� � �c�y � c�q �c�q � c�p � k�| �B� � B�  �"� � "� �"� �*� �"�r � "�� ��r � 
�� � 
�� � 
�� � #"�� �$�q � 
�� � 
��9 
� �3 
� �/)� / 
� �, 
� �( 
� �`  "D ~T  "H �8 /"D ~X  "K �X  "K � � 2*P�P  *RpP  *Rl 5*Fl6*t07*
tP  *C\ 9*Fl:*t0;*
tP  *C\P  *C\P  *C\X  *Kt                                                                                                                                                                                                                         �� P        �     @ 
        �     W P E g  ���� Z    	            	�������������������������������������� ���������	�
��������                                                                                          ��    ��1�� ��������������������������������������������������������   �4, 6� B 	� ?�  F	� Q��� {� ւ@a��6�������� ���	�                                                                                                                                                                                                                                                                                                       @��                                                                                                                                                                                                                                               �        � �   H�J      �                             ������������������������������������������������������                                                                                   	                                                        �             �        �    �   t          
 	  
	 
 	 	 ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� �������            x                 _    (    ��  D�J    	  wI                             ������������������������������������������������������                                                                                                                                     {     �      �        �        � �          	  
 	 
 	 	 ��  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���           t                                                                                                                                                                                                                                                                                                     
        �             


             �  }�         ��������������������  's������������  vo����������������    ������������  's����������������������������                                           R�                    N�               ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" R > / 	               	                 � �Ф� �o�                                                                                                                                                                                                                                                                                     �1n  EY                c      m      l                                                                                                                                                                                                                                                                                                                                                                                                                                        ( s  (s  J�  
�  �  Cm�  ����)��d����� O�#��������̎�U����L����r�          <        �"��         	�   &  AG� �   �                 K��                                                                                                                                                                                                                                                                                                                                      C B   �                     !��                                                                                                                                                                                                                            Y   
�� �� Ѱ��      �� @      ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� ���������  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���   �� �                                                                                                                                                                                                                                                                                                                                                                              