GST@�                                                           @c�                                                      &  �   ��                   ����e � 
 ʱ����������P���z���        �h     #    z���                                d8<n    �  ?     2g����  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"     �j�
�   ��
                                                                                 ����������������������������������       ��    =b 0Qb 4 114  4c  c  c      	 
      	   
       ��G �� � ( �(                 Enn )1         88�����������������������������������������������������������������������������������������������������������������������������o=  0  o4   1  +      '           �                    	�  7�  V�  	�                  n  	          : �����������������������������������������������������������������������������                                �         R�   @  #   }   �                          �                                                     '    E)n1n  	n    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������     4ILo�2K�q/�PNZ|,�áAP�'�H0
p�@hm3�T0 k� �<�@U2d   2$ ! ��O    � <�� 0ILo�3K�q/�RNZ|,�áAP�'�D0
p�@hm3�T0 k� �<�@U2d   2$ ! ��O    � <�� ,JLo�4K�p/�SNZ|,���AP�'�@0
p�@hm3�T0 k� �<�@U2d   2$ ! ��O    � <�� ,JLo�5K�p/�UNZ|,���AP�'�@0
p�@hm3�T0 k� �<�@U2d   2$ ! ��O    � <�� (JLo�7K�o/�WNZ|,���AP�'�<0
p�@hm3�T0 k� L@�DU2d   2$ ! ��O    � <�� $KLo�8K��o��YNZ|,���AP�'�80
p�@hm3�T0 k� L@�DU2d   2$ ! ��O    � <��  KLo�9K��n��[NZ|,���AP�'�80
p�@hm3�T0 k� L@�DU2d   2$ ! ��O    � <�� KLo�:K��n��\NZ|,���AP�'�4/
p�@hm3�T0 k� L@ �D U2d   2$ ! ��O    � <�� KLo�:K��m��^NZ|,���AP�'�0/
p�@hm3�T0 k� L@!�D!U2d   2$ ! ��O    � <�� LLo�;K��m��`NY|,���AP�'�0/
p�@hn3�T0 k� ,@"�D"U2d   2$ ! ��O    � <�� LLo�=K��l��cNY|,���AP�'�(/
p�@hn3�T0 k� ,D#�H#U2d   2$ !  -�O    � <�� MLo�>K��l�|eNY|,���AP�'�(/
p�@hn3�T0 k� ,D$�H$U2d   2$ !  ��O    � <��MLo�?K��k�|fNY|,���AP�'�$/
p�@hn3�T0 k� ,D%�H%U2d   2$ !  ��O    � <��MLo�@K��k�xh>Y|,���AP�'�$/
p�@hn3�T0 k� �D&�H&U2d   2$ !  ��O    � <��NLo�AK��j�xi>Y|,���AP�'� /
p�@hn3�T0 k� �D'�H'U2d   2$ !  ��O    � <��NLo�BK��j�tk>Y|,���AP�'�.
p�@hn3�T0 k� �H(�L(U2d   2$ ! ��O    � <�� NLo�CK��j�tl>Y|,���AP|'�.
p�@hn3�T0 k� �H)�L)U2d   2$ ! ��O    � <���NLo�DK��i�tn>Y|,���AP|'�.
p�@hn3�T0 k� �H*�L*U2d   2$ ! ��O    � <����OLo�DK��i�po>Y|,���AP|'�.
p�@hn3�T0 k� �H*�L*U2d   2$ ! ��O    � <����OLo�EK��h�pq�Y|,���AP|'�.
p�@ln3�T0 k� �H+�L+U2d   2$ ! ��O    � <����OLo�FK��h�lr�Y|,���AP|'�.
p�@ln3�T0 k� ,H,�L,U2d   2$ ! ��O    � <����OLo�GK��h�lt�Y|,���APx'�.
p�@ln3�T0 k� ,L-�P-U2d   2$ ! ��O   � <����PLo�HK��g�hu�Y|,���APx'�.
p�@ln3�T0 k� ,L.�P.U2d   2$ ! ��O    � <���PL_�HK��g�hv�Y|,���APx'�.
p�@ln3�T0 k� ,L/�P/U2d   2$ ! ��O    � <���PL_�IK��g�hx�Y|,���APx'�.
p�@ln3�T0 k� ,L0�P0U2d   2$ ! ��O    � <���PL_�JK��f�dy� Y|,���APx'�-
p�@lo3�T0 k� �L0�P0U2d   2$ ! ��O   � <���QL_�KK��f�dz� Y|,���APx'�-
p�@lo3�T0 k� �L1�P1U2d   2$ ! ��O    � <���QL_�KK��f�`|� Y|,���APt'�-
p�@lo3�T0 k� �L2�P2U2d   2$ ! ��O    � <���QL_�LK��e�`}� Y|,���APt'�-
p�@lo3�T0 k� �P3�T3U2d   2$ !  ��O    � <���QD��MK��e�`~� Y|,���APt'� -
p�@lo3�T0 k� �P4�T4U2d   2$ !  ��O    � <���RD��NK��e�\� X|,���APt'� -
p�@lo3�T0 k� �P5�T5U2d   2$ !  ��O    � <���RD��NK��d�\���X|,���APt'��-
p�@lo3�T0 k� �P6�T6U2d   2$ !  ��O    � <���RD��OK��d�\���X|,���APt'��-
p�@lo3�T0 k� ,P7�T7U2d   2$ !  ��O    � <��/�RD��PK��d�X���X|,���APp'��-
p�@lo3�T0 k� ,P7�T7U2d   2$ !  /�O    � <��/�RE��QK��d�X���X|,���APp'��-
p�@lo3�T0 k� ,T8�X8U2d   2$ !  ��O    � <��/�SE��RK��c�X��X|,���APp'��-
p�@lo3�T0 k� ,T9�X9U2d   2$ !  ��O    � <��/�SE��SK��c�T��X|,���APp'��-
p�@lo3�T0 k� ,T:�X:U2d   2$ !  ��O    � <��/�SE�|TK��c�T��X|,���APp'��-
p�@lo3�T0 k� �T;�X;U2d   2$ !  ��O    � <��/�SE�|UK��b�T��X|,���APp'��,
p�@lo3�T0 k� �T<�X<U2d   2$ !  ��O    � <��/�SL_|VK��b�P~��X|,���APp'��,
p�@lo3�T0 k� �T=�X=U2d   2$ !  ��O    � <��/�TL_|WK��b�P~��X|,���APl'��,
p�@lo3�T0 k� �X=�\=U2d   2$ !  ��O    � <��/�TL_xWK��b�P~��X|,���APl'��,
p�@lo3�T0 k� �X>�\>U2d   2$ !  ��O    � <��/�TL_xXK��b�L~��X|,���APl'��,
p�@lo3�T0 k� �X?�\?U2d   2$ !  ��O    � <��/�TL_xYCO�b�L}��X|,���APl'��,
p�@lo3�T0 k� �X@�\@U2d   2$ !  ��O    � <��/�TL_xZCO�b�L}��X|,���APl'��,
p�@lo3�T0 k� �XA�\AU2d   2$ !  ��O    � <��/�UL_x[CO�b�H}��X|,���APl'��,
p�@lo3�T0 k� �XB�\BU2d   2$ !  ��O    � <��/�UL_x\CO�a�H}��X|,���APl'��,
p�@lp3�T0 k� �XB�\BU2d   2$ !  ��O    � <��/�UL_t\CO�a�H|��X|,���APh'��,
p�@lp3�T0 k� �\C�`CU2d   2$ !  ��O    � <��/�UL_t]CO�a�H|��X|,���APh'��,
p�@pp3�T0 k� �\D�`DU2d   2$ !  ��O    � <��/�ULot^CO�a�D|��X|,���APh'��,
p�@pp3�T0 k� �\E�`EU2d   2$ !  ��O    � <��/�ULot_CO�a�D|��X|,���APh'��,
p�@pp3�T0 k� �\F�`FU2d   2$ !  ��O    � <��/�VLot_CO�a�D|��X|,���APh'��,
p�@pp3�T0 k� �\G�`GU2d   2$ !  ��O    � <��/�VLop`CO�a�D{��X|,���APh'��,
p�@pp3�T0 k� �\G�`GU2d   2$ !  ��O    � <��/�VLopaCO�a�@{��X|,���APh'��,
p�@pp3�T0 k� �`H�dHU2d   2$ !  ��O    � <��/�VLopa@��a�@{��X|,���APh'��,
p�@pp3�T0 k� �`I�dIU2d   2$ !  ��O    � <��/�VLopb@��a�@{��X|,���APh'��+
p�@pp3�T0 k� �`J�dJU2d   2$ !  ��O    � <��/�VLopc@��a�@z��X|,���APd'��+
p�@pp3�T0 k� �`K�dKU2d   2$ !  ��O    � <��/�VLopd@��a�<z��X|,���APd'��+
p�@pp3�T0 k� �`L�dLU2d   2$ !  ��O    � <��/�WLold@��a�<z��X|,���APd'��+
p�@pp3�T0 k� �`L�dLU2d   2$ !  ��O    � <��/�WLoleA�a�<z��X|,���APd'��+
p�@pp3�T0 k� �`M�dMU2d   2$ !  ��O    � <��/�WLoleA�a�<z��X|,���APd'��+
p�@pp3�T0 k� �dN�hNU2d   2$ !  ��O    � <��/�WLolfA�a�8z��X|,���APd'��+
p�@pp3�T0 k� �dO�hOU2d   2$ !  ��O    � <��/�WLolgA�a�8y��X|,���APd'��+
p�@pp3�T0 k� �dP�hPU2d   2$ !  ��O    � <��/�WLolgA�a�8y��X|,���APd'��+
p�@pp3�T0 k� �dQ�hQU2d   2$ !  ��O    � <��/�WLolhA�a�8y��X|,���APd'��+
p�@pp3�T0 k� �dQ�hQU2d   2$ !  ��O    � <��/�XLohiA�a o8y��X|,���APd'��+
p�@pp3�T0 k� �dR�hRU2d   2$ !  ��O    � <��/�XLohiA�a o4y��X|,���AP`'��+
p�@pp3�T0 k� �hS�lSU2d   2$ !  ��O    � <��/�XLohjA�a o4y��X|,���AP`'��+
p�@pp3�T0 k� �hT�lTU2d   2$ !  ��O    � <��/�XLohjA�a o4x��X|,���AP`'��+
p�@pp3�T0 k� �hU�lUU2d   2$ !  ��O    � <��/�XLohkA_�a o4x��W|,���AP`'��+
p�@pp3�T0 k� �hU�lUU2d   2$ !  ��O    � <��/�XLohkA_�a 8x��W|,���AP`'��+
p�@pp3�T0 k� �hV�lVU2d   2$ !  ��O    � <��/�XLohlA_�a 8x��W|,���AP`'��+
p�@pp3�T0 k� �hW�lWU2d   2$ !  ��O    � <��/�XLohlA_�a 8w��W|,���AP`'��+
p�@pp3�T0 k� �hX�lXU2d   2$ !  ��O    � <��/�XLohlA_�a 8w=�W|,���AP`'��+
p�@pp3�T0 k� �lY�pYU2d   2$ !  ��O    � <���YLollA_�a 8w=�W|,���AP`'��+
p�@pp3�T0 k� �lY�pYU2d   2$ !  ��O    � <���YLollA_�a�8w=�W|,���AP`'��+
p�@pp3�T0 k� �lZ�pZU2d   2$ !  ��O    � <���YLollA_�a�8w=�W|,���AP`'��+
p�@pq3�T0 k� �l[�p[U2d   2$ !  ��O    � <���YLolmA_�a�8w=�W|,���AP`'��+
p�@pq3�T0 k� �l\�p\U2d   2$ !  ��O    � <���YLolmA_�a�8w=�W|,���AP\'��+
p�@pq3�T0 k� �l]�p]U2d   2$ !  ��O    � <���YLopmA_�a�8w=�W|,���AP\'��*
p�@pq3�T0 k� �l]�p]U2d   2$ !  ��O    � <���YLopmA_�a�<w=�W|,���AP\'��*
p�@pq3�T0 k� �p^�t^U2d   2$ !  ��O    � <���YLopmA_�a�<w=�W|,���AP\'��*
p�@pq3�T0 k� �p_�t_U2d   2$ !  ��O    � <���YLotmA_�a�<w=�W|,���AP\'��*
p�@pq3�T0 k� �p`�t`U2d   2$ !  ��O    � <���YLotmA_�a�<w=�W|,���AP\'��*
p�@pq3�T0 k� �pa�taU2d   2$ !  ��O    � <���YLotmA_�a�<v=�W|,���AP\'��*
p�@pq3�T0 k� �pa�taU2d   2$ !  ��O    � <���YLoxmA_�a�@v=�W|,���AP\'��*
p�@pq3�T0 k� �pb�tbU2d   2$ !  ��O    � <���YLoxmA_�a�@v=�W|,���AP\'��*
p�@pq3�T0 k� �pc�tcU2d   2$ !  ��O    � <���YLoxmL�a�@uM�W|,���AP\'��*
p�@pq3�T0 k� �td�xdU2d   2$ !  ��O    � <���YLo|mL�a�DuM�W|,���AP\'��*
p�@tq3�T0 k� �td�xdU2d   2$ !  ��O    � <���YLo|mL�a�DuM�W|,���AP\'��*
p�@tq3�T0 k� �te�xeU2d   2$ !  ��O    � <���YL_|mL�a�DuM�W|,���AP\'��*
p�@tq3�T0 k� �tf�xfU2d   2$ !  ��O    � <���YL_�mL�a�DuM�W|,���AP\'��*
p�@tq3�T0 k� �tg�xgU2d   2$ !  ��O    � <���YL_�mL�a�DuM�W|,���AP\'��*
p�@tq3�T0 k� �th�xhU2d   2$ !  ��O    � <���YL_�mL�a�DtM�W|,���APX'��*
p�@tq3�T0 k� �th�xhU2d   2$ !  ��O    � <���YL_�mL�a�HtM�W|,���APX'��*
p�@tq3�T0 k� �xi�|iU2d   2$ !  ��O    � <���YL_�lL�a�HsM�W|,���APX'��*
p�@tq3�T0 k� �xj�|jU2d   2$ !  ��O    � <���YE��lL�a�LsM�W|,���APX'��*
p�@tq3�T0 k� �xk�|kU2d   2$ !  ��O    � <���YE��lL�a�LrM�W|,���APX'��*
p�@tq3�T0 k� �xk�|kU2d   2$ !  ��O    � <���YE��mL�a�LrM�W|,���APX'��*
p�@tq3�T0 k� �xl�|lU2d   2$ !  ��O    � <���YE��lL�a�LrM�W|,���APX'��*
p�@tq3�T0 k� �xm�|mU2d   2$ !  ��O    � <���YE��lL�a�LqM�W|,���APX'��*
p�@tq3�T0 k� �xn�|nU2d   2$ !  ��O    � <���YL_�lL/�a�PpM�W|,���APX'��*
p�@tq3�T0 k� �|n��nU2d   2$ !  ��O    � <���YL_�lL/�a�PpM�W|,���APX'��*
p�@tq3�T0 k� �|o��oU2d   2$ !  ��O    � <���YL_�lL/�a�ToM�W|,���APX'��*
p�@tq3�T0 k� �|p��pU2d   2$ !  ��O   � <���YL_�lL/�a�XnM�W|,���APX'��*
p�@tq3�T0 k� �|q��qU2d   2$ !  ��O    � <��/�YL_�lL/�a�XmM�W|,���APX'��*
p�@tq3�T0 k� �|q��qU2d   2$ !  ��O    � <��/�YL_�lL/�a�\lM�W|,���APX'��*
p�@tq3�T0 k� �|r��rU2d   2$ !  ��O    � <��/�YL_�lL/�a�\lM�W|,���APX'��*
p�@tq3�T0 k� �|s��sU2d   2$ !  ��O    � <��/�YL_�lL/�a�\kM�W|,���APX'��*
p�@tq3�T0 k� ��t��tU2d   2$ !  ��O    � <��/�YL_�lL/�a�`jM�W|,���APX'��*
p�@tq3�T0 k� ��t��tU2d   2$ !  ��O    � <��/�YL_�lL/�a�diM�W|,���APX'��*
p�@tq3�T0 k� ��u��uU2d   2$ !  ��O    � <��/�YL_�lL/�a�diM�W|,���APX'��*
p�@tq3�T0 k� ��v��vU2d   2$ !  ��O    � <��/�YLo�lL/�a�hhM�W|,���APX'��*
p�@tq3�T0 k� ��w��wU2d   2$ !  ��O    � <��/�YLo�lL/�a�hhM�W|,���APX'��*
p�@tq3�T0 k� ��w��wU2d   2$ !  ��O    � <��/�YLo�lL/�a�lhM�W|,���APT'��*
p�@tq3�T0 k� ��x��xU2d   2$ !  ��O    � <��/�YLo�lL/�a�lhM�W|,���APT'��*
p�@tq3�T0 k� ��y��yU2d   2$ !  ��O    � <��/�XLo�lL/�a�lhM�W|,���APT'��*
p�@tq3�T0 k� ��z��zU2d   2$ !  ��O    � <��/�XLo�lL/�a�phM�W|,���APT'��*
p�@tr3�T0 k� ��z��zU2d   2$ !  ��O    � <��/�WLo�lL/�a�thM�W|,���APT'��*
p�@tr3�T0 k� ��{��{U2d   2$ !  ��O    � <��/�WLo�lL/�a�thM�W|,���APT'��*
p�@tr3�T0 k� ��|��|U2d   2$ !  ��O    � <��/�VLo�lL/�a�xhM�W|,���APT'��*
p�@tr3�T0 k� ��}��}U2d   2$ !  ��O    � <��/�VLo�lL/�`�|gM�W|,���APT'��*
p�@tr3�T0 k� ��}��}U2d   2$ !  ��O    � <��/�VLo�mL/�`�|gM�W|,���APT'��*
p�@tr3�T0 k� ��~��~U2d   2$ !  ��O    � <��/�ULo�mL/�`��gM�W|,���APT'��*
p�@tr3�T0 k� ����U2d   2$ !  ��O    � <��/�ULo�mL/�`��gM�W|,���APT'��*
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�ULo�mL/�`��gM�W|,���APT'��*
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�TLo�mL/�`��gM�W|,���APT'��*
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�TLo�mL/�`��gM�W|,���APT'��*
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�SLo�mL/�`��g=�W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�SLo�mL/�`��g=�W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�SLo�mL/�_��g=�W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�RLo�nL/�_��g=�W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�RLo�nL/�_��g=�W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�RLo�nL/�_��g=�W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�QLo�nL/�_ߐg��W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�QLo�nL/�_ߐg��W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�QLo�nL/�_ߔg��W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�QLo�nL/�_ߔf��W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�PLo�nL/�_ߘf��W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�PLo�nL/�_ߘf��W|,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�PLo�nL/�_ߜe��W!�,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�OLo�oL/�^ߠe��W!�,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�OLo�oL�^ߠd��W!�,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�OLo�oL�^ߤd��W!�,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�OLo�oL�^�d��W!�,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <��/�NLo�oL�^�c��W!�,���APT'��)
p�@tr3�T0 k� ������U2d   2$ !  ��O    � <���NLo�oL�^�c��W!�,���APT'��)
p�@tr3�T0 k� ����U2d   2$ !  ��O    � <���NLo�oL�^�c��W!�,���APT'��)
p�@tr3�T0 k� ����U2d   2$ !  ��O    � <���MLo�oL�^�c��W!�,���APP'��)
p�@tr3�T0 k� ����U2d   2$ !  ��O    � <���MLo�oL�^�b��W!�,���APP'��)
p�@tr3�T0 k� ����U2d   2$ !  ��O    � <���MLo�oL�^�b��W!�,���APP'��)
p�@tr3�T0 k� ����U2d   2$ !  ��O    � <���MLo�oA_�^�b��W|,���APP'��)
p�@tr3�T0 k� ��~��~U2d   2$ !  ��O    � <����MLo�oA_�^�b��W|,���APP'��)
p�@tr3�T0 k� ��~��~U2d   2$ !  ��O    � <����LL_�pA_�^�b��W|,���APP'��)
p�@tr3�T0 k� ��~��~U2d   2$ !  ��O    � <����LL_�pA_�^�b��W|,���APP'��)
p�@tr3�T0 k� ��~��~U2d   2$ !  ��O    � <����LL_�pA_�^��b��W|,���APP'��)
p�@tr3�T0 k� ��~��~U2d   2$ !  ��O    � <����KL_�pC��^��b��W|,���APP'��)
p�@tr3�T0 k� ��~��~U2d   2$ !  ��O    � <����KL_�pC��^��b��W|,���APP'��)
p�@tr3�T0 k� ��}��}U2d   2$ !  ��O    � <����KL_�pC��^��b��W|,���APP'��)
p�@tr3�T0 k� ��}��}U2d   2$ !  ��O    � <����KA��pC��^��b��W|,���APP'��)
p�@tr3�T0 k� ��}��}U2d   2$ !  ��O    � <����KA��pC��^O�b��W|,���APP'��)
p�@tr3�T0 k� ��}��}U2d   2$ !  ��O    � <����KA��pC��^O�b��W|,���APP'��)
p�@tr3�T0 k� ��}��}U2d   2$ !  ��O    � <����KA��qC��^O�b��W!�,���APP'��)
p�@tr3�T0 k� ��}��}U2d   2$ !  ��O    � <����KA��qC��^O�b��W!�,���APP'��)
p�@tr"��T0 k� ��|��|U2d   2$ !  ��O    � <����KF�qC��^O�b��W!�,���APP'��)
p�@tr"��T0 k� ��|��|U2d   2$ !  ��O    � <����KF�rC��^O�b��W!�,���APP'��)
p�@tr"��T0 k� ��|��|U2d   2$ !  ��O    � <����KF�rC��^O�b��W!�,���APP'��)
p�@tr"��T0 k� ��|��|U2d   2$ !  ��O    � <����KF�rC��^O�b��W!�,���APP'��)
p�@tr"��T0 k� ��|��|U2d   2$ !  ��O    � <��O�KF�rC��^O�b��W!�,���APP'��)
p�@tr"��T0 k� ��|��|U2d   2$ !  ��O    � <��O�KE��sC��^O�b��W!�,���APP'��)
p�@tr"��T0 k� ��|��|U2d   2$ !  ��O    � <��O�KE��sC��^O�b��W!�,���APP'��)
p�@tr"��T0 k� ��{��{U2d   2$ !  ��O    � <��O�KE��sC��^O�b��W!�,���APP'��)
p�@tr"��T0 k� ��{��{U2d   2$ !  ��O    � <��O�KE��tA_�^O�b��W!�,���APP'��)
p�@tr"��T0 k� ��{��{U2d   2$ !  ��O    � <�� �KE� tA_�^O�b��W|,���APP'��)
p�@tr"��T0 k� ��{��{U2d   2$ !  ��O    � <�� �KE�tA_�^O�b��W|,���APP'��)
p�@tr3�T0 k� ��{��{U2d   2$ !  ��O    � <�� �KE�tA_�^O�b��W|,���APP'��)
p�@tr3�T0 k� ��{��{U2d   2$ !  ��O    � <�� �KE�tA_�^�b��W|,���APP'��)
p�@tr3�T0 k� ��z��zU2d   2$ !  ��O    � <�� �KE�tA_�^�b��W|,���APP'��)
p|@tr3�T0 k� ��z��zU2d   2$ !  ��O    � <���jA��@��vqpX!_�|,�˃Bèz�/���BC4|�T0 k� ��p� pU2d   2$ !  ��     � ; �jA��@��vqpZ![�|,�ӄBð|�/���B�8|�T0 k� ��n��nU2d   2$ !  ��     � < �jA��@��vqp\!W�|,�ۄBø}�0���B�8|�T0 k� ��m��mU2d   2$ !  ��     � < �kD3�@��vqp^!W�|,��Bü~�0���B�8|�T0 k� ��l��lU2d   2$ !  ��     � < � kD3�@��vqp_!S�|,��B���1���B�<{�T0 k� ��k��kU2d   2$ !  ��     � < ��lD3�CB�uqpc!O�|,���IЀ�2���B�<{�T0 k� ��k��kU2d   2$ !  ��     � < ��lD3�CB�u	Qpe!O�|,��IԀ�2���B�D{�T0 k� ��j��jU2d   2$ !  ��     � < ��mD3߳CB�u	Qpf�K�|,��I��2���B�Lz�T0 k� ��k��kU2d   2$ !  ��     � < ��mD3ߴCB�t	Qph�K�|,��I��3���B�Tz�T0 k� ��k��kU2d   2$ !  ��     � < ��mD3ߴCB�t	Qpi�K�|,��I�~�3���B�\z"T0 k� ��k��kU2d   2$ !  ��     � < ��mDC۴E��s	Qpk�G�|,�#�I#�~ �3���B�dz"T0 k� ��f��fU2d   2$ !  ��     � < ��nDC׵E��r	Qpn�G�|,�3�I#�} �4���B�ty"T0 k� ��b��bU2d   2$ !  ��     � < ���nDC׶E��q	apo�G�|,�;�I#�| �4���B�|y"T0 k� ��_��_U2d   2$ !  ��     � < ��nDCӷE��q	app�G�|,�C�I#�{ �5���B��y"T0 k� ��]��]U2d   2$ !  �     � < �#�nDCϷE��p	apr�G�|,�K�I�{25���B��y"T0 k� ��\��\U2d   2$ !  ��    � < �#�nDCϸE��o	aps�G�|,�O�I�z26���O��y"T0 k� ��Z��ZU2d   2$ ! �    � < �#�kDCǹE��m!pu�G�|,�_�I�y27���O��x"T0 k� �hV�lVU2d   2$ ! ��    � < �#�jDCǺE��l!pvG�|,�g�I�x28���O��x"T0 k� �\T�`TU2d   2$ ! ��/    � < �S�iDCûE��l!pxC�|,�k�I#�x"8���O��x�T0 k� �PR�TRU2d   2$ ! ��/    � < �S�hE�EB�k!tyC�|,�s�I#�w"9���O��w�T0 k� �DP�HPU2d   2$ ! ��/    � < �S�eE�EB�i!txC�|,��I#�v";���O��w� T0 k� �,L�0LU2d   2$ ! ��/    � < �S�dE�EB�h!txC�|,Ç�I#�v";���O��w��T0 k� � K�$KU2d   2$ ! ��/    � < �S�cE�EB�g!xxC�|,Ë�I�u<���O��v�T0 k� �I�IU2d   2$ ! ��/    � < �c�bE��E2�exwC�|,Ï�I�u=���O��v�T0 k� �G�GU2d   2$ ! ��/    � < �c�aE��E2�d|wC�|,×�I�u>���O��v�T0 k� ��E� EU2d   2$ ! ��/    � < �c�_E��E2�b�wC�|,ß�I t?���O��u�T0 k� ��A��AU2d   2$ ! ��/    � < �c�^E��E2�a�vC�|,ã�I$ t@���O��u�T0 k� ��?��?U2d   2$ ! ��/    � < �c�\D���CB�_�vC�|,ç�I$ t @���O��u�T0 k� ��=��=U2d   2$ ! ��/    � < �c�[D���CB�^�vC�|,ë�I$ t A���O��t�T0 k� ��;��;U2d   2$ ! ��/    � < �s�ZD���CB�]��uC�|,ï�I$ t$B���O��t�T0 k� ��:��:U2d   2$ ! ��/    � < �s�XD���CB�Z��uC�|,ӷ�I s,C b��O��s�T0 k� ��6��6U2d   2$ ! ��/    � < �s�XD���CB�X��t?�|,ӻ�Is0D b��O��s�T0 k� ��4��4U2d   2$ ! ��/    � < �s�WD���CB�W��t?�|,ӻ�Is4D b��O��s�T0 k� ��2��2U2d   2$ ! ��/    � < �s�VD���CB�U��t?�|,ӿ�Is8E b��O��r�T0 k� �|0��0U2d   2$ ! ��/    � < �s�UD���CB�Tќs?�|,�ïIs<E b��O��r�T0 k� �p.�t.U2d   2$ ! ��/    � < �s�TD���CB�RѠs?�|,�ðE�s�@F b��O��r3�T0 k� �d,�h,U2d   2$ ! ��/    � < �s�RD���CB�OѨq!?�|,�ǳE�s�HG b��O��q3�T0 k� �P+�T+U2d   2$ ! ��(    � < �s�QD���CR�MѬq!?�|,�ǴE�s�LG ���E��q3�T0 k� �X,�\,U2d   2$ ! ��(    � < �s�PD���CR�KѰp!?�|,�ǶE�s�PH ���E��q3�T0 k� �`-�d-U2d   2$ ! ��(    � < �s�OD���CR�IѴo!?�|,�˷E�r�TH ���E��p�T0 k� �d/�h/U2d   2$ ! ��(    � < �s�ND��CR�FѼn!?�|,�˺E�$r�`I ���E��p�T0 k� �p0�t0U2d   2$ !  ��(    � < �s�MI�{�CR�D��m!?�|,�˻E�(q�dI ���E��o�T0 k� �t0�x0U2d   2$ !  .�(    � < �s�LI�{�CR�B��l!?�|,�˼E�,q�hI ���E��o�T0 k� �x1�|1U2d   2$ !  ��(   � < �s�KI�w�CR�@��k!?�|,�˽E�0q�pI ���E��o�T0 k� ��1��1U2d   2$ !  ��(    � < �s�JI�w�CR�>��k!C�|,�˿E�4p�tI ���E��n�T0 k� ��1��1U2d   2$ !  ��(    � < �s�IEcs�CR�:��i�C�|,���E�<or|I ���E��n�T0 k� ��1��1U2d   2$ !  ��(    � < �s�HEco�Cb�8��h�C�|,���E�@or�I ���E��m�T0 k� ��1��1U2d   2$ !  ��(    � < �s�GEck�Cb�6��g�G�|,���E�@nr�I ���E��m�T0 k� ��1��1U2d   2$ !  ��(    � < �s�GEck�Cb�4��f�G�|,���E�Dmr�I ���E��l�T0 k� ��1��1U2d   2$ !  ��(   � < �s�EEcc�Cb�0��d!K�|,��E�Llr�H ���E��k�T0 k� ��0��0U2d   2$ !  $�(    � < �s�DEcc�Cb�.��c!O�|,��E�Pkr�H ���E��j�T0 k� ¤0��0U2d   2$ !  ��(    � < �s�DEc_�E2�,� b!O�|,��E�Tjr�H ���E��j�T0 k� ¨0��0U2d   2$ !  ��(    � < �s�CEc[�E2�*�a!S�|,��E�Xir�G ���E��i�T0 k� °/��/U2d   2$ !  ��(    � < �s�BESW�E2�'r`!S�|,��E�Xhr�G ���E��h�T0 k� ´/��/U2d   2$ !  ��(    � < �s�AESO�E2�#r]!W�|,��E�`fr�F ���E� g�T0 k� ��.��.U2d   2$ !  ��(    � < �s�@ESK�E2�!r\![�|,��E�`eb�E ���E�f�T0 k� ��/��/U2d   2$ !  ��(    � < �s�@ES?�E2�r [!_�|,��E�ddb�E ���E�e�T0 k� ��/��/U2d   2$ !  ��(    � < �s�?C�7�E2�r$Y!c�|,��E�dcb�D��E�d�T0 k� ��0��0U2d   2$ !  ��(    � < �s�>C�( E2�r,X`|,��E�hbb�C��E�c�T0 k� ��0��0U2d   2$ !  ��(    � < �s�=C�( E2�r4Uh|,��E�h`b�B��E�a�T0 k� ��/��/U2d   2$ !  ��(    � < �s�=C� E"�r8Tl|,��E�l_b�A��E�`�T0 k� ��.��.U2d   2$ !  ��(    � < �s�<OSE"�r@Rl|,��E�l^b�@���E�_�T0 k� ��-��-U2d   2$ !  ��(    � < �s�;OSE"�rDQ	p|,��E�l\b�?���E�^�T0 k� ��,��,U2d   2$ !  ��(    � < �s�:OSE"�rLM	t	|,��E�pZb�>���E�\�T0 k� ��+��+U2d   2$ !  ��(    � < �s�:OS
E"�bPL	t
|,�{�E�pYR�=���C�[�T0 k� ��1��1U2d   2$ !  ��(    � < �s�9OS
E"�bTJ	x|,�w�E�pXR�<ҿ�C�Y�T0 k� ��5��5U2d   2$ !  ��(    � < �s�8OSE"�bXH ax|,�s�C�lWR�;һ�C�X�T0 k� ��8��8U2d   2$ !  ��(    � < �s�7OR�E"�	b`E a||,�g�C�lTR�:ҳ�C�V�T0 k� ��9��9U2d   2$ !  ��(    � < �s�7OR�E"�bdC a�|,�_�C�lSR�9ҫ�E�U�T0 k� ��;��;U2d   2$ !  ��(    � < �s�6OR�E"�bhA a�|,[�C�lRR�8R��E�S�T0 k� ��;��;U2d   2$ !  ��(    � < �s�5OR�E�bl>��|,O�C�hPR�6R��E�Q�T0 k� ��:��:U2d   2$ !  ��(    � < �s�5OR�E�bp<��|,G�C�dOB�6R��E�P�T0 k� ��=��=U2d   2$ !  ��(    � < �s�4OR�E�bp:��|,?�C�dNB�5R��E�N�T0 k� ��>��>U2d   2$ !  ��(    � < �s�4OR�E�bt8��|,7�C�`MB�5B��E�M�T0 k� ��?��?U2d   2$ !  ��8    � < �s�3OR�E� Rt5��|,+�C�\KB�4B��E�J�T0 k� ��@��@U2d   2$ !  ��8    � < �s�2OR�E��Rx3��|,#�C�XJ�3B�E�I�T0 k� ��A��AU2d   2$ !  ��8    � < �s�2OR�E��Rx1��|,�C�XI�3Bw�E�H�T0 k� ��A��AU2d   2$ !  ��8    � < �s�1OR�E��Rx.��|,�C�PG�2Bk�E�E�T0 k� ��A��AU2d   2$ !  ��8    � < �s�0OR�E��R|,�� |,�C�PG�2Bg�E�D�T0 k� ��@��@U2d   2$ !  ��8    � < �s�0OR�E��R|*��!|,��C�LF�1B_�E�C�T0 k� ��@��@U2d   2$ !  ��8    � < �s�/OR�E��R|)��#|,��C�LF�1BW�E�A�T0 k� ��@��@U2d   2$ !  ��8    � < �s�/OR� E��Rx'��$|,��C�HE�12S�E�@�T0 k� ��@��@U2d   2$ !  ��8    � < �s�.ER� E��Rx$��'|,��C�HE"�22G�E��>�T0 k� ��@��@U2d   2$ !  ��8    � < �s�.ER� E��Rx"��)|,��C�DD"�22?�E��=�T0 k� ��@��@U2d   2$ !  ��8    � < �s�-ER�!E��Rx!��+|,���D@C"�32;�E��<�T0 k� ��A��AU2d   2$ !  ��8    � < �s�-ER�!E��Bt��,|,���D<B"�323�E��:�T0 k� ��B��BU2d   2$ !  ��8    � < �s�,ER�"@b��Bp��0|,���D4A"�42+�E��8�T0 k� ��C��CU2d   2$ !  ��8    � < �s�,ER�"@b��Bpѐ1|,һ�D0@"�52#�E��7�T0 k� ��C��CU2d   2$ !  ��8    � < �s�+EB�"@b��Bpѐ3|,��D,?"�52�E��6�T0 k� ��D��DU2d   2$ !  ��8    � < �s�+EB�#@b��Bhь6|,��D$="�62�E��5�T0 k� ��E��EU2d   2$ !  ��8    � < �s�*EB�#E���Bhь7|,��D <2�72�E��4�T0 k� ��G��GU2d   2$ !  ��8    � < �s�*EB�#E���Bd�9|,��D<2�8"�D3�4�T0 k� �|H��HU2d   2$ !  ��8    � < �s�(EB�#E����`�<|,2��D:2�9!��D3�3�T0 k� �xI�|IU2d   2$ !  ��8    � < �s�(EB�#E����\�>|,2��D:2�:!��D3�3�T0 k� �tJ�xJU2d   2$ !  ��8    � < �s�'EB�#E����X�?|,2�D:2�;!��D3�2�T0 k� �pK�tKU2d   2$ !  ��8    � < s�&EB�#E��T�xB|,2s�D9Ҝ=!��E��2�T0 k� �lG�pGU2d   2$ !  ��8    � < |s�%EB�#E��P�tC|,Rk�D9Ҕ=!��E��1�T0 k� �lD�pDU2d   2$ !  ��8    � < ys�$E2�"E��L�pE|,Rc�D 9Ґ>!��E��1�T0 k� �hB�lBU2d   2$ !  ��8    � < ws�#E2x"E��D�hG|,RS�D 9҈@!��E�1�T0 k� �`B�dBU2d   2$ !  ��8    � < ts�"E2p"E��@�dI|,RK�D�8҄@!��E�0�T0 k� �\A�`AU2d   2$ !  ��H    � < qs�"E2l!E҇��<A`J|,RC�D�8ҀA!��E�0�T0 k� �XA�\AU2d   2$ !  ��H    � < ns� CBd E҃��4AXM|,�3�D�7�tC��E�0�T0 k� �LB�PBU2d   2$ !  ��H    � < ks� CB` E���0ATN|,�+�C��7�pC��E�0�T0 k� �HA�LAU2d   2$ !  ��H    � < hs�CBXE���,
APP|,�#�C��7�hD��E�0�T0 k� �@B�DBU2d   2$ !  ��H    � < es�CBTC�{��(
ALQ|,��C��6�dE��E�0�T0 k� �<C�@CU2d   2$ !  ��H    � < bs�CBLC�s��	A@T|,��C��6�XF�E�0�T0 k� �0D�4DU2d   2$ !  ��H    � < _s|CBHC�o��A<V|,���C��5�PG�E�1�T0 k� �(E�,EU2d   2$ !  ��H    � < \s|CBDC�k��A8X|,���C��5�LH��E�1�T0 k� �$F�(FU2d   2$ !  ��H    � < YsxCR@C�g���0Y|,���C��5�DH��E�x1�T0 k� �F� FU2d   2$ !  ��H    � < VsxCR8C�_���(\|,���C�5�8J��E�l2�T0 k� �H�HU2d   2$ !  ��H    � < S�tCR4C�[��� ^|,���C�5�0J��E�h2�T0 k� �H�HU2d   2$ !  ��H    � < P�tCR0C�W���`|,���C�5b(K��E�d2�T0 k� ��I��IU2d   2$ !  ��H    � < M�pCR,C�O���a|,���C�4b K��E�\3�T0 k� ��J��JU2d   2$ !  ��H    � < J�pCR,C�G���e|,��C�4bM��FT4�T0 k� ��K��KU2d   2$ !  ��H    � < G�lCR(C�C���f|,��C�4bM��FL4�T0 k� ��K��KU2d   2$ !  ��H    � < D�lCR$C�;���� h|,��C�3bN��FH5�T0 k� ��L��LU2d   2$ !  ��H    � < A�lCR$C�7�Q���i|,��C�3a�N��	FD6�T0 k� ��M��MU2d   2$ !  ��H    � < >�hCb C�3�Q���k|,��C�3a�O��	F<6�T0 k� ��M��MU2d   2$ !  ��H    � < ;chCb C�+�Q���m|,��C�3a�P��	F87�T0 k� ��N��NU2d   2$ !  ��H    � < 8chCbC�'�Q���n|,��C�3a�P��
F48�T0 k� ��N��NU2d   2$ !  ��H    � < 5cdCbC��Q���r|,�o�C�t2a�Q��F,9�T0 k� ��P��PU2d   2$ !  ��H    � < 2cdCbC��Q���s|,g�Dl2q�R��F(:3�T0 k� �|Q��QU2d   2$ !  ��H    � < /c`CbE��Q���u|,_�Dh2q�R��F$;3�T0 k� �xS�|SU2d   2$ !  ��H    � < ,c`CbE��Q���w|,W�D`2q�S��F ;3�T0 k� �tT�xTU2d   2$ !  ��H    � < )c`CbE���Q���x|,O�DX2q�S��E�<3�T0 k� �lU�pUU2d   2$ !  ��H    � < &c\CbE���Q���z|,G�DP1q�T��E�=3�T0 k� �dU�hUU2d   2$ !  ��H    � < #c\CbE���Q�м{|,�;�DL1ѤT��E�>�T0 k� �dU�hUU2d   2$ !  ��H    � <  S\CrE���Q�и}|,�3�DD1јU��E�>�T0 k� �dT�hTU2d   2$ !  ��H    � < SXCrE���Q�Ь�|,�#�D41шV��B�@�T0 k� �XT�\TU2d   2$ !  ��H    � < STCr E���Q�Ф�|,��D,1рV��B�A�T0 k� �PT�TTU2d   2$ !  ��H    � < STCr E���Q�Р|,��D$0�xW��B�A3�T0 k� �LT�PTU2d   2$ !  ��H    � < SPCq�
E���Q�И|,1�D0�pW��B�B3�T0 k� �HP�LPU2d   2$ !  ��H    � < SLCq�	E��Q�Д|,1�D0�hX��B�C3�T0 k� �DL�HLU2d   2$ !  ��H    � < CLCq�	E��Q�Ќ~|,0��D0�`X��B�C3�T0 k� �<I�@IU2d   2$ !  ��H    � < CDCq�E��Q�Ѐ}|,0��D�0�LY��B�E3�T0 k� �,H�0HU2d   2$ !  ��H    � < 
C@Cq�E��Q��x}|,0��D�/�DY��B�E3�T0 k� � F�$FU2d   2$ !  ��H    � < C@CA�E����p}|,0��D�/�<YфB�F3�T0 k� �E�EU2d   2$ !  ��H    � < �<CA�E����h||,0��D�/�4YфB�G3�T0 k� �D�DU2d   2$ !  ��H    � < �8CA�E����d||,0��D�/�,YфB�G3�T0 k� �D�DU2d   2$ !  ��H    � <���4CA�E����\||,0��D�/�$YфB�H3�T0 k� � C�CU2d   2$ !  ��H    � <���0CA� D1w���T{|,0��D�/�YшB�I3�T0 k� ��C��CU2d   2$ !  ��H    � <���(E���D1g���D{|,0��C�.�Y1�B�J3�T0 k� ��C��CU2d   2$ !  ��H    � <���$E���D1_���<{|,@��C�.� Y1�B�J3�T0 k� ��C��CU2d   2$ !  ��H    � <���E���D1W���4z|,@��C�.��Y1�B�K3�T0 k� ��C��CU2d   2$ !  ��H    � <���E���D1O���,z|,@��C�.��Y1�E�L3�T0 k� ��C��CU2d   2$ !  ��H    � <���
E���D1G���$z|,@��C�.��Y1�E�L3�T0 k� ��C��CU2d   2$ !  �H    � <���
E���D1?�A��y|,@�AR�.��Y
q�E�M3�T0 k� ��B��BU2d   2$ !  �H    � <���
E���D17�A��y|,�w�AR|.��Y
q�E�M3�T0 k� ��B��BU2d   2$ !  ��H    � <����
E���D1#�A��x|,�g�ARl-`�X
q�E�N3�T0 k� ��C��CU2d   2$ !  ��H    � <����
E���D1�A|��x|,�_�ARd-`�X
q�E�O3�T0 k� ��C��CU2d   2$ !  ��H    � <����
E���DA��t��w|,�[�AR\-`�W
q�E�O3�T0 k� ��D��DU2d   2$ !  ��H    � <����	E���DA��p��w|,�S�ARP-`�W
q�E�P3�T0 k� ��D��DU2d   2$ !  ��H    � <����	E���DA��l��v|,�K�ARH-`�W
q�E�P3�T0 k� ��D��DU2d   2$ !  ��H    � <����	E���D@���h��v|,�C�AR@-`�V
q�@Q3�T0 k� �tC�xCU2d   2$ !  ��H    � <����	E���D@���d��u|,�;�AR8-`�V
q�@Q3�T0 k� �hC�lCU2d   2$ !  ��H    � <����	E���D@���`��u|,�7�AR0-`�U
q�@R3�T0 k� �`B�dBU2d   2$ !  ��H    � <����	Eѳ�D@���\��t|,�/�AR,-`�U
q�@R3�T0 k� �XB�\BU2d   2$ !  ��H    � <��B�	Eѯ�E����X��t|,�'�AR$,`|T
q�@ S3�T0 k� �PA�TAU2d   2$ !  ��H    � <��B�	Eѫ�E����T��s|,�#�AR,`tS
q�@ S3�T0 k� �DA�HAU2d   2$ !  ��H    � <��B�	Eѧ�E����P��s|,��AR,`lS
q�@ T3�T0 k� �<@�@@U2d   2$ !  ��H    � <��B�	Eѣ�E����L��r|,��AR,`dR
q�@$T3�T0 k� �4?�8?U2d   2$ !  ��H    � <��B�	Eџ�E���H��r|,��AR,`\Q
q�@$U3�T0 k� �,?�0?U2d   2$ !  ��H   � <��B�	Eћ�E���D��q|,��AR ,`TQ
q�@$U3�T0 k� �$>�(>U2d   2$ !  ��H    � <��B�	Eѓ�E��D��q|,��AQ�,`LP
q�@(V3�T0 k� �=� =U2d   2$ !  ��H    � <��B�	Eя�E��@��p|,���AQ�,`DO
q�@(V3�T0 k� �=�=U2d   2$ !  ��H    � <��B�	Eы�E���<��p|,���AQ�,`<O
q�@(V3�T0 k� �<�<U2d   2$ !  ��H    � <��B�
Eу�E���8�xp|,��AQ�,`4N
q�@(W3�T0 k� �;�;U2d   2$ !  ��H   � <���x
E��E���4�po|,��AQ�,P,M
q�@,W3�T0 k� � A�AU2d   2$ !  ��H    � <���t
E�w�E���0�lo|,��AQ�+P$M
q�@,X3�T0 k� ��F� FU2d   2$ !  ��H    � <���lE�s�E�{�,�dn|,�߻AQ�+PL
q�@,X3�T0 k� ��I��IU2d   2$ !  ��H    � <���dE�o�E�s�,�`n|,�ۻAQ�+PK
q�@,X"s�T0 k� ��K��KU2d   2$ !  ��H    � <���\E�g�E�k�(�Xn|,�ӺAQ�+PK
q�@0Y"s�T0 k� ��M��MU2d   2$ !  ��H    � <���TD1c�E�c�$�Tm|,�ϺAQ�+PJ
q�@0Y"s�T0 k� ��M��MU2d   2$ !  ��H    � <���LD1[�E�[� �Lm|,�˹AQ�+_�I
q�@0Y"s�T0 k� ��M��MU2d   2$ !  ��H    � <���DD1W�E�W� �Hm|,�ǹAQ�+_�I
q�@0Z"s�T0 k� ��N��NU2d   2$ !  ��H    � <���<D1O�E�L �@l|,���AQ�+_�H
q�@4Z"s�T0 k� ��N��NU2d   2$ !  ��H    � <���4D1G�E�D�<l|,���AQ�+_�G
q�@4["s�T0 k� ��M��MU2d   2$ !  ��H    � <���,D1C�D�<�4k|,���AQ�+O�G
q�@4["s�T0 k� ��P��PU2d   2$ !  ��H    � <���$D1;�D�8�0k|,���AQ�+O�F
q�@4["s�T0 k� ��Q��QU2d   2$ !  ��H    � <���D17�D�0�,k|,���AQ�+O�F
q�@8\"s�T0 k� ��R��RU2d   2$ !  ��H    � <���D1/�D�(�$j|,���AQ�+O�E
q�@8\"s�T0 k� ��R��RU2d   2$ !  ��H    � <���E�+�D�$� j|,���AQ�*O�E
q�@8\3�T0 k� ��S��SU2d   2$ !  ��H    � <���E�#�D�	�j|,���AQ�*O�E
q�@8]3�T0 k� ��T��TU2d   2$ !  ��H    � <����E��D��i|,���AQ�*O�D
q�@<]3�T0 k� ��S��SU2d   2$ !  ��H    � <����E��D��i|,���AQ�*O�D
q�@<]3�T0 k� �|S��SU2d   2$ !  ��H    � <����E��D� �i|,���AQx*O�D
q�@<^3�T0 k� �tS�xSU2d   2$ !  ��H    � <����E��D� ��h|,���AQt*ϐD
q�@<^3�T0 k� �pR�tRU2d   2$ !  ��H    � <����E��D�  �� h|,���AQp*ψC
q�@<^3�T0 k� �hQ�lQU2d   2$ !  ��H    � <����E���D�� ���h|,���AQl*�|C
q�@@^3�T0 k� �`P�dPU2d   2$ !  ��H    � <����E���D�� ���h|,���AQh*�tC
q�@@_3�T0 k� �XP�\PU2d   2$ !  ��H    � <����E���D�� ���g|,��AQd*�lC
q�@@_3�T0 k� �PP�TPU2d   2$ !  ��H    � <����E���D�� ���g|,�{�AQ`*�dC
q�@@_3�T0 k� �HL�LLU2d   2$ !  ��H    � <����E���D�� ���g|,�w�AQX*�\C
q�@@`"��T0 k� �<I�@IU2d   2$ !  ��H    � <����E���D�� ���f|,�s�AQT*�TC
q�@D`"��T0 k� �4G�8GU2d   2$ !  ��H   � <����E���D�� ���f|,�o�AQP*�LC
q�@D`"��T0 k� �,E�0EU2d   2$ !  ��H    � <����D���D�� ���f|,�k�AQL*�@C
q�@D`"��T0 k� �$D�(DU2d   2$ !  ��H    � <����D���D�� ���f|,�g�AQH*�8C
q�@Da"��T0 k� �C� CU2d   2$ !  ��H    � <����D���D��! ���e|,�c�AQD*�0C
q�@Da"��T0 k� �B�BU2d   2$ !  ��H    � <����D���D��# ���e|,�_�AQ@)�(C
q�@Da"��T0 k� �A�AU2d   2$ !  ��H   � <����D���D��% ���e|,�[�AQ<)� C
q�@Ha"��T0 k� � A�AU2d   2$ !  ��H    � <����D���D��& ���e|,�[�AQ8)�C
q�@Hb"��T0 k� ��A��AU2d   2$ !  ��H    � <����D���D��( ���d|,�W�AQ4)�C
q|@Hb"��T0 k� ��<��<U2d   2$ !  ��H    � <��ѼD���D��* ���d|,�S�AQ4)�C
qx@Hb"��T0 k� ��8��8U2d   2$ !  ��H    � <���D���D��, ���d|,�O�AQ0)��C
qt@Hb3�T0 k� ��5��5U2d   2$ !  ��H    � <���D���D��.����d|,�K�AQ,)��C
qt@Hc3�T0 k� ��3��3U2d   2$ !  ��H    � <���D���E��0����d|,�K�AQ()��C
qp@Lc3�T0 k� ��1��1U2d   2$ !  ��H    � <��� D���E��2����c|,�G�AQ$)��B
ql@Lc3�T0 k� ��1��1U2d   2$ !  ��H    � <��� D���E��3����c!�,�C�AQ )��B
qh@Lc3�T0 k� ��2��2U2d   2$ !  ��H    � <���!D���E��5����c!�,�?�AQ)��B
qd@Lc3�T0 k� ��2��2U2d   2$ !  ��H    � <���!D��E��7����c!�,�?�AQ)��B
q`@Ld3�T0 k� ��2��2U2d   2$ !  ��H    � <���"D�{�E��9����b!�,�;�AQ)��A
q\@Ld3�T0 k� ��1��1U2d   2$ !  ��H    � <���"D�w�E��;����b!�,�7�AQ)��A
q\@Ld3�T0 k� ��1��1U2d   2$ !  ��H    � <���#D�s�E��=����b!�,�3�AQ)��A
qX@Pd3�T0 k� ��1��1U2d   2$ !  ��H    � <���#D�k�E��?����b!�,�3�AQ)��@
qT@Pd3�T0 k� �|0��0U2d   2$ !  ��H    � <���#D�g�F�A����b!�,�/�AQ)��@
qP@Pe3�T0 k� �t0�x0U2d   2$ !  ��H    � <���#D�c�F|C����a!�,�+�AQ).�@
qL@Pe3�T0 k� �h1�l1U2d   2$ !  ��H    � <���$D�_�F|E����a!�,�+�AQ).�?
qH@Pe3�T0 k� �`1�d1U2d   2$ !  ��H    � <���$D�[�FxG����a!�,�'�AQ ).�?
qD@Pe3�T0 k� �X2�\2U2d   2$ !  ��H    � <���|%D�W�FtI����a|,�#�AQ ).�>
qD@Pe3�T0 k� �P1�T1U2d   2$ !  ��H    � <���x%D�S�FpK����a|,�#�AP�).x>
q@@Pf3�T0 k� �H1�L1U2d   2$ !  ��H    � <��Ap&D�O�FpM����a|,��AP�).p>
q<@Tf3�T0 k� �@1�D1U2d   2$ !  ��H    � <��Al'D�K�FlO����`|,��AP�)>h=
q8@Tf3�T0 k� �80�<0U2d   2$ !  ��H    � <��Ad'D�G�FlQ����`|,��AP�)>`=
q4@Tf3�T0 k� �00�40U2d   2$ !  ��H    � <��A`(D�C�FhS��	�|`|,��AP�(>X=
q4@Tf3�T0 k� �(0�,0U2d   2$ !  ��H    � <��AX)D�?�FhU��	�|`|,��AP�(>P<
q0@Tf3�T0 k� � /�$/U2d   2$ !  ��H    � <��AT*D�;�FdW��
�x`|,��AP�(>L<
q,@Tg3�T0 k� �/�/U2d   2$ !  ��H    � <��AL*D�7�FdY��
�t`|,��AP�(ND<
q(@Tg3�T0 k� �/�/U2d   2$ !  ��H    � <���H+D�3�E�d[���t_|,��AP�(N<;
q(@Tg3�T0 k� �.�.U2d   2$ !  ��H    � <���@,D�/�E�d]���p_|,��AP�(N4;
q$@Xg3�T0 k� �.�.U2d   2$ !  ��H    � <���<-D�+�E�`_���p_!�,��AP�(N0;
q @Xg3�T0 k� ��.� .U2d   2$ !  ��H    � <���4.D�'�E�`a���l_!�,��AP�(N(;
q @Xg3�T0 k� ��.��.U2d   2$ !  ��H    � <���,/D�#�E�`b���h_!�,��AP�(N :
q@Xh3�T0 k� ��.��.U2d   2$ !  ��H    � <���(/D��E�`d���h_!�,��AP�(N:
q@Xh3�T0 k� ��.��.U2d   2$ !  ��H    � <��� 0D��E�`f���d_!�,��AP�(N:
q@Xh3�T0 k� ��.��.U2d   2$ !  ��H    � <���1D��E�`h�|�d^!�,��AP�(N9
q@Xh3�T0 k� ��-��-U2d   2$ !  ��H    � <���2D��E�dj�x�`^!�,���AP�(N9
q@Xh3�T0 k� ��-��-U2d   2$ !  ��H    � <���2D��E�dk�t�`^!�,���AP�(N9
q@Xh3�T0 k� ��-��-U2d   2$ !  ��H    � <���3D��E�dm�l�\^!�,���AP�(M�9
q@Xh3�T0 k� ��,��,U2d   2$ !  ��H    � <���4D��E�do�h�X^!�,���AP�(M�8
q@\i3�T0 k� ��,��,U2d   2$ !  ��H    � <���5D��E�hp�d>X^!�,���AP�(M�8
q@\i3�T0 k� ��,��,U2d   2$ !  ��H    � <���5D��E�hr�`>T^|,���AP�(M�8
q@\i3�T0 k� ��,��,U2d   2$ !  ��H    � <���6D��E�hs�X>T]|,��AP�(=�7
q@\i3�T0 k� ��+��+U2d   2$ !  ��H    � <���7D��E�lu�T>P]|,��AP�(=�7
q @\i3�T0 k� ��+��+U2d   2$ !  ��H    � <���7D���E�lv@P>P]|,��AP�(=�7
q @\i3�T0 k� ��+��+U2d   2$ !  ��H    � <���8D���E�px@H>L]|,��AP�(=�7
p�@\i3�T0 k� ��+��+U2d   2$ !  ��H    � <���9D���E�py@D>L]|,��AP�(=�7
p�@\i3�T0 k� ��*��*U2d   2$ !  ��H    � <���9D��E�tz@@>H]|,��AP�(-�6
p�@\j3�T0 k� ��*��*U2d   2$ !  ��H    � <���:D��E�t{@8>H]|,��AP�(-�6
p�@\j3�T0 k� ��*��*U2d   2$ !  ��H    � <���:D��E�x|@4>H]|,��AP�(-�6
p�@\j3�T0 k� ��*��*U2d   2$ !  ��H    � <���;D��E�|}@, >D]|,��AP�(-�6
p�@`j3�T0 k� ��)��)U2d   2$ !  ��H    � <���;D��E�|~@(!>D\|,��AP�(-�5
p�@`j3�T0 k� �x(�|(U2d   2$ ! �H    � <���<D��
E��@ ">@\|,��AP�(�5
p�@`j3�T0 k� �d'�h'U2d   2$ ! ��O    � <�� �=D��E���@$>@\|,��AP�(�5
p�@`j3�T0 k� �T%�X%U2d   2$ ! ��O    � <�� �=L_�E���0%N<\|,��AP�(�5
p�@`j3�T0 k� �@$�D$U2d   2$ ! ��O    � <�� �>L_�E��0&N<\|,�ߤAP�(�5
p�@`k3�T0 k� �0#�4#U2d   2$ ! ��O    � <�� �>L_�E��0(N<\|,�ߣAP�(�4
p�@`k3�T0 k� �!� !U2d   2$ ! ��O    � <�� �?L_�E��0)N8\|,�ߣAP�(�4
p�@`k3�T0 k� � � U2d   2$ ! ��O    � <�� �?L_�CO�~0 +N8\|,�ۣAP�(�4
p�@`k3�T0 k� ����U2d   2$ ! ��O    � <�� �@L_�CO�~?�,N4\|,�ۣAP�'�4
p�@`k3�T0 k� ����U2d   2$ ! ��O    � <�� �@L_�CO�}?�.N4\|,�ۣAP�'�4
p�@`k3�T0 k� ����U2d   2$ ! ��O   � <�� �AL_�CO�}?�/N4[|,�ףAP�'�3
p�@`k3�T0 k� ����U2d   2$ ! ��O   � <�� �AL_�CO�|?�1N0[|,�ףAP�'�3
p�@`k3�T0 k� ����U2d   2$ ! ��O    � <�� |BL_�CO�{?�2N0[|,�ףAP�'�3
p�@`k3�T0 k� ����U2d   2$ ! ��O    � <�� xBLo�Kߘ{O�4N,[|,�ӣAP�'�3
p�@dk3�T0 k� ����U2d   2$ ! ��O    � <�� tBLo�KߜzO�5N,[|,�ӢAP�'|3
p�@dl3�T0 k� �|��U2d   2$ ! ��O    � <�� pCLo� KߜyO�7N,[|,�ӢAP�'x3
p�@dl3�T0 k� �l�pU2d   2$ ! ��O    � <�� lCLo�!KߠyO�8N([|,�ϢAP�'t2
p�@dl3�T0 k� �X�\U2d   2$ ! ��O    � <�� hDLo�#KߠxO�:N([|,�ϢAP�'t2
p�@dl3�T0 k� �H�LU2d   2$ ! ��O    � <�� dDLo�$Kߤx?�;N([|,�ϢAP�'p2
p�@dl3�T0 k� �4�8U2d   2$ ! $�O    � <�� `ELo�%Kߤw?�=N$[|,�ϢAP�'l2
p�@dl3�T0 k� <4�8U2d   2$ ! ��O    � <�� XELo�&Kߨv?�?N$[|,�ˢAP�'h2
p�@dl3�T0 k� <4�8U2d   2$ ! ��O    � <�� TELo�(Kߨv?�@N$[|,�ˢAP�'d2
p�@dl3�T0 k� <8�<U2d   2$ ! ��O   � <�� PFLo�)K߬u?�BN$[|,�ˢAP�'`1
p�@dl3�T0 k� <8�<U2d   2$ ! ��O   � <�� PFLo�*K߬u?�DN Z|,�ǡAP�'\1
p�@dl3�T0 k� <8�<U2d   2$ ! ��O   � <�� LGLo�+K߬t?�EN Z|,�ǡAP�'\1
p�@dl3�T0 k� �8�<U2d   2$ ! ��O   � <�� HGLo�-K߰t?�GN Z|,�ǡAP�'X1
p�@dl3�T0 k� �8�<U2d   2$ ! ��O    � <�� DGLo�.K߰s/�INZ|,�ǡAP�'T1
p�@dm3�T0 k� �8�<U2d   2$ ! ��O    � <�� @HLo�/K�s/�JNZ|,�áAP�'�P1
p�@dm3�T0 k� �<�@U2d   2$ ! ��O    � <�� <HLo�0K�r/�LNZ|,�áAP�'�L1
p�@dm3�T0 k� �<�@U2d   2$ ! ��O    � <�� 8HLo�1K�r/�NNZ|,�áAP�'�L0
p�@hm3�T0 k� �<�@U2d   2$ ! ��O    � <��                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��C� ]�#`#_ � �� Kb
      
	  ����     Kb
���                        Z���         .      ���   0
 
          t��  Z Z    � ��     t�c �     D9            P  Z��          ��     ��� 0
% 	           ^)�    
	   ���4     ^)����4                   	 Z���        ��     ���   8

           b�+   � �    ��h�     b�+��h�           	           	 Z��          � �     ���  8          W�Y     
   .�w@�     W�Y�wCv      ��               Z��          �@     ���   P
	
          1�  ��
	    B��     1���                             �^              �  ���    P             ��A9    	     V��+"    ��A9��-       ��                	 i =         �     ��@   8	 

          '*(         j ��     '*( �}      ��                   o <         �p     ��@   0

!           )��   �	    ~�&�[     )���&�      �m                  ��          �     ��H   H	
          ~#  � �
      � �     ~#  '      ��                      �         	 ڠ
`     ��P   (
          r��  `      � ��B     r�� ��B                        
 A �         
  �P     ��@   X           � ��
      � ��3     � ��3                                ���                ��@   0

 
2
 
                 ��      �                                                                           �                               ��        ���          ��                                                                 �                          z�g  ��        ��(�\     z�r�(�i    ���                    x                j  �   �   �                          z    ��        ��)       z  �)           "                                                 �                         �� �����w��� �&  � ����(�)  
 	              
   �   �h� ���N       �d �c@ �d 0d@ �� d� ��  d� ˤ _� �� `  �� �`� �� a� � a� �$ b  �D b  �d b@���X � �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0� ���� ����� ����� � � �m@ � n@ ބ �r@���� � |  d� |D  e  N e@ GD `j� H 0k� Hd k� H� l  9$ �e� :$  f� :d g  JD �m@ KD 0n@ K�  n� :� `[� ;D  \� ;� \� ;� \� ;� `o� <� p� <� p� <�  p� K� �`� L�  a� #� `^@ $d _  
�\ U� 
�� V  
�\ V  
�\ V� 
�� V� 
�| W  
�\ W� 
�� W� 
�\ W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������� <��   ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"     �j
��   �
� �  �  
�  5��  ��     ��n  �    W��  ��     ��w       )��  ��     ��&          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �O      ��T ��        � �T ��        �        ��        �        ��        �   �     q� 
��        ��                         ���    ����                                     �                ����            ����%��   <����               25 Terry Yake rson y   4:21                                                                        1  1     �C
2�C
� �SC.k C6 �B� �C �C" � C% �	C& �
K � K �J�2 � J�2 � J�* � J�" �kj � � kr � �c� � �c� � � c� �u"�u "�e"�e*� q *Ht �  *GtI *2tI *2tA )�t �)�t � *Jt) * |A )�tA "*FdA )�t9$*lA %*FdI *2t9  *>| � (*Et) )*Pd)***|9+*lA ,*FdI *2tA )�t � /*Jt)0* |A )�tA 2*FdA )�tA )�t!5)�tY  *Jt* )�t8"|- )�t � :*Gd � ;*Et<"|0 )�t � >*Et "|                                                                                                                                                                                                                         h� R         �     @ 
        �     a P E f  ��                   	 
�������������������������������������� ���������	�
��������                                                                                          ��    �"�� ��������������������������������������������������������   �4, :� 6 �@"�@���@�@��A)���������                                                                                                                                                                                                                                                                                                                    �                                                                                                                                                                                                                                                    d    7      �  D�J    	  $m                             ������������������������������������������������������                                                                               
                                                           �     �      �        �        �  �          	  
 	 
 	 	 ��������������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� �           x                        #    � �   R�J    
  �                             ������������������������������������������������������                                                                         	                                                                  �� 0        �      �      �  �              	 	 
  	 	 	 ����� ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� �������������                                                                                                                                                                                                                                                                                                                               �             


           �   }�                                                                          N�               ����������������������������   ����������������   ������������  *��������������������������������������ww�ww333wwwwwwww�ww�ww�ww�ww333wwww N @ 0 
              	 
                 � -/� �c@                                                                                                                                                                                                                                                                                   E)n1n  	n                    b                  l            m                                                                                                                                                                                                                                                                                                                                                                                                          
 �  � ��  � ��  � (��  �  ��  EZm�  �N ��H�r����������������h�����W���������*         :  ���> : ~��        
 	 
�   & AG� �   R              �r�                                                                                                                                                                                                                                                                                                                                      p B J   �      ��                !��                                                                                                                                                                                                                            Y   �� �� ����      �� B 	     ��������������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ������ ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� �������������   ��       ���������������������������������������������������f��ff�fff�ff���������l�ff�ffffl��ff˼fllf������l��̼�ʗ���˹�ffjz�fkyl�l��fƨ�����������������������̼��̉������������������������������f���f�fff�ff�ffl�ff�flfl�l��xl�wwl���l̻�����˺��fl����l�xx��w��̻���l�f�f�ƻ�fl�����ffl�ffffffff���f���̚���ffflffflfffffffffflfffff������������������������l���l������f����������������������������l��lf��f�fff�f��l˪���ww��w�����flflffffffff�̼̙��fww��w��fx�̻�llffff�ffff���fl���f�l�l�˶����fffl��fflfll����ff��ff��lfl�lf��l���l�����������l�������l�������ʼ�j˚��̩��ʨ��ɘ���xxxȈ��ɉ�x���̇�̺������www��ww��xw���x��xk�����������wx��������������x����l�ƈ��Ƈ���w��Ɨ��̩z�̩yf̪�f�������������������������������̙i���ɖ�yɌ��ˌȉ̚ə̩���ə��Ɉ����x�̹x�̹�����������ƺ�������������������ˈ������˙������̫��̺�������˪�������������̸��̗�����̇��̇�����������������������̈���xx����x���w���ɉ��̨���k���̛̻�������������l��Ʀl�Ɗl�l���̻�lk��̺�f̩�l��f�ɫ�ˉ�lɊ�˙���ʚ���˙�˫̼���ɬ�̚��̼�����̼���̬������̼�����˻������������f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff���m�    E      5   �  z                       B     �   �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �r@  �    � �N ^$   �̞   8  ��  ��   �   �   ��Ҝ     �f ��     �� p���� ���� p���� �$��   `d     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@     | 
f� ��  | 
f� �$ ^$   l c@ �d �� c@ �d �$ & �  ��&  �      �  ��   ���� e�����   g���  �     f ^�         �� � <            ��D$���2�������J���p���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            "! "   "      ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "!  " ! " ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       "! "   "      ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   �   ��  � � ��      �    �     ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                              	�    �     �                                                                                                                                                                                                 �  �  ��  8�  5I  5U  3U  DT  EZ UJ T� �J� ����+�""""�""//��          ��wɪ�pɪ��ɪ��̙�н��н̽Ѝɚݣ��"�<̲�;���0"�0  ="  ""  "/  /�� ���  �����                               �� �� �� ���          �.���       �  �      �  ��  �  ��  �              �                                   ����  �   �             ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                       �   ���                            �   �                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw     �  �  ��  �   �   �                         ���                                                                                                                                                                            �� ̽ ̽��۽ }�  wz  � ��������ɜ���̚��̸ ��  ��  �  �  T�  T�  H� �E �E �D�[ ˻  ˸  ��  
� ,"�"" �"  �"              "   *�  ��� ��� �ة��ڋ�̽� ��  ��  ̻� ̻� ��� ��@ ��@ DD0 T30 B3� ��  ��  ��  
� +� �"" �"� �" ��� ����  ��          ���    �                       
 "� ""� ""� "                       �                             ���                         �  ��                    �����                                  �  �˰ ��� �wp ���                                                                                                                                                                 �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��        �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                  �       �                        �   ��  ���  � �    �                                                                                                                                            �   �  �  �� �� �� �� T� EJ  4T  3E  E   4   �         �   �   �               �̚���ɀ��̰��� ��� �ɘ���˸������⌄@���D�J�ЉZ�یT��ۻ� ��� ͹� ͹� ؛��۝��������۹�"۲                    �   �   �   �   ��  ��  Ș����� �  �    �  �           �      �   ��   �  �  ��  �   �                     �� �� �� �� �݉���̙�  ���                              �������  �                     �  �   �  �  ��  �  ��  �                                                                                                                                                                                                    �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                �   ���                                                                                                                                                                                                      	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                        �          �   � � �  ��� ��  �                       �   �                      �������  ���    �              �  �� ��  �    � ���                                                                                                                                                                                              �  ��  ��  ��  �  �w 
�w Ț� ̹� ��� ��� �ͼ �� �� 
��  �-  "  3"  3$ 33 �33 �30*� ""  ""��"/����   �              �   �   �   �   ڀ  z�  ��� ��� ��� ��ɠ̽��̸���������ܼ���ۉ�����4EX EU� EU� U� TX K�  ��  �� �� " �"" "  �"/  ���            �  �  �" �.�� "            �   �   �  �  �  �           �   ��  �   ��  �                    �� ��� ��� ����                            �                               � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                     �  �  �  �  �� 
�w ��p������˚��̸���̽��̍̽��̽�����̘�������J�ST�C UJ� Z�  J�  ۼ �� ʨ "�� "+� "" �""   ���   ��  ��  �p  }`  g`  w                   �   �   �   �   �   �   ""  "   ". 0  �@  �   �   �               "�  "/  ����  �       �       �        ���                    ������������                        �                         �   �                      �������  ���    �                    ��  ��  ���                    � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         �  ��� ��� }�� wݪ �� 	�� �� �ͼ ��� ��� ̘� �ͻ +���"�8"8  8� �� �U��EU��3 ̻�"̰""�" ��" �"                             �   ��� �˹��˚���ڍ�̽���ͽ��ͽ���ݼ��л�� ��D �UT EUT UU0 C3  2"  ""  -�  ��  ��  �   � ��"/ �" � ���    �        �   ��  ��  ��  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ���                 ��                                                                                                                                                                                             �� ̻ ��˛��  �� �˚̻���ۚ����I���䘼�^���^�٘�:�^�� ^�� D�( �) �) �) ��) ˹� ț�+��,��,����  �𫝝 ��� �ɍ ��ݨ��ډ�݊�� ��D@ �D�  J�� ݩ� ��� �ۻ �ک �ڹ�ɻ��̸���������� ����������            �   ��  ��  ��  ��  ��                                          �� ��� ��� ��  �                         �   �                    �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��   �  �   
�  �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                             "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwww""""wwwwwwwGwqGwGwDGwG""""wwwwwwqAqwAwG""""wwwwwwwwDDwwwwwwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwqDDDG""""wwwwwqqADAqq""""wwwwwwqwwwqwqwq""""wwwwqDDDwGq"""$www4ww4Gw4DGw4www4ww4wwwwwwwwwwtwww333DDDGwGGwqwDDwtwwww3333DDDDwGtqGwADqDGwDwwww3333DDDDwwqwwwwDwwDGwwwwww3333DDDDADAGqGqtGwDwwww3333DDDDGqGqGqGqtGwDwwww3333DDDDGqqqwwtDDwwww3333DDDDDDqwqqqwAwtDGwwww3333DDDDwqwqwGqDDGwwwww3333DDDDDGwAwwwwDDtDwwww3333DDDDww4Gw4Gw4Gw4Dww4www43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
2�C
� �SC.k C6 �B� �C �C" � C% �	C& �
K � K �J�2 � J�2 � J�* � J�" �kj � � kr � �c� � �c� � � c� �u"�u "�e"�e*� q *Ht �  *GtI *2tI *2tA )�t �)�t � *Jt) * |A )�tA "*FdA )�t9$*lA %*FdI *2t9  *>| � (*Et) )*Pd)***|9+*lA ,*FdI *2tA )�t � /*Jt)0* |A )�tA 2*FdA )�tA )�t!5)�tY  *Jt* )�t8"|- )�t � :*Gd � ;*Et<"|0 )�t � >*Et "|3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.����������������������������������������� ��=�K�X�X�_��B�G�Q�K� � � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������6�+� � ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� ��#�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                