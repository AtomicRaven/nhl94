GST@�                                                           �t�                                                      U���      �  >      
      ����e J���J�������̸��`�������        �g     #    ����                                d8<n    �  ?     ����  �
fD�
�L���"����D"� j   " B   J  jF�"     "�j  " ���
��
�"    B�jl �   B ��
  ��                                                                              ����������������������������������       ��    =b 0Qb 4 114  4c  c  c        	 
      	   
       ��G �� � ( �(                 nn 
)1         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                  +       �   @  &   }   �                                                                                 '      
)n1n  �    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E + �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��Z C�A���BM�0�o��L�ތNA�����l��Z3��T0 k� ���#[P "�2't �8t B ��_    ����8��[ C�A���BM�0�o��L�ތNL<����l��Z3��T0 k� ���#[P "�2't �8t B ��_    ����8��[ C�A���BM�0�o��L�ތNL<����l��Z3��T0 k� ���#[P "�2't �8t B ��_    ����8��[ C�A���BM�0�o��L�ތOL<����l��Z3��T0 k� ���#kP "�2't �8t B ��_    ����8��[ C�A���BM�0�o��L�ތOL<����l��Z3��T0 k� ���#kP "�2't �8t B ��_    ����8��\ G�A���BM�0�o��L�ސOL<����\��Z3��T0 k� ���#kP "�2't �8t B ��_    ����8��\ G�A���BM�0�o��L� ��OL<����\��Z3��T0 k� ���#kP "�2't �8t B ��_    ����8��\ G�A���BM�0�o��L� ��PL<����\��Z3��T0 k� ���#kP "�2't �8t B ��_    ����8��\ G�A���BM�0�o��L� ��PL<����\��Z3��T0 k� ���#{P "�2't �8t B ��_    ����8��] G�A���BM�0�o��L� ��PL<����\��Z3��T0 k� ���#{P "�2't �8t B ��_    ����8��] G�A���BM�0�o��L� ��PL<����\��Z3��T0 k� ���#{P "�2't �8t B ��_    ����8��] G�A���BM�0�o��L� ��QL<�������Z3��T0 k� ���#{P "�2't �8t B ��_    ����8��] G�A���BM�0�o��L� ��QL<�������Z3��T0 k� ���#{P "�2't �8t B ��_    ����8��^ G�A���BM�0�o��L� ��QL<�������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��^ G�A���BM�0�o��L� ��QL<�������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��^ G�A���BM�0�o��L� ��RLL�������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��^ G�A���BM�0�o��L� ��RLL�������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��^ G�A���BM�0�o��L� ��RLL�������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��_ G�A���BM�0�o��L� ��RLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��_ G�A���BM�0�o��L� ��SLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��_ G�A���BM�0�o��L� ��SLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��_ G�A���BM�0�o��L� ��SLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��` G�A���BM�0�o��L� ��SLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��` G�A���BM�0�o��L� ��SLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��` G�A���BM�0�o��L� ��TLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��` G�A���BM�0�o��L� ��TLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��` G�A���BM�0�o��L� ��TLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��a G�A���BM�0�o��L� ��TLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��a G�A���BM�0�o��L� ��TLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��a G�A���BM�0�o��L� ��ULL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��a G�A���BM�0�o��L� ��ULL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��a G�A���BM�0�o��L� ��ULL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��a G�A���BM�0�o��L� ��ULL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��b G�A���BM�0�o��L�� ��ULL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��b G�A���BM�0�o��L�� ��VLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��b G�A���BM�0�o��L�� ��VLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��b G�A���BM�0�o��L�� ��VLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��b G�A���BM�0�o��L�� ��VLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��b G�A���BM�0�o��L�� ��VLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��c G�A���BM�0�k��L�� ��VLL������Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��c G�A���BM�0�k��L�� ��WLL�,�����Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��c G�A���BM�0�k��L�� ��WLL�,�����Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��c G�A���BM�0�k��L�� ��WLL�,�����Z3��T0 k� ���#�P "�2't �8t B ��_    ����8�c G�A���BM�0�k��L�� ��WLL�,�����Z3��T0 k� ���$P "�2't �8t B ��_    ����8�c G�A���BM�0�g��L�� ��WLL�,�����Z3��T0 k� ���$P "�2't �8t B ��_    ����8�c G�A���BM�0�g��L�� ��WLL�,�����Z3��T0 k� ���$P "�2't �8t B ��_    ����8�d G�A���BM�0�g��L�� ��WLL�,�����Z3��T0 k� ���$P "�2't �8t B ��_    ����8�d G�A���BM�0�g��L�� ��XLL�,�����Z3��T0 k� ���$P "�2't �8t B ��_    ����8�d G�A���BM�0�g��L�� ��XLL� l�����Z3��T0 k� ���#;P "�2't �8t B ��_    ����8�d G�A���BM�0�g��L�� ��XLL� l�����Z3��T0 k� ���#;P "�2't �8t B ��_    ����8�d G�A���BM�0�c��L�� ��XLL� l�����Z3��T0 k� ���#;P "�2't �8t B ��_    ����8�d G�A���BM�0�c��L�� ��XLL� l�����Z3��T0 k� ���#;P "�2't �8t B ��_    ����8��d G�A���BM�0�c��L�� ��XLL� l�����Z3��T0 k� ���#;P "�2't �8t B ��_    ����8��e G�A���BM�0�c��L�� ��XLL�������Z3��T0 k� ���#KP "�2't �8t B ��_    ����8��e G�A���BM�0�c��L�� ��YLL�������Z3��T0 k� ���#KP "�2't �8t B ��_    ����8��e G�A���BM�0�c��L�� ��YLL�������Z3��T0 k� ���#KP "�2't �8t B ��_    ����8��e G�A���BM�0�_��L�� ��YL<�������Z3��T0 k� ���#KP "�2't �8t B ��_    ����8��e G�A���BM�0�_��L�� ��YL<�������Z3��T0 k� ���#KP "�2't �8t B ��_    ����8��e G�A���BM�0�_��L�� ��YL<�������Z3��T0 k� ���#kP "�2't �8t B ��_    ����8��e G�A���BM�0�_��L�� ��YL<�������Z3��T0 k� ���#kP "�2't �8t B ��_    ����8��e G�A���BM�0�_��L�� ��YL<�������Z3��T0 k� ���#kP "�2't �8t B ��_    ����8N�e G�A���BM�0�_��L�� ��YL<�������Z3��T0 k� ���#kP "�2't �8t B ��_    ����8N�f G�A���BM�0�_��L�� ��ZA��������Z3��T0 k� ���#kP "�2't �8t B ��_    ����8N�f G�A���BM�0�[��L�� ��ZA��̻����Z3��T0 k� ���#{P "�2't �8t B ��_    ����8N�f G�A���BM�0�[��L�� ��ZA��̻����Z3��T0 k� ���#{P "�2't �8t B ��_    ����8��2 ���@� @o8# o;�|  �+��(2P�<  ����#Z3� T0 k� �  � "�2't �8t B  ��/    �   2��2 ���@� @o8# o;�|  �+��(2AP<  ����#Z3� T0 k� �  � "�2't �8t B  /�/    �   6��2 ���@� @o8# o;�|  �+��(2AP<  ����#Z3� T0 k� �$ �( "�2't �8t B  ��/    �   :��2 ���B�� @o8# o;�|  �+��(2A�<  ����#Z3� T0 k� �, �0 "�2't �8t B  ��/    �   >��2 ���B�� @o8# o;�|  +��(2A�< �����#Z3� T0 k� �4 �8 "�2't �8t B ��/    �   B��2 ���B�� @o8# o;�|   +��(2A�< �����#Z3� T0 k� �@ �D "�2't �8t B ��/    �   F��2 ���B�� @o8# o;�|   +��(2A�< �����#Z3� T0 k� �H �L "�2't �8t B ��/    �   I��1 ���B�� @o8# o;�|   +��(1A�< �����#Z3� T0 k� �P �T "�2't �8t B ��/    �   L��1_��B�� @8# o;�|$  +��(1P�< �����#Z3� T0 k� �X �\ "�2't �8t B ��/    �   O��1_��B�� @8# �;�|$ P+��(1P�< �����#Z3� T0 k� �` �d "�2't �8t B ��/    �   R��0_��B�� @8# �;�|$ P+��(0P�< �����#Z3� T0 k� �l �p "�2't �8t B ��/    �   U��0_��B�� @8# �;�|$ P+��(0P�< �����#Z3� T0 k� �t �x "�2't �8t B ��/    �   X��0_��B�� @8# �;�|( P+��(/P�@ ���@�#Z3� T0 k� �| �� "�2't �8t B ��/    �   [��/���B�� BO8# �;�|( P+��(/P�D ���@�#Z3� T0 k� �� �� "�2't �8t B ��/    �   ^��.���B�� BO8#O;�|( �+��(.P�D 0��@�#Z3� T0 k� �� �� "�2't �8t B ��/    �   a��.���B�� BO8#O;�|( �+��(-P�H 0��@�#Z3� T0 k� � �� "�2't �8t B ��/    �   d�-���B�  BO8#O;�|( �+��(,P�L 0��@�#Z3� T0 k� � �� "�2't �8t B  ��/    �   d�,���B� BO8#O;�|( �+��(,P�L 0����#Z3� T0 k� �����"�2't �8t B  ��)    �   d�,���B� A�8#O;�|( �+��(+P�P 0����#Z3� T0 k� �����"�2't �8t B  ��)    �   c�+���B� A�8#�;�|( �+��(*P�T 0����#Z3� T0 k� �����"�2't �8t B  ��)    �   b�*���B� A�8#�;�|( �+��()P�T 0����"Z3� T0 k� �����"�2't �8t B  /�)    �   a�)���B� A�8#�;�|( �+��((P�X 0����"Z3� T0 k� �����"�2't �8t B  ��)    �   `�)���B� A�8#�;�|( �+� ('P�X  ����"Z3� T0 k� �����"�2't �8t B  ��)    �   _�(���B� A�8#�;�|( �+� (&P�\  ����"Z3� T0 k� �����"�2't �8t B  ��)    �   ^�'���B� A�8#�7�|( �+� ($P�`  ����!Z3� T0 k� �����"�2't �8t B  ��)    �   ]�&���B� A�8$�7�|( �+� (#P�`  ����!Z3� T0 k� �����"�2't �8t B  ��)    �   \��%���B� A�8$�7�|( �/� ("P�d  ����!Z3� T0 k� �����"�2't �8t B  ��)    �   [��$���B� A�8$�7�|( �/��,!Epd  �� � Z3� T0 k� �����"�2't �8t B  ��)    �   Z��#O��B� A�8$�3�|( �/��, Eph  �� � Z3� T0 k� �����"�2't �8t B  ��)    �   Y��!O��B�  A�4$�3�|( p/��,Epl �� �Z3� T0 k� �����"�2't �8t B  ��)    �   X� O��B�$ Eo4%�/�|( p/��,Epl �� �Z3� T0 k� �����"�2't �8t B  ��)    �   W�O��B�( Eo4%�/�|( p/�	�0E`l����Z3� T0 k� �����"�2't �8t B  ��)    �   W����B�, Eo0%�+�|( p/�	�0E`l����Z3� T0 k� �����"�2't �8t B  ��)    �   W����B�, Eo,&�'�|( `/�	�8E`p  ����Z3� T0 k� ������"�2't �8t B  ��)    �   W����B�0 E_,&�'�|( `/�	�8E`t  ����Z3� T0 k� ������"�2't �8t B  ��)    �   W����B�4 E_('�#�|( `/�
 <D0t  ����Z3� T0 k� ������"�2't �8t B  ��)    �   W����B�4 E_('��|( `3�
 @D0x  ����Z3� T0 k� ������"�2't �8t B  ��)    �   W����B�8 E_$'��|( `3�
 DD0x  ����Z3� T0 k� ����"�2't �8t B  ��)    �   W  ���B�8 E_(��|( `3�
 HD0|  ����Z3� T0 k� ����"�2't �8t B  ��)    �   W ���B�8 EO(��|( `3� LD0|  ����Z3� T0 k� ����"�2't �8t B  ��)    �   W ���B�< EO(��|( P7� PD0|  ����Z3� T0 k� ����"�2't �8t B  ��)    �   W ���B�@ EO)��|( P7� PD0�  ����Z3� T0 k� ���#�"�2't �8t B  ��)    �   W ���B�@ EO)��|( P7� PD0�  ����Z3� T0 k� �#��'�"�2't �8t B  ��)    �   W ���B�H EO)��|( P7� PD0�  ����Z3� T0 k� �'��+�"�2't �8t B  ��)    �   W ���B�H EO)���|( P3� TD0� 0����Z3� T0 k� �/��3�"�2't �8t B  ��)    �   W ���B�S�E? )���|( P3��TD0� 0����Z3� T0 k� �;��?�"�2't �8t B  ��)    �   W ���B�[�E>�)���|( �3��TD@�	 0����Z3� T0 k� �G��K�"�2't �8t B  ��)    �   W ���B�_�E>�(���|( �3��XD@�	 0����Z3� T0 k� �O��S�"�2't �8t B  ��)    �   W ���Pc�E>�(���|( �3��XD@�
 0����Z3� T0 k� �S��W�"�2't �8t B  ��)    �   W ��Pg�E>�(���|( �3��\D@� 0����Z3� T0 k� �W��[�"�2't �8t B  ��)    �   W ��Po�E>�'���|( �3��\D@� 0��� Z3� T0 k� �_��c�"�2't �8t B  ��)    �   W  ��Ps�E>�'���|( �/��\E`� 0��� Z3� T0 k� �c��g�"�2't �8t B  ��)    �   W ���Pw�E>�&���|( �/��`E`� 1  �Z3� T0 k� �k��o�"�2't �8t B  ��)    �   W ���P�E.�%���|( �/��dE`� 1�Z3� T0 k� �s��w�"�2't �8t B  ��    �   W ��P ��E.�%���|( �/��hE`� A�Z3� T0 k� �x �| "�2't �8t B  ��    �   W ��P ��E.�$���|(  /��hEP� A�Z3� T0 k� �| �� "�2't �8t B  ��    �   W ��P ��E.�$���|(  /��hEP� A �Z3� T0 k� ���"�2't �8t B  ��    �   W #��P ��E.�#���|(  /��lEP� A$�Z3� T0 k� ���"�2't �8t B  ��    �   W #��P ��B��"���|(  /��lEP� A,1Z3� T0 k� ���"�2't �8t B  ��    �   W #�#�P ��B��!���|(  /��pEP� A41Z3� T0 k� ���"�2't �8t B  ��    �   W '�'�P ��B��!���|(  /��tC� A<1Z3� T0 k� ���"�2't �8t B  ��    �   W '�+�P ��B�� ���|(  /��tC� A@1Z3� T0 k� ���"�2't �8t B  ��    �   W +�/�P ��B�����|(  3��tC� AH1 Z3� T0 k� ���"�2't �8t B  ��    �   W /�;�P��B�����|(  3��xC� AX1"Z3� T0 k� ���"�2't �8t B  ��    �   W /��?�P��B�����|(  7��|C� Q`1"Z3� T0 k� ����"�2't �8t B  ��    �   X 3��C�P��B�����|(  7��|C� Qh	!#Z3� T0 k� ����"�2't �8t B  ��    �   Y�7��K�P��B�����|( �7��|C� Qp
!$Z3� T0 k� ����"�2't �8t B  ��    �   Z�7��O�P��B�����|( �;���C� Qx
!%Z3� T0 k� ��	��	"�2't �8t B  ��    �   [�;��S�P��C�ދ�|( �;� �C� Q�! &Z3� T0 k� ��	��	"�2't �8t B  ��    �   \�?��[�P��C�އ�|( �?� �C� Q�! 'Z3� T0 k� ��
��
"�2't �8t B  ��    �   ]�C��_�P��C�އ�|( �C� � C� Q�!$(Z3� T0 k� ��
��
"�2't �8t B  ��)    �   ^�G�g�P��C�ރ�|( �C� �!C� Q�!$)Z3� T0 k� ��� "�2't �8t B  ��)    �   _�K�k�B���C���|( �G� �"EP� Q�!(*Z3� T0 k� ��"�2't �8t B  ��)    �   `�O�s�B���E.��|( �K��#EP� Q�,+Z3� T0 k� ��"�2't �8t B  ��)    �   a�W��B���E.�{�|( �S��%EP� Q�0-Z3� T0 k� �� "�2't �8t B  ��)    �   b�W���B���E.�w�|( �W��&EP� !�0.Z3� T0 k� �$�("�2't �8t B  ��)    �   c�[���B���E.�w�|( �[��'E@� !�4/Z3� T0 k� �,�0"�2't �8t B  ��)    �   d�_���B���E��s�|( �_��(E@� !��80Z3� T0 k� �4�8"�2't �8t B  ��)    �   e�c���B���E��s�|( �c��)E@� !��<1Z3� T0 k� �<�@"�2't �8t B  ��)    �   f�g���P��E��s�|( �g��*E@� !��@2Z3� T0 k� �D�H"�2't �8t B  ��)    �   g�k����P��E�
�s�|( �k���+E@� !��D3Z3� T0 k� �L�P"�2't �8t B  ��)    �   h�s����P�E��o�|( �s���-E0� !��H4Z3�T0 k� �\�`"�2't �8t B  ��)    �   i�w����P�E��o�|( �{���.E0� "�P5Z3�T0 k� �d�h"�2't �8t B  ��)    �   j�{����P�E��o�|( ����/E0� "�T6Z3�T0 k� �l�p"�2't �8t B  ��)    �   k�����P!�E��s�|( ���	�0E0� "�X7Z3�T0 k� �t�x"�2't �8t B  ��)    �   l������P!�E��s�|( ���	�0E0� " �\8Z3�T0 k� �|��"�2't �8t B  ��)    �   n������P!�E��s�|( ���	�1E � 2(�`9Z3�T0 k� ���"�2't �8t B  ��)    �   p������P!�E��s�|( �	�2E � 20�d9Z3�T0 k� ���"�2't �8t B  ��)    �   r�����P!'�E����w�|( �	 �3E � 2@�p;Z3�T0 k� ���"�2't �8t B  ��)    �   t����P!+�E���w�|( ���	 �3E � 2H�t<Z3�T0 k� ���"�2't �8t B  ��)    �   v����P!/�E���w�|( ���	 �4B� 2P�x<Z3�T0 k� ���"�2't �8t B  ��)    �   x����P!3�E���{�|( ���	 �4B� 2\�|=Z3�T0 k� ����"�2't �8t B  ��)    �   z���#�P7�E���{�|( ���	 �5B� 2d��>Z3�T0 k� ����"�2't �8t B  ��)    �   |���+�P;�E����|( ���	�5B� 2l��?Z3�T0 k� ����"�2't �8t B  ��)    �   ~���3�P?�E����|( �Ä	�5B�
 2t��?Z3�T0 k� ����"�2't �8t B  ��)    �   � ���;�PC�E����|( �Ǆ	�6B�	 2|��@Z3�T0 k� ����"�2't �8t B  ��)    �   � ���G�PG�E�#����|( �τ	�6B� B���AZ3�T0 k� ����"�2't �8t B  ��)    �   � ���O�@K�E�'����|( �ӄ	�6B� B���AZ3�T0 k� ����"�2't �8t B  ��)    �   � ���W�@O�E+����|( �ۄ	 �6B� B���BZ3�T0 k� ����"�2't �8t B  ��)    �   � ���_�@O�E/����|( ��	 �6B� B���CZ3�T0 k� � �"�2't �8t B  ��)    �   � ���g�@S�E3�N��|( ��	 �6B� B���CZ3�T0 k� ��"�2't �8t B  ��)    �   � ���w�@[�E?�N��|( ��	! 7B� B���EZ3�T0 k� �� "�2't �8t B  ��)    �   � ����@_�EC�N��|( ���	 7E � B���EZ3�T0 k� �$�("�2't �8t B  ��)    �   � ����@c�EG�N��|( ���	 7E �  B���FZ3�T0 k� �,�0"�2't �8t B  ��)    �   � ����@g�EK�.��|( ��	7E �� B���GZ3�T0 k� �4�8"�2't �8t B  ��)    �   ����@g�EO�.��|( ��	7E �� B���GZ3�T0 k� �<�@"�2't �8t B  ��)    �   �����@k�ES�.��|( ��	7E �� R���HZ3�T0 k� �D�H"�2't �8t B  ��)    �   �����@o�D�W�.��|( ��	!7E �� R���HZ3�T0 k� �P�T"�2't �8t B  ��)    �   �����@s�D�[�.��|( ��	!7E �� R���IZc�T0 k� �X�\"�2't �8t B  ��)    �   �����@w�D�_���|( �#�	!7E �� R���JZc�T0 k� �`�d"�2't �8t B  ��)    �   �'��ý@w�D�c���|( �'�	!7E �� S� JZc�	T0 k� �h�l"�2't �8t B  ��)    �   �/��˽@{�D�g���|( �+�	!7E�� S�KZc�	T0 k� �p�t"�2't �8t B  ��)    �   �3��Ӽ@�D�k���|( �/� 7E�� S�KZc�
T0 k� �x�|"�2't �8t B  ��)    �   �C���@��D�s����|( �7� 7E�� S$� LZc�
T0 k� ���"�2't �8t B  ��) 	   �   �K���@��D�w����|( �;� 7E�� S0�(MZc�T0 k� ���"�2't �8t B  ��) 	   �   �S����@��D�{����|( �?� 7B��� S8�0MZc�T0 k� ���"�2't �8t B  ��) 	   �   �[����@��D�����|( �C��7B��� S@�4NZc�T0 k� ���"�2't �8t B �) 	   �   �c���@��D�����|( �G��7B���CH�<NZc�T0 k� ���"�2't �8t B ��/ 	   �   �k���@��D������|( �K��7B���CP�DOZc�T0 k� �t�x"�2't �8t B ��/ 	   �   �s���@��D������|( �K��7B���CX�LOZc�T0 k� �d�h"�2't �8t B ��/ 	   �   �{��#�@��D������|( �O��7B���C`�TPZc�T0 k� �X�\"�2't �8t B ��/ 	   �   ��{��+�@��D�� ���|( �S��7B���Ch�\PZc�T0 k� �L �P "�2't �8t B	 ��/ 	   �   �����3�@��D�����|( �S��7B���Cp�dQZc�T0 k� �@!�D!"�2't �8t B ��/ 	   �   �����C�@��F����|( �W��7B���3� �tRZc�T0 k� �("�,""�2't �8t B ��/ 	   �   �����K�@��F����|( �[��7B���3� |RZc�T0 k� �#�#"�2't �8t B ��/ 
   �   }����W�@��F����|( �[��7B���3� �SZc�T0 k� �#�#"�2't �8t B ��/ 
   �   x����_�@��F����|( �[�� 7B���3� �SZc�T0 k� � $�$"�2't �8t B ��/ 
   �   t����g�@��F����|( �_��$7B��3�!�SZc�T0 k� ��%��%"�2't �8t B ��/ 
   �   p����o�@��F����|( �_��(7E�#�!�TZc�T0 k� ��%��%"�2't �8t B ��/ 
   �   l����w�@��E��	���|( �_��,7E�#�!�TZc�T0 k� ��&��&"�2't �8t B ��/ 
   �   h�����@��E��
��|( �_��07E�#�!�UZc�T0 k� �'��'"�2't �8t B ��/ 
   �   d������@��E����|( �_��47E�#�!�UZ3�T0 k� �'��'"�2't �8t B ��/ 
   �   `������@��E����|( �_��<7E'�#�"�UZ3�T0 k� �(��("�2't �8t B ��/    �   \������@��E����|( �_��D7E�3�#�"��VZ3�T0 k� �*��*"�2't �8t B �/    �   \���B��@��E���'�|( �_��H7E�;�#�"��WZ3�T0 k� �*��*"�2't �8t B �/    �   \���B��@��E���+�|( A[��P7E�C�#�"��WZ3�T0 k� �+��+"�2't �8t B ��/    �   \���B��@��E���3�|( A[��T7E�K�#�"��WZ3�T0 k� t,�x,"�2't �8t B  ��/    �   \���Bë@��@��7�|( A[��X7E�S�#�#��WZ3�T0 k� h,�l,"�2't �8t B" ��/    �   \ a��B˪@��@� ?�|( A[��`7E�[�#�#��XZ3�T0 k� \-�`-"�2't �8t B# ��/    �   \ b�BӪ@��@� C�|( AW��d8E�_�#�#��XZ3�T0 k� �P.�T."�2't �8t B$ ��/    �   \ b�B۩@��@� K�|( AW��l8E�g�#�#� XZ3�T0 k� �D.�H."�2't �8t B% ��/    �   \ b�B�@��@� O�|( AS��p8E�o�#�$�XZ3�T0 k� �4/�8/"�2't �8t B& ��/    �   \ b�B�@��@� W�|( AS��x9E�w�$ $�XZ3�T0 k� �(0�,0"�2't �8t B' ��/    �   \ b�B�@��@  [�|( AO��|9E��$%�XZ3�T0 k� �1� 1"�2't �8t B( ��/    �   \ b'�B��@� @ _�|( AO���:Eq��$%sXZ3�T0 k� �1�1"�2't �8t B) ��/    �   \ b+�B��@� @ g�|( 1K���:Eq��$&s$XZ3�T0 k� �2�2"�2't �8t B* ��/    �   \ b3�C�@� @ k�|( 1K���;Eq��$&s,XZ3�T0 k� ��3��3"�2't �8t B* ��/    �   \ b7�C�@�@ o�|( 1G���<Eq�� &s4XZ3�T0 k� ��3��3"�2't �8t B+ ��/    �   \ b?�C�@�@ s�|( 1G���=Eq�� 's<WZ3�T0 k� ��4��4"�2't �8t B, ��/    �   \ bC�C�@�@ {�|( 1C���=Eq��  'sDWZ3�T0 k� ��5��5"�2't �8t B- ��/    �   \ bK�C�@�@ �|( 1C���>Eq�� $'sHWZ3�T0 k� ��5��5"�2't �8t B. ��/    �   \ bO�C'�@�@  ��|( 1?���?Eq�� ,(sPVZ3�T0 k� ��6��6"�2't �8t B. ��/    �   \ bW�C+�@�@$ ��|( 1?���@Eq�� 0(sXVZ3�T0 k� ��7��7"�2't �8t B/ ��/    �   \ b[�C3�@�@( ��|( 1;���AEq�� 4)s\UZ3�T0 k� ��7��7"�2't �8t B0 ��/    �   \ bc�C7�@�@,  ��|( A;���BD��� 8)cdUZ3�T0 k� �8��8"�2't �8t B0 ��/    �   \ bg�C?�@�@0! ��|( A7���CD��� <)clTZ3�T0 k� �9��9"�2't �8t B1 ��/    �   \ bk�CC�@�@4" ��|( A7���DD��� @*cpTZ3�T0 k� x:�|:"�2't �8t B2 ��/    �   \ bs�CK�@�@8" ��|( A3���ED��� D*cxSZ3�T0 k� l:�p:"�2't �8t B2 ��/    �   \ bw�CO�@�@<# ��|( A3���GD��� H*c|SZ3�T0 k� `;�d;"�2't �8t B3 ��/    �   \ b{�CW�@�@@$ ��|( A3���HD��� L+c�RZ3�T0 k� P<�T<"�2't �8t B3 ��/    �   \ b��C[�@�@D$ ��|( A/���ID��� P+c�RZ3�T0 k� D<�H<"�2't �8t B4 ��/    �   \ b��Cc�@ @H% ��|( A/���JD��� T+c�QZ3�T0 k� 8=�<="�2't �8t B4 ��/    �   \ b��Cg�@ @H& ��|( A+���LLQ�� T+c�PZ3�T0 k� ,>�0>"�2't �8t B5 ��/    �   \ b��Ck�@ @L& ��|( A+���MLR� P,c�PZ3�T0 k�  >�$>"�2't �8t B5 ��/    �   \ b��Cs�@@P' ��|( A'���NLR� P,c�OZ3�T0 k� �?�?"�2't �8t B6 ��/    �   \ b��Cw�@@T' ��|( A'���PLR� P,S�NZ3�T0 k� �@�@"�2't �8t B6 ��/    �   \ b��C{�@@X( ��|( Q'���QLR� P-S�MZ3�T0 k� ��@��@"�2't �8t B6 ��/    �   \ b��C�@@\) ��|( Q#���RLR� P-S�MZ3�T0 k� ��A��A"�2't �8t B7 ��/    �   \ b��C��@@\) ��|( Q#���TLR� L-S�LZ3�T0 k� ��B��B"�2't �8t B7 ��/    �   \ b��C��@@`* ��|( Q#���ULR'� L.S�KZ3�T0 k� ��C��C"�2't �8t B7 ��/    �   \ b��C��@@d* ��|( Q���VLR+� L.S�KZ3�T0 k� ��C��C"�2't �8t B8 ��/    �   \ b��C��@@h+ ��|( Q���WLR/� L.S�JZ3�T0 k� иD��D"�2't �8t B8 ��/    �   \ b��C��@@h+ ��|( Q���YLR3� H.S�IZ3�T0 k� ЬE��E"�2't �8t B8 ��/    �   \ b��C��@@l, ��|( Q���ZLR;� H/S�IZ3�T0 k� РE��E"�2't �8t B8 ��/    �   \ b��C��@@p- ��!�( Q���[LR?� H/�Hb��T0 k� ��F��F"�2't �8t B8 ��/    �   \ b��C��@	@p- ��!�( Q���\LRC� H/�Gb��T0 k� ��G��G"�2't �8t B8 ��/    �   \ b��C��@	@t. ��!�( Q���]LbG� H/�Gb��T0 k� �|G��G"�2't �8t B8 ��/    �   \ b��C��@	@x. ��!�( a���^LbK� H0�Fb��T0 k� �lH�pH"�2't �8t B9 ��/    �   \ b��C��@	@x/ ��!�( a���`LbO� D0�Fb��T0 k� �`I�dI"�2't �8t B9 ��/    �   \ b��C��@
@|/ ��!�( a���aLbS� D0�Eb��T0 k� �TI�XI"�2't �8t B9 ��/    �   \ b��C��@
@�0 ��!�( a���bLb[� D0�Db��T0 k� �HJ�LJ"�2't �8t B9 ��/    �   \ b��C��@
@�0 ��!�( a��cLb_� D1�Db��T0 k� �<K�@K"�2't �8t B8 ��/    �   \ b��CÖ@
@�1 ��!�( a��dLbc� D1�Cb��T0 k� �0L�4L"�2't �8t B8 ��/    �   \ b��Cǖ@ 
@�1 ��!�( a��eLbg� @1�Cb��T0 k� � L�$L"�2't �8t B8 ��/    �   \ b��C˕@ @�1 ��!�( a��fLbk� @1�Bb��T0 k�  M�M"�2't �8t B8 ��/    �   \ b��Cϕ@ @�2 �|( a
��gLbo� @1�BZ3�T0 k�  N�N"�2't �8t B8 ��/    �   \ b��Cӕ@$@�2 �|( a��hLbs� @2�AZ3�T0 k� �N� N"�2't �8t B8 ��/    �   \ b��Cה@$@�3 �|( a��iLbw� @2�AZ3�T0 k� �O��O"�2't �8t B8 ��/    �   \ b��Cה@$@�3 �|( q��jLb{� @2�@Z3�T0 k� �P��P"�2't �8t B7 ��/    �   \ b��C۔@$@�4 �|( q��kLb� <2�@Z3�T0 k� ��P��P"�2't �8t B7 ��/    �   \ b��Cߔ@(@�4 �|( q��kLb�� <2�?Z3�T0 k� ��Q��Q"�2't �8t B7 ��/   �   \ b��C�@(@�4 �|( q��lLb�� <3�?Z3�T0 k� �R��R"�2't �8t B7 ��/    �   \ b��C�@(@�5 �|( q��mLb�� <3�>Z3�T0 k� �R��R"�2't �8t B6 ��/    �   \ c�C�@,@�5 �|( 1 ��nLb�� <3�>Z3�T0 k� �S��S"�2't �8t B6 ��/    �   \ c C�@,@�6 �|( 1 ��nLb�� <3�=Z3�T0 k� ϘT��T"�2't �8t B5 ��/    �   \ c C�@,@�6 �|( 1  ��oLb�� <3�=Z3�T0 k� ψU��U"�2't �8t B5 ��/    �   \ c C�@,@�6 �!�( 1 "�oLb�� <4�=bs�T0 k� �|U��U"�2't �8t B5 ��/    �   \ c C��@0@�7 #�!�( 0�%�pLb�� 84�<bs�T0 k� �pV�tV"�2't �8t B4 ��/    �   \ c C��@0@�7 #�!�( 0�'�pLb�� 84�<bs�T0 k� �dW�hW"�2't �8t B4 ��/    �   \ cC��@0@�8 '�!�( 0�)�pLb�� 84�;bs�T0 k� �XW�\W"�2't �8t B3 ��/    �   \ cC��@0@�8 '�!�( 0�+�qLb�� 84�;bs�T0 k� �LX�PX"�2't �8t B3 ��/    �   \ cD�@4@�8 +�!�( 0�-�qLb�� 85�:bs�T0 k� �<Y�@Y"�2't �8t B2 ��/    �   \ cD�@4@�9 /�!�(  �0�qLb�� 85�:bs�T0 k� �0Y�4Y"�2't �8t B1 ��/    �   \ cD�@4@�9 /�!�(  �2�qLb�� 85�:bs�T0 k� �$Z�(Z"�2't �8t B1 ��/    �   \ c D�@4@�9 3�!�(  �4�qLb�� 45�9bs�T0 k� �[�["�2't �8t B0 ��/    �   \ c$D�@8@�: 3�!�(  �6�qLb�� 45�9bs�T0 k� �[�["�2't �8t B/ ��/    �   \ c$D�@8@�: 7�!�(  �8��qLb�� 45�8bs�T0 k� � \�\"�2't �8t B/ ��/    �   \ c(D�@8@�: 7�|(  �;��qLb�� 45�8Z3�T0 k� ��]��]"�2't �8t B. ��/    �   \ c(D�@8@�: ;�|(  �=��pLb�� 46�8Z3�T0 k� ��^��^"�2't �8t B- ��/    �   \ c,D�@8@�: ;�|(  �?��pLb�� 46|7Z3�T0 k� ��^��^"�2't �8t B, ��/    �   \ c0D�@<@�: ?�|(  �A��pLb�� 46x7Z3�T0 k� ��_��_"�2't �8t B, ��/    �   \ c0D�@<@�: ?�|(  �D�|oLb�� 46t7Z3�T0 k� ��`��`"�2't �8t B+ ��/   �   \ c4D�@<@�; C�|(  �F�xoLb�� 46t6Z3�T0 k� ��`��`"�2't �8t B* ��/    �   \ c4D�@<@�; C�|( ! H�tnLb�� 46p6Z3�T0 k� ��a��a"�2't �8t B) ��/    �   \ c8D�@<@�; C�|( ! J�pnLb�� 07l6Z3�T0 k� �b��b"�2't �8t B( ��/    �   \ c8D�@@@�< G�|( L�lmLb�� 07h5Z3�T0 k� �b��b"�2't �8t B' ��/    �   \ c<D�@@@�< G�|( N�hlLb�� 07d5Z3�T0 k� �c��c"�2't �8t B& ��/    �   \ c<D�@@@�< K�|( P�hlLR�� 07d5Z3�T0 k� �td�xd"�2't �8t B% ��/    �   \ c@D�@@@�< K�|( R�dkLR�� 07`4Z3�T0 k� �he�le"�2't �8t B$ ��/    �   \ c@D�@@@�= O�|( T�`jLR�� 07\4Z3�T0 k� �Xe�\e"�2't �8t B# ��/    �   \ cDD�@D@�= O�|( V�\iLR�� 07#X4Z3�T0 k� �Lf�Pf"�2't �8t B" ��/    �   \ cDD�@D@�= O�|( X�XhLR�� 07#X4Z3�T0 k� �@g�Dg"�2't �8t B! ��/    �   \ cHD�@D@�> S�|( Z�TgLR�� 08#T3Z3�T0 k� �4g�8g"�2't �8t B  ��/    �   \ cHD�@D@�> S�|( \�PfD��� 08#P3Z3�T0 k� �(h�,h"�2't �8t B ��/    �   \ cLD�@D@�> W�|( �\�TeD��� 08#L3Z3�T0 k� i� i"�2't �8t B ��/    �   \ cLD�@D@�> W�|( �]�TeD��� ,8#L2Z3�T0 k� i�i"�2't �8t B ��/    �   \ cPD�@H@�? W�|( �^QTeD��� ,8#H2Z3�T0 k�  j�j"�2't �8t B ��/    �   \ cPD#�@H@�? [�|( �_QXdD��� ,8#D2Z3�T0 k� �k��k"�2't �8t B ��/    �   \ cTD#�@H@�? [�|( �_QXdD��� ,8#D2Z3�T0 k� �k��k"�2't �8t B ��/    �   \ cTD#�@H@�? _�|( �`QXdD��� ,8#@1Z3�T0 k� ��l��l"�2't �8t B ��/    �   \ cXD#�@H@�? _�|( �aQ\cEr���,9#<1Z3�T0 k� ��m��m"�2't �8t B ��/    �   \ cXD#�@H@�@ _�|( �bQ\cEr���,9#<1Z3�T0 k� ��n��n"�2't �8t B ��/    �   \ cXD'�@H@�@ c�|( �cQ\cEr���,9#81Z3�T0 k� ݴn��n"�2't �8t B ��/    �   \ c\D'�@L@�@ c�|( �cQ\bEr���,9#80Z3�T0 k� ݨo��o"�2't �8t B ��/    �   \ c\D'�@L@�@ c�|( �dQ`bEr���,9#40Z3�T0 k� ��p��p"�2't �8t B ��/    �   \ c`D'�@L@�A g�|( �eQ`bEr���,9#00Z3�T0 k� ��p��p"�2't �8t B ��/    �   \ c`D'�@L@�A g�|( �fa`aEr� �,9#00Z3�T0 k� ��q��q"�2't �8t B ��/    �   \ c`D'�@L@�A g�|( � fadaEb��,9#,/Z3�T0 k� �xr�|r"�2't �8t B ��/    �   \ cdD+�@L@�A k�|( � gadaEb��(9#,/Z3�T0 k� �hr�lr"�2't �8t B
 ��/    �   \ cdD+�@L@�A k�|( ��had`Eb��(9#(/Z3�T0 k� �\s�`s"�2't �8t B ��/    �   \ cdD+�@P@�B k�|( ��had`Eb��(:#(/Z3�T0 k� �Pt�Tt"�2't �8t B ��/    �   \ chD+�@P@�B k�|( ��iah`Ec �(:#$/Z3�T0 k� �Dt�Ht"�2't �8t B ��/    �   \ chD+�@P@�B o�|( ��jah`D3 �(:# .Z3�T0 k� �8u�<u"�2't �8t B ��/    �   \ clD+�@P@�B o�|( ��jah_D3 �(:# .Z3�T0 k� �,v�0v"�2't �8t B ��/    �   \ clD/�@P@�B o�|( ��kah_D3 	�(:#.Z3�T0 k� �w� w"�2't �8t B  ��/    �   \ clD/�@P@�B s�|( ��lQh_D3 
�(:#.Z3�T0 k� �w�w"�2't �8t B  ,�/    �   \ cpD/�@P@�C s�|( ��lQl_D3 �(:#.Z3�T0 k� �x�x"�2't �8t B  ��/    �   \ cpD/�@P@�C s�|( ��mQl^D3 �(:#-Z3�T0 k� ��y��y"�2't �8t B ��/    �   \ cpD/�@T@�C s�|( ��mQl^D3 �(:#-Z3�T0 k� ��y��y"�2't �8t B ��/    �   \ ctD/�@T@�C w�|( ��nQl^D3 �(:#-Z3�T0 k� �z��z"�2't �8t B ��/    �   \ ctD/�@T@�C w�|( ��oQp^D3 �(:#-Z3�T0 k� �{��{"�2't �8t B ��/    �   \ ctD3�@T@�C w�|( ��oQp]D2��(;#-Z3�T0 k� �{��{"�2't �8t B ��/    �   \ ctD3�@T@�D w�|( ��pQp]DB��(;#,Z3�T0 k� �|��|"�2't �8t B ��/    �   \ cxD3�@T@�D {�|( ��pQp]DB��(;#,Z3�T0 k� �}��}"�2't �8t B ��/    �   \ cxD3�@T@�D {�|( ��q�p]DB��(;#,Z3�T0 k� �}��}"�2't �8t B ��/    �   \ cxD3�@T@�D {�|( ��q�t]DB��(;#,Z3�T0 k� �~��~"�2't �8t B ��/    �   \ c|D3�@T@�D {�|( ��r�t]DB��$;#,Z3�T0 k� ���"�2't �8t B ��/    �   \ c|D3�@X@�D �|( ��r�t]DB��$;#,Z3�T0 k� x��|�"�2't �8t B ��/    �   \ c|D3�@X@�E �|( ��s�t]DB��$;#,Z3�T0 k� l��p�"�2't �8t B ��/    �   \ c|D7�@X@�E �|( ��s1t]DB��$;#-Z3�T0 k� �`��d�"�2't �8t B	 ��/    �   \ c�D7�@X@�E �|( ��t1t]DB��$;#-Z3�T0 k� �T��X�"�2't �8t B	 ��/    �   \ c�	D7�@X@�E ��|( ��t1t]DB��$;.Z3�T0 k� �H��L�"�2't �8t B
 ��/    �   \ c�	D7�@X@�E ��|( ��u1t]DB��$; .Z3�T0 k� �<��@�"�2't �8t B
 *�/    �   \ c�	D7�@X@�E ��|( ��u1t]DR��$; .Z3�T0 k� �0��4�"�2't �8t B
 ��/    �   \ c�	D7�@X@�E ��|( ��v1t]DR��$; /Z3�T0 k� �$��(�"�2't �8t B
 ��/    �   \ c�	D7�@X@�F ��|( ��v1t]DR� �$< /Z3�T0 k� ����"�2't �8t B	 ��/    �   \ c�	D7�@X@�F ��|( ��w1t]DR�!�$< 0Z3�T0 k� ��"�2't �8t B	 ��/    �   \ c�	D;�@\@�F ��|( ��w1t]DR�"�$<��0Z3�T0 k� �~�~"�2't �8t B	 ��/    �   \ c�	D;�@\@�F ��|( ��x1t]DR�#�$<��1Z3�T0 k� ��}��}"�2't �8t B ��/    �   \ c�	D;�@\@�F ��|( ��xt]DR�#�$<��1Z3�T0 k� ;�|��|"�2't �8t B ��/   �   \ c�	D;�@\@�F ��|( ��xt]DR�$�$<��2Z3�T0 k� ;�{��{"�2't �8t B ��/    �   \ c�	D;�@\@�F ��|( ��yt]DR�&�$<��2Z3�T0 k� ;�y��y"�2't �8t B ��/    �   \ c�	D;�@\@�F ��|( ��yt]DR�'�$<��2Z3�T0 k� ;�x��x"�2't �8t B ��/    �   \ c�	D;�@\@�G ��|( ��zt]DR�(�$<��3Z3�T0 k� ;�v��v"�2't �8t B ��/    �   \ c�	D;�@\@�G ��|( ��zt]Db�)�$<��3Z3�T0 k� ��t��t"�2't �8t B ��/    �   \ c�
D;�@\@�G ��|( ��zt]Db�*�$<��4Z3�T0 k� ��r��r"�2't �8t B ��/    �   \ c�
D;�@\@�G ��|( ��{t]Db�+�$<��4Z3�T0 k� ��q��q"�2't �8t B ��/    �   \ c�
D?�@\@�G ��|( ��{t]Db�,�$<��4Z3�T0 k� ��o��o"�2't �8t B ��/    �   \ c�
D?�@\@�G ��|( ��|t]Db�-�$<��5Z3�T0 k� ��m��m"�2't �8t B ��/    �   \ c�
D?�@`@�G ��|( ��|t]Db�0�$<��5Z3�T0 k� +�i��i"�2't �8t B ��/    �   \ c�
D?�@`@�G ��|( ��}
�t]Db�1�$=��6Z3�T0 k� +�h��h"�2't �8t B ��/    �   \ c�
D?�@`@�H ��|( ��}
�t]Db�2� =��6Z3�T0 k� +�f��f"�2't �8t B ��/    �   \ c�
D?�@`@�H ��|( ��}
�t]Db�4� =��7Z3�T0 k� +�d��d"�2't �8t B  ��/    �   \ c�
D?�@`@�H ��|( ��~
�t]Db�5� =��7Z3�T0 k� +�b��b"�2't �8t B  ,�/    �   \ c�
D?�@`@�H ��|( �~
�t]D2|7� =��7Z3�T0 k� ��`��`"�2't �8t B  ��/    �   \ c�
D?�@`@�H ��|( �~
�t]D2t8� =��8Z3�T0 k� �|^��^"�2't �8t B  ��/    �   \ c�
D?�@`@�H ��|( �
�t]D2p9� =��8Z3�T0 k� �x\�|\"�2't �8t B  ��/   �   \ c�
DC�@`@�H ��|( �
�t]D2h;� =��8Z3�T0 k� �xZ�|Z"�2't �8t B  ��/    �   \ c�
DC�@`@�H ��|( �
�t]D2d<� =�8Z3�T0 k� �tX�xX"�2't �8t B  ��/    �   \ c�
DC�@`@�H ��|( ��
�t]Eb\>� =�9Z3�T0 k� �pV�tV"�2't �8t B  ��/    �   \ c�
DC�@`@�H ��|( ��
�t]EbX?  =�9Z3�T0 k� �pT�tT"�2't �8t B  ��/    �   \ c�
DC�@`@�H ��|( ��
�t]EbPA  =�9Z3�T0 k� �lR�pR"�2't �8t B  ��/    �   \ c�
DC�@`@�I ��|( ��
�t]EbLB  =�:Z3�T0 k� �lP�pP"�2't �8t B  ��/    �   \ c�
DC�@d@�I ��|( ��
�t]EbDC  =�:Z3�T0 k� �hN�lN"�2't �8t B  ��/    �   \ c�
DC�@d@�I ��|( ��
�t]Eb@E  =�:Z3�T0 k� �hL�lL"�2't �8t B  ��/    �   \ c�DC�@d@�I ��|( ��
�t]Eb8F  =�;Z3�T0 k� �hJ�lJ"�2't �8t B  ��/    �   \ c�DC�@d@�I ��|( ��
�t]Eb4H  =�;Z3�T0 k� �hH�lH"�2't �8t B  ��/    �   \ c�DC�@d@�I ��|( ��~
�t]Eb,I  =�;Z3�T0 k� �dF�hF"�2't �8t B  ��/    �   \ c�DC�@d@�I ��|( ��~
�t]ER(K  =�;Z3�T0 k� �dD�hD"�2't �8t B  ��/    �   \ c�DC�@d@�I ��|( ��~
�t]ER L  =�<Z3�T0 k� �dC�hC"�2't �8t B  ��/    �   \ c�DG�@d@�I ��|( ��}
�t]ERM  =�<Z3�T0 k� �dA�hA"�2't �8t B  ��/    �   \ c�DG�@d@�I ��|( ��}
�t]ERO  >x<Z3�T0 k� �d?�h?"�2't �8t B  ��/    �   \ c�DG�@d@�I ��|( ��}
�t]ERP  >t<Z3�T0 k� �d=�h="�2't �8t B  ��/    �   \ c�DG�@d@�I ��|( ��|
�t]C�Q  >l=Z3�T0 k� �d;�h;"�2't �8t B  ��/    �   \ c�DG�@d@�J ��|( ��|
�t]C� S  >h=Z3�T0 k� �d:�h:"�2't �8t B  ��/    �   \ c�DG�@d@�J ��|( ��{
�t]C��T  >R`=Z3�T0 k� �d8�h8"�2't �8t B  ��/    �   \ c�DG�@d@�J ��|( ��z
�t]C��U  >RX=Z3�T0 k� �d6�h6"�2't �8t B  ��/    �   \NH3 7�A��BM�/�o��L�ߚ��LL��g�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NH3 7�A��BM�/�o��L�ߚ��LL��g�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NH3 7�A��BM�/�o��L�ߚ��LL��k�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NH3 7�A�� BM�/�o��Lߚ��LL��k�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NH3 7�A�� BM�/�o��Lߚ��LL��k�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NL3 ;�A�� BM�0�o�"�Lߚ� LL��k�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NL3 ;�A���BM�0�o�"�Lߚ�LL��k�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NL3 ;�A���BM�0�o�"�Lߚ�LL��o�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NL3 ;�A���BM�0�o�"�Lߚ�LL��o�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NL3 ;�A���BM�0�o�"�Lߚ> LL��o�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NL3 ;�A���BM�0�o�"�Lߚ> #LL��o�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NL3 ;�A���BM�0�o�"�Lߚ>$%LL��o�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8NL3 ;�A���BM�0�o�"�Lߚ>$%LL��s�l�bs��T0 k� ���#�P "�2't �8t B �_    ����8�P4 ;�A���BM�0�o�"�Lߚ>$&LL�|s�l�bs��T0 k� ���#�P "�2't �8t B ��_    ����8�P5 ;�A���BM�0�o�"�Lߚ>('LL�|s�l�
bs��T0 k� ���#�P "�2't �8t B ��_    ����8�T6 ;�A���BM�0�o�"�Lߚ>,(LL�|s�l�
bs��T0 k� ���#�P "�2't �8t B ��_    ����8�T7 ;�A���BM�0�o��Lߚ>,)LL�|s�l�
bs��T0 k� ���#�P "�2't �8t B ��_    ����8�X8 ;�A���BM�0�o��Lߚ>0*LL�|s�l�	bs��T0 k� ���#�P "�2't �8t B ��_    ����8�\8 ;�A���BM�0�o��Lߚ>0*LL�|w�l�	bs��T0 k� ���#�P "�2't �8t B ��_    ����8�\9 ;�A���BM�0�o��Lߚ>4+LL�Lw�l�	bs��T0 k� ���$P "�2't �8t B ��_    ����8�`: ;�A���BM�0�o��Lߚ>4,L<�Lw�l�bs��T0 k� ���$P "�2't �8t B ��_    ����8�`; ;�A���BM�0�o��Lߚ>8-L<�Lw�l�bs��T0 k� ���$P "�2't �8t B ��_    ����8�d; ;�A���BM�0�o��Lߚ>8.L<�L{�l�bs��T0 k� ���$P "�2't �8t B ��_    ����8�d< ;�A���BM�0�o��Lߚ></L<�L{�l�Z3��T0 k� ���$P "�2't �8t B ��_    ����8�h= ;�A���BM�0�o��Lߚ></L<���l�Z3��T0 k� ���#KP "�2't �8t B ��_    ����8�h> ;�A���BM�0�o��Lߚ>@0L<���l�Z3��T0 k� ���#KP "�2't �8t B ��_    ����8�l> ?�A���BM�0�o��Lߚ>@1A�����l�Z3��T0 k� ���#KP "�2't �8t B ��_    ����8�l? ?�A���BM�0�o�"�Lߚ>D2A�����l�Z3��T0 k� ���#KP "�2't �8t B ��_    ����8�p@ ?�A���BM�0�o�"�Lߚ>D2A�����l�Z3��T0 k� ���#KP "�2't �8t B ��_    ����8�pA ?�A���BM�0�o�"�Lߚ>H3A�����l�Z3��T0 k� ���#[P "�2't �8t B ��_    ����8�tA ?�A���BM�0�o�"�Lߚ>H4A�����\�Z3��T0 k� ���#[P "�2't �8t B ��_    ����8�tB ?�A���BM�0�o�"�Lߚ>L4A�����\�Z3��T0 k� ���#[P "�2't �8t B ��_    ����8�xC ?�A���BM�0�o�"�Lߚ>L5A�����\�Z3��T0 k� ���#[P "�2't �8t B ��_    ����8�xC ?�A���BM�0�o�"�Lߚ>L6A�����\�Z3��T0 k� ���#[P "�2't �8t B ��_    ����8�|D ?�A���BM�0�o�"�Lߚ>P6A�����\�b���T0 k� ���#kP "�2't �8t B ��_    ����8�|D ?�A���BM�0�o�"�Lߚ>P7A�����\�b���T0 k� ���#kP "�2't �8t B ��_    ����8��E ?�A���BM�0�o�"�Lߚ>T8A�����\�b���T0 k� ���#kP "�2't �8t B ��_    ����8��F ?�A���BM�0�o�"�Lߚ>T8A�����\�b���T0 k� ���#kP "�2't �8t B ��_    ����8��F ?�A���BM�0�o��Lߚ>T9A�����\�b���T0 k� ���#kP "�2't �8t B ��_    ����8��G ?�A���BM�0�o��Lߚ �X:A�����\�b���T0 k� ���#{P "�2't �8t B ��_    ����8��G ?�A���BM�0�o��Lߚ �X:A�����\�b���T0 k� ���#{P "�2't �8t B ��_    ����8��H ?�A���BM�0�o��Lߛ �\;A�����\�b���T0 k� ���#{P "�2't �8t B ��_    ����8��I ?�A���BM�0�o��L� �\;A�����\�b���T0 k� ���#{P "�2't �8t B ��_    ����8��I ?�A���BM�0�o��L� �\<A�����\�b���T0 k� ���#{P "�2't �8t B ��_    ����8��J ?�A���BM�0�o��L�� �`<A�����\�b���T0 k� ���#�P "�2't �8t B ��_    ����8��J ?�A���BM�0�o��L�� �`=A��̧�\�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��K ?�A���BM�0�o��L�� �`>A��̧�\�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��K ?�A���BM�0�o��L�� �d>A��̫�\�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��L ?�A���BM�0�o��L�� �d?A��̫�\�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��L ?�A���BM�0�o��L�� �d?A��̫�\�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��M ?�A���BM�0�o��L�� �h@A��̫�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��M ?�A���BM�0�o��L�� �h@A��̫�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��N ?�A���BM�0�o��L�� �hAA��̫�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��N C�A���BM�0�o��L�� �lAA��̫�l�Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��O C�A���BM�0�o��L�� �lBA��̫�l�Z3��T0 k� ���#�P "�2't �8t B ��_   ����8��O C�A���BM�0�o��L�� �lBA��̫�l� Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��P C�A���BM�0�o��L�� �pCA��̫�l� Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��P C�A���BM�0�o��L� �pCA��̯�l� Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��P C�A���BM�0�o��L� �pCA��̯�l� Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��Q C�A���BM�0�o��L� �pDA��̯�l� Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��Q C�A���BM�0�o��L� �tDA��̯�l� Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��R C�A���BM�0�o��L� �tEA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��R C�A���BM�0�o��L� �tEA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��R C�A���BM�0�o��L� �xFA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��S C�A���BM�0�o��L��xFA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��S C�A���BM�0�o��L��xFA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��T C�A���BM�0�o��L��xGA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��T C�A���BM�0�o��L��|GA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��T C�A���BM�0�o��L��|HA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��U C�A���BM�0�o��L��|HA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��U C�A���BM�0�o��L��|HA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��V C�A���BM�0�o��L�ހIA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��V C�A���BM�0�o��L�ހIA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��V C�A���BM�0�o��L�ހJA��̯�l��Z3��T0 k� ���#�P "�2't �8t B ��_    ����8��W C�A���BM�0�o��L��JA��̯�l��Z3��T0 k� ���$P "�2't �8t B ��_    ����8��W C�A���BM�0�o��L��JA��̯�l��Z3��T0 k� ���$P "�2't �8t B ��_    ����8��W C�A���BM�0�o��L��KA��̯�l��Z3��T0 k� ���$P "�2't �8t B ��_    ����8��X C�A���BM�0�o��L��KA��̳�l��Z3��T0 k� ���$P "�2't �8t B ��_    ����8��X C�A���BM�0�o��L��KA��̳�l��Z3��T0 k� ���$P "�2't �8t B ��_    ����8��X C�A���BM�0�o��L��LA��̳�l��Z3��T0 k� ���#;P "�2't �8t B ��_    ����8��X C�A���BM�0�o��L��LA��̳�l��Z3��T0 k� ���#;P "�2't �8t B ��_    ����8��Y C�A���BM�0�o��L��LA��̳�l��Z3��T0 k� ���#;P "�2't �8t B ��_    ����8��Y C�A���BM�0�o��L��MA��̳�l��Z3��T0 k� ���#;P "�2't �8t B ��_    ����8��Y C�A���BM�0�o��L�ވMA��̳�l��Z3��T0 k� ���#;P "�2't �8t B ��_    ����8��Z C�A���BM�0�o��L�ވMA��̳�l��Z3��T0 k� ���#[P "�2't �8t B ��_    ����8��Z C�A���BM�0�o��L�ތMA��̳�l��Z3��T0 k� ���#[P "�2't �8t B ��_    ����8                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��� ]�$�$� � �� [|          � ��     T. 拭     n �                  5          `     ���   @

"         ��m   $ $       �f�    ���eV�    � �            � 5�        �p     ���   8	(          zZ            ��,     p� ���     � �                7          j`     ���    	
'
           J8�         ;:o     J%� ;+�     �               ���           �0     ���   8		          ��.k          . 'o�    ��'� 'R�     a�   
                          ��     ���   X	           �^  ��      B�
>�      �^�
>�           
                   ����               O  ���    0 0	           z�  N N      V ;k�     {� :��    ���             Z \         �`�  	  ��@  0

 
          ]  � �	     j ]�^     ] ]�^                     	 Z \            
`     ��P   8�          U� > >      ~ }�     T�7 �    ���           	 Z \          0�   
  ��`  (
            >=y   b     �la     >3Pp�     ���            U  Z \         	  ��     ��H   (            =�-  U U  	   � ���     =�' �}    ���             / Z \         
 L�b     ��@ P
B          ���
	      � �S�     � �Cn     - �                       ���_              O  ��@    8	 1	                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          6��  ��        ����D     8l����    �                    x        �       j  �   �	   �                          6    ��        ���       8  ��           "                                                �                          � � ; '�
 ; ] } � �������   
        	      
  y   �A ���A       4� `j� 5d k� 5� k� >D `o� ? @p� ?� q  %� `t� &d u� &� u����  ����. ����< ����J ����X ����X � �� p� �d �t� �d u� � �r@ �  s@ 
�\ V� 
�� V� 
�\ W  
�< W� 
�� W� 
�\ W� �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� � }`���� ����� ����� � � �^@ � _@  � �[� � \� ä }@ � �j� � k�  � �m@ � n@ �� �o� �� p� � �r@ �  s@���� � D� \� $� �j� %� k� �� ^@ �� �^` �� _` �$ }@ GD `t� H 0u� Hd u� H� v  JD �r@ KD 0s@ K�  s� 
�� U� 
�\ V  
�| V  
�< V� 
�� V� 
� W  
�� W� 
�\ W� 
�| W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� \   ����  ������  
�fD
��L���"����D" � j  "  B   J jF�"     "�j  " ��
��
��"    B�j l �  B �
� �  �  
�  ��  ��     � �  �        ��     � �       >��  ��     �          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �/'      �� T ���        �> �  ��        �        ��        �        ��        �  	   w�     ��e���        ��                         ���    	 ���                                    �                  ����            	  �	���%��     \��                 27 Jeremy Roenick y    1:33                                                                        7  5     � �
�1C. � �cVq � c\s c]i �KA �cjV � crV � 	csW � 
k�D �c�9 �c�1 �K NB� \B� �"�
 � "� �"� � *� � *� � *� � *� �"� � *� �"� � *� � *� � *� � *� � *� � *� ] � ] 
�  y ""�# i#� i 
�  t 
�  � 
� �'� � 
� � )"� �*� � 
� 
� � 
� � 
� �H /*P�X  *H�H 1*P�X  *H� � 3"�] 4�G 5
�V@  "H �X  *H�H 8*P�X  *H� �:*:s � ;*Gs �  *As � =*Fs �>*:s �  *Gs                                                                                                                                                                                                                         L� R @       �    ` 
             _ P E `  ������   	            �������������������������������������� ���������	�
��������                                                                                          ��    �~� #  ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, 8  < >��� S� � ��@=���@c�@���A���F�r���&��                                                                                                                                                                                                                                                                                                              h�@�                                                                                                                                                                                                                                          	    n    ; !   ��  4�J     �h  	                           ������������������������������������������������������                                                                                                                                     �  �     h       j          ��               	 
     ��������������������� ���������������������������� � ���� ���������������� ����� ������������������ ���� ������������ ���� � ����� ��� ��� �������� ������ ����������� ������� ��������  ��� �� �� ���� �������������� �������� ���           R                     6 !    �  L�J      .$                             ������������������������������������������������������                                                                   	                                                             �    �4             �          �4 R               	 	 ����  ��������� ������� ����������������� ������� ����� �������� ����� �� ��� � �  �� ��� ������������ ������������������ ������������������ ������������������������������� ���������� ���� �������� ����� ����� ��� ������� ���                                                                                                                                                                                                                                                                                                                      �             


             �  }�         ��������       ��������   ����������������  R|������������������������  'p����������������������������               y�                                          +  '�                  ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 2 G :                                 �  ��] �t�       	t�S$
�C$+TA                                                                                                                                                                                                                                                             
)n1n  �        e            k      k      k                  a                                                                                                                                                                                                                                                                                                                                                                                                          @   	>�  J�  2�  2�  Fa�  ��v�X��� �������̞���̞�*�̞�d��������@�        6   x�B :�� |		         �   & AG� �   �              ���                                                                                                                                                                                                                                                                                                                                       N I   �                      !�� !��                                                                                                                                                                                                                        Y��   �� � ���      �� 8      ��������������������� ���������������������������� � ���� ���������������� ����� ������������������ ���� ������������ ���� � ����� ��� ��� �������� ������ ����������� ������� ��������  ��� �� �� ���� �������������� �������� �������  ��������� ������� ����������������� ������� ����� �������� ����� �� ��� � �  �� ��� ������������ ������������������ ������������������ ������������������������������� ���������� ���� �������� ����� ����� ��� ������� ���   ��      $����������������˪�������������������������������������f��ff��ff�������̺�ff�fffffffffffffffffff����ƹ��ffʻfff�fffjffffffffffff��������������������ʺ��l���f˪������������������������������������������������������������������fff�fff�fff�ffk�ffi�ff��ff��ff�ffffffff�fff�x�����w��xx�������wfffffff�ffff�fffww��ww�x����wx��fk��ff��ff��ffʹffj��fʪ�f�ˊ�k������������ʚ��������������������������������������������˫��ʫ��ff��fl��fl��ff̫fff�ffʬ�f���f�����������wu���w��l������f����W��������xww��Wy�l����x������k���W�fi���j���j���f����˘�����y�y�y����������������������������������������������������ʻ����ʫɚ�����l���ƨ�lƘ�j���k���̜i���j���kxx���wx������wx������������ƈx����������������wW����w�������������������������z����������˫��̺������������������������������������������������������������ʺ������k������������������������������������������x�j���˙�x�˘��̩�x������x���xx�x������x������wx���˫��ʫ����������˪�����ʻ��������������������������������������ʻ�ʻ�����ʪ̫����˺��������������������˪�����f���k��f��fǶW�g���k���̻���f������������������x�������˩f̺�����uw�����w��x�wXx��˪�����������l����l���i��ƹx�f�������������������ʫUW��UUU�UUUX      C   &   F   +�  8                       8     �   �����J����      ��     ��   �     � �   �      � �     �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �t� � ���t� � �$ ^$    ���        ��   �   �    >     �f ��        p���� ��   p���� �$     `d ��     `d �$ ^$ �@          �� �      W   � 
�� ��    ����� ��  ����� �$ ^$��    �  �         ��  ^@   * .j  �E t� = �� t� = N�] �  ��U  �      �   d   ���� e����J g���        f ^�         ���              ���h�������J���J��r����      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  "  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��  DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰ wwwywww�www�www�www�www�www�www����������!��������������������a��������݈����������a������������(-�a������!�-���www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�www�������������������������������������!�����!�-����������!-�����������!������www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�www������m����������݈����������������a݈�����m����!�����������a�-������www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�wwwy-��������!�����������������������������������!��������                                          �      �  a r!   f�"""""*��**"*�"�""�""v""*f   "  ""- ��"�"*"-""z"""""����            n   �  "  q  ��                          �  �                                 � gv"!g�vg�vggfvv|�b��r""gb"�vr�rgb��v���g���v���***�*q!q�"!a�!vwfqqr~� qw��q�~~q�����~~~�w~~w�w            �   ~   ��  ~~  �w      v    �                ggj�vvggvvgg!vg�g֪vvg�r�r��⢪rq**gjb�v�q*gjj*vv��gg�z�/�"!�"�*�""*z����qw�~q~ww��q~qwvq�w�`� ��� �w �~p w�p  ��                    �                        lggz�v��g        �       ggbvvrgggavvvqggav� �      ���w!z�w"""�!""*�"! ��        q� q�        `               �        �                      wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            "! "   "      ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """"! "   "      ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       "! "   "      ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                              	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           "� /���  �       �   �   �                                              �  � �              "                           ��  ����� ��                           �   ���                            "  "  "                            ���                          ����                  �   �� �       �  �  "�  "   "                                                 �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   �   " � ��      �    �   �   �"  ""  !� �� ��  �               �   " ��.�  ��                                               �".��".  ���    �                    �   ���                                                                                                                                                                                                       �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �               �   �       �       Ț  ��  ��" �"��"/��"���  �             "   "      �  �                         �  ���               �".��".  ���    �    �   �                            �   �                        �   �   .   .�   �       �         � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                          �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �"  "�  ���        �                              �  ��  ��  ww  &'  vv  w                   �   �                      �".��".  ���    �              .  ". ""  "    � ���                                    ""  "".  . �    �                                                                                                                                        �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �           "   "   �  �                              �          �   � � /  �"" �"  �                       �   �                      �".��".  ���    �                    ".  ".  ���              �  �˰ ��� �wp �&                                                                                                                                                                                    �� �����ݼڜ��ک��ک��z�	��� 
�� 
�� 	�� ̘ ɪ  ��  �  �� �� ������������ ���  � � � �� "� "��"�/ ��                      �   ��  ��  �̰ ��� ��˰�̻��̻���������ˉ�U��EP�ET �I� ٕ  �D� �L� ��� ��" ����/�"�"�""�����                         �"  �". �.  �                                        �� ��                  �          �         �   �  �  �   �     �  .   .     �   �  ��  �                                                                                                                    �  �  "   "                                                                     ˰ ̻ ̻ �� {�  �� 
�� ��� ��� ������
���	��ܻ̍ݻ���"� 8"  8  �  D�  H�  X�  ��  �   �          "  "     �                        ��  ��� �̺�̻����ۻ�˽��̽��̝ ̙� �30 �EP �U@ �T0 EC0 T3  C:  K�  �"  �"/ ����˽� �"� "" �""� � �� ��      �   �  .�  ."  �            �   �"  ""  !� �� ��  �               �   " ��.�  ��           �   �    �   �       �   �   �                .                         � ��                  �  �˰ ��� �wp �&                                                                                                                                                                   ̻  ��  rb  wg 
�w ���
���ɛ������̽�̪��̙���̻̽̽���٘"#3 ""DR�U� T� �� 	��  ��  ,� "� "� ""��""�������� �  ��   �   p   z   ��  ��  ��� �̹ �ؚ �ک ��������������32"�D2" UR" EU@ EU@ 4U@ K˰ 
�� ��  �   "   ""  "" ��"/���� �� �     ��  "�  "�  "�  "�  ��  �                             �� ̽                       "  �"  �                    �   �                      �".��".  ���    � "� "     �  �   �   �         ��   �  ��  �  �  �         � ".��".��/����  �                                �   "                                                                                                    � 
��	�˽���w��rb��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            .  .     �   �           .          �  ��  �".���.  ��                           "  "  "  "                       �  ��  ��  ww  &'  vv  w                �                        ��"� �"� ����                              "  .���"    �     �                                                                                                                                                                                     �w ��� ɪ�����̻����̙���̍�̻�� �� ��� �DD
UUD
C33
UC D� ̀  ��  ��  +�  "  "/���/ ���   �   ��  ��  ��  ˠ  ��  ��  �   �   �0  D0  ED  5T  4T@ D@ �� ��  ��  ��  "" �" �����               �� �� �� �� ��         "   "                            ,  �.�+��+    ��             �       �   �                   �   �       "  "  �"  ̰  ˰  ��  ��  �               �   �                             �"  �""� "�       "   "   "�  �                            �   ���                            �   "                                                                                                                       �  ɪ� ɪ� ̚� �ȍ ͷ  "�  "� .( 3># �4�
�T��T�"�UN"�UN(�Dɜ� ʨ����, � /�������� � ��                                ��  ��  ��  g}  &'� vz� gz� ̊� �ɩ 8̜ D<� T� @��  �� ɀ ��  ��  "   .          �  ��  �".���.  ��                           "  "  "  "                  D   L   �   �   �   ��  .�"." "."   /�  �  �              � ��         �� �� �� g} &' vw                       "  .���"    �     �                                                                                                                                                                                           �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ����))������؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� ����"  �". �.  �                                        �� ��                  �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                   2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                            @  A   �  D   D                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=""""��������AA�A    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ADA�LL��L�D����3333DDDD x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(XxLL����������D����3333DDDD w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""����������A������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(""""�������I�I������ �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�""""�������I��D���I������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`�D�M�D���M������3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(MD�M�A�����MD�����3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(�""""�����AMAD������ � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(�""""������������������ � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(""""wwwwwwwGGwGGwGwGw �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((�UQUUQUUQUUQUUUDUUUUU3333DDDD ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`DEQQUUDUTEUUUU3333DDDD M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M""""������������������������ � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(�""""�������DAADAI � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(��A�AM�M�DM��M334CDDDD 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5DD����M��DM�����3333DDDD x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x""""wwwwwwDGqGq w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwwGwwDGwwwwwwww + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+ADAH�DJ�H�H�����3333DDDD � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(��H��J�AD�DH�D����3333DDDD � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(�""""�������DD����� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
�1C. � �cVr c^j �KA �cjV � crV � csW �	k~L � 
k�D �c�9 �c�1 �K NB� \B� �"�
 � "� �"� � *� � *� � *� � *� �"� � *� �"� � *� � *� � *� � *� � *� � *� ] � ] 
�  y ""�# i#� i 
�  t 
�  � 
� �'� � 
� � )"� �*� � 
� 
� � 
� � 
� �H /*P�X  *H�H 1*P�X  *H� � 3"�] 4�G 5
�V@  "H �X  *H�H 8*P�X  *H� �:*:s � ;*Gs �  *As � =*Fs �>*:s �  *Gs3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������ �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� � � � � � � � � � � � � � � � � � � � ����������������������������������������������������<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ���������������������������������������������������� � � � � � � � � � � � � � � � � � � � ���������������������������������������������������� � � � � � � � � � � � � � � � � � � � �����������������������������������������!��9�G�Z��6�G�0�U�T�Z�G�O�T�K� � � � � � �,�>�0����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0�����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ��"�������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�2�3� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            