GST@�                                                            \     �                                               d  �                         ���2���r�	 J�������ĸ��p�������        i      #    ����                                d8<n    �  ?     |�����  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"     "�j��   * ��
  ?                                                                               ����������������������������������       ��    =b 0Qb 4 114  4c  c  c      	 
      	   
       ��G �� � ( �(                 Ehp )1         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                ��  �       �   @  #   }   �                                                                                '    E)h1p  �    H   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������     ��A��N���0'���Y|?�/f�@RA_ SL.�`^�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA^�SL.�`^�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA^�SL.�`^�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA^�SL.�`^�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@SA^�SL.�`^�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@SA^�SL�`^�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@SA^�SL�`^�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@TA^�SL�`^�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@TA^�SL�a^�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@TA^�SL�a^�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@UA^�SL�a�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@UA^�SL�a�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@UA^�SA^�a�"s��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@UA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@UA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@VA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@VA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@VA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@VA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@VA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@VA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@VA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@VA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@VA^�SA^�a�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�<VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�<VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�<VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�<VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�<VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�<VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�f�8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�f�8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�f�8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�f8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� �d�dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� �d� dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� �d� dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� �d� dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� �d� dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� �d� dcQ�t B(e1't   �� 	   � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� �d� dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� �d� dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� � d�$dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f8VA^�SA^�a.�3��T0 k� � d�$dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� � d�$dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� � d�$dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� � d�$dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� � d�$dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� � d�$dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� � d�$dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� �$d�(dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� �$d�(dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� �$d�(dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� �$d�(dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� �$d�(dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� �$d�(dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� �$d�(dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a.�3��T0 k� �(d�,dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a�3��T0 k� �(d�,dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a�3��T0 k� �(d�,dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a�3��T0 k� �(d�,dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a�3��T0 k� �(d�,dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a�3��T0 k� �(d�,dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a�3��T0 k� �(d�,dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f/8VA^�SA^�a^�3��T0 k� �(d�,dcQ�t B(e1't   ��    � �� �o�A���N�� "���Y|?��[/dDEo<[L 4u_+�3��T0 k� �7��;�cQ�t B(e1't   ��    � �� �o�A���N�� "���Y|?��]/`DEo8\L 0u_'�3��T0 k� �3��7�cQ�t B(e1't   ��    � �� �k�A���N�� "���Y|?��^/\CEo8\L ,u_'�3��T0 k� �3��7�cQ�t B(e1't   ��    � �� �k�A���Nߋ�"���Y|?��`/\CEo8]L $u_'�3��T0 k� �/��3�cQ�t B(e1't   ��    � �� �k�A���Nߋ�!���Y|?��a/XCEo4^L  u_'�3��T0 k� �+��/�cQ�t B(e1't   ��    � �� �g�A���Nߌ�!���Y|?��b/TBE_4^L u_#�3��T0 k� �'��+�cQ�t B(e1't   ��    � �� �g�A���Nߌ�!���Y|?��d/TBE_0_L u_#�3��T0 k� �#��'�cQ�t B(e1't   ��    � �� �c�A���Nی�!���Y|?��e/PBE_,`L u#�3��T0 k� ���#�cQ�t B(e1't   ��    � �� �c�A���Nی�!���Y|?��e/LAE_,`L u#�3��T0 k� ����cQ�t B(e1't   ��    � �� �c�A���Nی� ���Y|?��f/LAE_(aL v�3��T0 k� ����cQ�t B(e1't   ��    � �� �_�A���Nۍ� ���Y|?��f/HAE_$aL w�3��T0 k� ����cQ�t B(e1't   ��    � �� �_�A���N׍� ���a�?��g/DAE_ bL  x�3��T0 k� ����cQ�t B(e1't   ��    � �� �_�A���N׍� ���a�?��g/D@E_bL  x�3��T0 k� ����cQ�t B(e1't   ��    � �� �[�A���N׍� ���a�?��h/@@E_cL/�y�3��T0 k� ����cQ�t B(e1't   ��    � �� �[�A���N׍� ���a�?��h/@@E_dL/�y�3��T0 k� ����cQ�t B(e1't   ��    � �� �[�A���N׍����a�?��i/<?EOdL/�z�3��T0 k� ����cQ�t B(e1't   ��    � �� �W�A���Nӎ����a�?��i/8?EOdL/�{�3��T0 k� �����cQ�t B(e1't   ��    � �� �W�A���Nӎ����a�?��i/8?EOeL/�{�3��T0 k� �����cQ�t B(e1't   ��    � �� �W�A���Nӎ����a�?��j/4?EOeL/�|�3��T0 k� ������cQ�t B(e1't   ��    � �� �S�A���Nӎ����a�?��j/4>EO eL/�}�3��T0 k� ������cQ�t B(e1't   ��    � �� �S�A���Nώ����a�?��k/0>L��fL/�}�3��T0 k� ������cQ�t B(e1't   ��    � �� �S�A���Nώ����a�?��k/0>L��fL/�~/�3��T0 k� ������cQ�t B(e1't   ��    � �� �O�A���NϏ����Y|?��k/,>L��fL/�~/�3��T0 k� ������cQ�t B(e1't   ��    � �� �O�A���NϏ����Y|?��l/,=L��gL/�/�3��T0 k� ������cQ�t B(e1't   ��    � �� �O�A���NϏ����Y|?��l/(=L��gL/�/�3��T0 k� ������cQ�t B(e1't   ��    � �� �K�A���Nˏ����Y|?��m/(=L��gL/Ԁ/�3��T0 k� ������cQ�t B(e1't   ��    � �� �K�A���Nˏ����Y|?��m/$=L��hL/Ѐ/�3��T0 k� ������cQ�t B(e1't   ��    � �� �K�A���Nˏ����Y|?��m/$=L��hL/�/�3��T0 k� ������cQ�t B(e1't   ��    � �� �K�A���Nˏ����Y|?��n/ <L��hL/�/�3��T0 k� ������cQ�t B(e1't   ��    � �� �G�A���Nː����Y|?��n/ <M�hL/�/�3��T0 k� ������cQ�t B(e1't   ��    � �� �G�A���Nː����Y|?��n/<M�iL/�/�3��T0 k� ������cQ�t B(e1't   ��    � �� �G�A���Nǐ����Y|?��o/<M�iL�~/�3��T0 k� ������cQ�t B(e1't   ��    � �� �G�A���Nǐ����Y|?��o/<M�iL�~/�3��T0 k� ������cQ�t B(e1't   ��    � �� �C�A���Nǐ����Y|?��o/;M�iL�~/�3��T0 k� ������cQ�t B(e1't   ��   � �� �C�A���Nǐ����Y|?��p/;M�jL�~/�3��T0 k� ������cQ�t B(e1't   ��    � �� �C�A���Nǐ����Y|?��p/;M�jL�~/�3��T0 k� ������cQ�t B(e1't   ��   � �� �C�A���Nǐ����Y|?��p/;M�jL�}/�3��T0 k� ������cQ�t B(e1't   ��    � �� �?�A���NÑ����Y|?���q;M�jC�}/�3��T0 k� ������cQ�t B(e1't   ��    � �� �?�A���NÑ����Y|?���q:L��kC�}/�3��T0 k� ������cQ�t B(e1't   ��    � �� �?�A���NÑ����Y|?���q:L��kC�}/�3��T0 k� ������cQ�t B(e1't   ��    � �� �?�A���NÑ����Y|?���r:L��kC�|/�3��T0 k� ������cQ�t B(e1't   ��    � �� �;�A���NÑ����Y|?���r:L��kC�|/�3��T0 k� ������cQ�t B(e1't   ��    � �� �;�A���NÑ����Y|?���r:L��lC�|/�3��T0 k� ������cQ�t B(e1't   ��    � �� �;�A���N������Y|?���r�:L��lC�|/�3��T0 k� ������cQ�t B(e1't   ��    � �� �;�A���N������Y|?���s�9L��lL�|/�3��T0 k� ������cQ�t B(e1't   ��    � �� �7�A���N������Y|?���s� 9L��lL�{/�3��T0 k� ������cQ�t B(e1't   ��    � �� �7�A���N������Y|?���t� 9EN�mL�{/�3��T0 k� ������cQ�t B(e1't   ��    � �� �7�A���N������Y|?���t^�9EN�mL�{/�3��T0 k� ������cQ�t B(e1't   ��    � �� �7�A���N������Y|?���t^�9EN�mL�{/�3��T0 k� ������cQ�t B(e1't   ��    � �� �3�A���N������Y|?���t^�8EN�mL�{/�3��T0 k� �� �� cQ�t B(e1't   ��   � �� �3�A���N������Y|?���t^�8EN�mL�z/�3��T0 k� ����cQ�t B(e1't   ��   � �� �3�A���N������Y|?���u^�8E>�lL�z/�3��T0 k� ����cQ�t B(e1't   ��    � �� �3�A���N������Y|?���uN�8E>�lL�z/�3��T0 k� ����cQ�t B(e1't   ��    � �� �3�A���N������Y|?���uN�8E>�lL|z.��3��T0 k� ����cQ�t B(e1't   ��    � �� �3�A���N������Y|?�?�uN�8E>|lLxz.��3��T0 k� �|��cQ�t B(e1't   ��    � �� �/�A���N������Y|?�?�uN�8E>xkLtz.��3��T0 k� �x�|cQ�t B(e1't   ��    � �� �/�A���N������Y|?�?�uN�9L�tkLty.��3��T0 k� �x�|cQ�t B(e1't   ��    � �� �/�A���N������Y|?�?�t>�9L�pkL/py.��3��T0 k� �t�xcQ�t B(e1't   ��   � �� �/�A���N������Y|?�?�t>�9L�pjL/ly.��3��T0 k� �p�tcQ�t B(e1't   ��    � �� �/�A���N������Y|?�?�t>�9L�ljL/hy.��3��T0 k� �l�pcQ�t B(e1't   ��    � �� �/�A���N������Y|?�?�t>�:L�hjL/hy.��3��T0 k� �h�lcQ�t B(e1't   ��    � �� �+�A���N������Y|?�?�t>�:L�diL/dy��3��T0 k� �h�lcQ�t B(e1't   ��    � �� �+�A���N������Y|?�?�t>�:L�diL/`y��3��T0 k� �d�hcQ�t B(e1't   ��    � �� �+�A���N������Y|?�?�t>�;L�`iL/`x��3��T0 k� �`	�d	cQ�t B(e1't   ��    � �� �+�A���N������Y|?�?�t>�<L�\hL/\x��3��T0 k� �\
�`
cQ�t B(e1't   ��    � �� �+�A���N������Y|?�?�t.�<L�XhL/Xx��3��T0 k� �\
�`
cQ�t B(e1't   ��    � �� �+�A���N������Y|?�?�s.�=L�XhL/Xx��3��T0 k� �X�\cQ�t B(e1't   ��    � �� �'�A���N������Y|?�?�s.�=L�TgL/Tx^��3��T0 k� �T�XcQ�t B(e1't   ��    � �� �'�A���N������Y|?�?�s.�>L�PgL/Px^��3��T0 k� �P�TcQ�t B(e1't   ��    � �� �'�A���N������Y|?�?�s.�?L�PgL/Px^��3��T0 k� �L�PcQ�t B(e1't   ��    � �� �'�A���N������Y|?�?�s.�?L�LgL/Lw^��3��T0 k� �L�PcQ�t B(e1't   ��    � �� �'�A���N������Y|?�?�s.�@L�HfL/Lw^��3��T0 k� �H�LcQ�t B(e1't   ��    � �� �'�A���N������Y|?�O�s.�AL�HfL/Hw^��3��T0 k� �D�HcQ�t B(e1't   ��   � �� �'�A���N������Y|?�O�s.�BL�DfL/Dw^��3��T0 k� �@�DcQ�t B(e1't   ��    � �� �'�A���N������Y|?�O�s.�CL�@fL/Dw^��3��T0 k� �@�DcQ�t B(e1't   ��    � �� �#�A���N������Y|?�O�s��DL�@eL/@w^��3��T0 k� �<�@cQ�t B(e1't   ��    � �� �#�A���N������Y|?�O�s��EL�<eL/@w^��3��T0 k� �8�<cQ�t B(e1't   ��    � �� �#�A���N������Y|?�O�s��EL�8eL/<w^��3��T0 k� �4�8cQ�t B(e1't   ��    � �� �#�A���N������Y|?�O�r��FL�8eL/<w^��3��T0 k� �4�8cQ�t B(e1't   ��    � �� �#�A���N������Y|?�O�r��GL�4dL/8v^��3��T0 k� �0�4cQ�t B(e1't   ��    � �� �#�A���N������Y|?�O�r.�HL�4dL/8v^��3��T0 k� �,�0cQ�t B(e1't   ��    � �� �#�A���N������Y|?�O�r.�IL�0dL/4v^��3��T0 k� �(�,cQ�t B(e1't   ��    � �� �#�A���N������Y|?�O�r.�JL�0dL/4v^��3��T0 k� �(�,cQ�t B(e1't   ��    � �� ��A���N������Y|?�O|r.�LE>,cL/0v^��3��T0 k� �$�(cQ�t B(e1't   ��    � �� ��A���N������Y|?�O|r.�ME>,cL/0v^��3��T0 k� � �$cQ�t B(e1't   ��    � �� ��A���N������Y|?�Oxr.�NE>(cL/,v^��3��T0 k� �� cQ�t B(e1't   ��    � �� ��A���N������Y|?�Oxr�OE>(bL/,v^�3��T0 k� �� cQ�t B(e1't   ��    � �� ��A���N������Y|?�Otr�PE>$bL/(v^�3��T0 k� ��cQ�t B(e1't   ��    � �� ��A���N������Y|?�Otr�QL�$aL/(v^�3��T0 k� ��cQ�t B(e1't   ��   � �� ��A���N������Y|?�Opr�RL�$aL/$u^�3��T0 k� ��cQ�t B(e1't   ��    � �� ��A���N������Y|?�Opr�SL� aL/$u^�3��T0 k� ��cQ�t B(e1't   ��    � �� ��A���N������Y|?�Olq��TL� `L/$u^�3��T0 k� ��cQ�t B(e1't   ��   � �� ��A���N������Y|?�Olq��UL� `L/ u^�"s��T0 k� ��cQ�t B(e1't   ��    � �� ��A���N������Y|?�Olq��VL�`L/ u^�"s��T0 k� ��cQ�t B(e1't   ��    � �� ��A���N������Y|?�Ohq��WL�_L/u^�"s��T0 k� ��cQ�t B(e1't   ��    � �� ��A���N������Y|?�Ohq��XL�_L/u^�"s��T0 k� � �cQ�t B(e1't   ��    � �� ��A���N������Y|?�Odq�YL�^L/u^�"s��T0 k� ��� cQ�t B(e1't   ��    � �� ��A��N������Y|?�Odq�ZL�^L/u^�"s��T0 k� ��� cQ�t B(e1't   ��    � �� ��A��N������Y|?�O`q�[L�^Lu^�"s��T0 k� ����cQ�t B(e1't   ��    � �� ��A��N������Y|?�O`q�\L�]Lu^�"s��T0 k� ����cQ�t B(e1't   ��    � �� ��A��N������Y|?�O`q�]L�]Lu^�"s��T0 k� �� �� cQ�t B(e1't   ��    � �� ��A��N������Y|?�O\q��^L�]Lt^�"s��T0 k� ��!��!cQ�t B(e1't   ��    � �� ��A��N������Y|?�O\q��^L�\Lt^�"s��T0 k� ��!��!cQ�t B(e1't   ��    � �� ��A��N������Y|?�OXq��_L�\Lt^�3��T0 k� ��"��"cQ�t B(e1't   ��    � �� ��A��N������Y|?�OXq��`L�\C�t^�3��T0 k� ��"��"cQ�t B(e1't   ��    � �� ��A��N��� ���Y|?�OXq��`L�\C�t^�3��T0 k� ��#��#cQ�t B(e1't   ��    � �� ��A��N��� ���Y|?�OTq��aL�[C�t^�3��T0 k� ��$��$cQ�t B(e1't   ��    � �� ��A��N��� ���Y|?�OTq��aL�[C�t^�3��T0 k� ��$��$cQ�t B(e1't   ��    � �� ��A��N��� ���Y|?�OTq��bL�[C�t^�3��T0 k� ��%��%cQ�t B(e1't   ��    � �� ��A��N��� ���Y|?�OPp��bL�ZEOt^�3��T0 k� ��%��%cQ�t B(e1't   ��    � �� ��A��N��� ���Y|?�OPp��bL�ZEO t^�3��T0 k� ��&��&cQ�t B(e1't   ��    � �� ��A��N��� ���Y|?�OPp��cL�ZEN�t^�3��T0 k� ��'��'cQ�t B(e1't   ��    � �� ��A��N��� ���Y|?�OLp~�cL�ZEN�s^�3��T0 k� ��'��'cQ�t B(e1't   ��    � �� ��A��N��� ���Y|?�?Lp~�cL�YEN�s^�3��T0 k� ��(��(cQ�t B(e1't   ��    � �� ��A��N��� ���Y|?�?Lp~�cL�YEN�s^�"���T0 k� ��(��(cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?Hp cE.YE>�s^�"���T0 k� ��)��)cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?HpcE.XE>�s^�"���T0 k� ��*��*cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?HpbE.XE>�s^�"���T0 k� ��*��*cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?DpbE.XE>�r^�"���T0 k� ��+��+cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?DpbE.WE>�r^�"���T0 k� ��+��+cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?DpaEWE>�r^�"���T0 k� ��,��,cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?@p_aEVE>�q^�"���T0 k� ��,��,cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?@p_aEVE.�q^�"���T0 k� ��-��-cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?<o_ `EUE.�p^�"���T0 k� ��.��.cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?<o_$`EUE.�p^�"���T0 k� ��.��.cQ�t B(e1't   ��    � �� ��A��N���!���Y|?�?<o_(_B�UE.�o^�3��T0 k� ��/��/cQ�t B(e1't   ��    � �� ��A��N���"���Y|?�?<o_,_B�TE.�n^�3��T0 k� ��/��/cQ�t B(e1't   ��    � �� ��A��N���"���Y|?�?8n_,^B�TB��n^�3��T0 k� ��0��0cQ�t B(e1't   ��    � �� ��A��N���"���Y|?�?8n_0^B�TB��m^�3��T0 k� ��1��1cQ�t B(e1't   ��    � �� ��A��N��� "���Y|?��4n_4]B�SB��l^�3��T0 k� ��1��1cQ�t B(e1't   ��    � �� ��A��N��� "���Y|?��4n_8]B�SB��l^�3��T0 k� ��2��2cQ�t B(e1't   ��    � �� ��A��N��� "���Y|?��0m_<\B�RB��k^�3��T0 k� ��2��2cQ�t B(e1't   ��    � �� ��A��N��� "���Y|?��,m_<\L�RB��j^�3��T0 k� ��3��3cQ�t B(e1't   ��    � �� ��A��N��� "���Y|?��,m_@[L� RB��i^�3��T0 k� ��3��3cQ�t B(e1't   ��    � �� ��A��N��� "���Y|?��(l_D[L� QB��i^�3��T0 k� ��4��4cQ�t B(e1't   ��    � �� ��A��N��� "���Y|?��$loDZL�$QB��h^�3��T0 k� ��5��5cQ�t B(e1't   ��    � �� ��A��N��� "���Y|?��$koHZL�(QB��g^�3��T0 k� ��5��5cQ�t B(e1't   ��    � �� ��A��N��� "���Y|?�� koLYL�(QC�f^�3��T0 k� ��6��6cQ�t B(e1't   ��    � �� ��A��N��� #���Y|?��joPYL�,PC�e^�3��T0 k� ��6��6cQ�t B(e1't   ��    � �� ��A��N��� #���Y|?��ioPXL�0PC�d^�3��T0 k� ��7��7cQ�t B(e1't   ��    � �� ��A��N��� #���Y|?��hoTXL�0PC�c^�3��T0 k� ��7��7cQ�t B(e1't   ��    � �� ��A��N��� #���Y|?��hoXWL�4OC�b^�3��T0 k� ��8��8cQ�t B(e1't   ��    � �� ��A��N��� #���Y|?��goXWL�8OC�a^�3��T0 k� �|8��8cQ�t B(e1't   ��    � �� ��A��N��� #���Y|?��go\VL�8OC�`^�3��T0 k� �|9��9cQ�t B(e1't   ��    � �� ��A��N��� #���Y|?��fo\VL�<NC�`^�3��T0 k� �x:�|:cQ�t B(e1't   ��    � �� ��A��N��� #���Y|?��fo`VL�@NC�_^�3��T0 k� �x:�|:cQ�t B(e1't   ��    � �� ��A��N���$#���Y|?��fodUL�@NC�^^�3��T0 k� �t;�x;cQ�t B(e1't   ��    � �� ��A��N���$#���Y|?��fodUL�DNC�^^�3��T0 k� �p;�t;cQ�t B(e1't   ��    � �� ��A��N���$#���Y|?��eohTL�DMC�]^�3��T0 k� �p<�t<cQ�t B(e1't   ��    � �� ��A��N���$#���Y|?��eohTL�HMC�\^�3��T0 k� �l<�p<cQ�t B(e1't   ��    � �� ��A��N���$#���Y|?��eolTL�HMC�\^�3��T0 k� �h=�l=cQ�t B(e1't   ��    � �� ��A��N���$#���Y|?��eopSL�LMC�[^�3��T0 k� �h=�l=cQ�t B(e1't   ��    � �� ��A��N���$#���Y|?��dopSL�PLC�[^�3��T0 k� �d>�h>cQ�t B(e1't   ��    � �� ��A��N���$#���Y|?��dotSL�PLC�[^�3��T0 k� �`?�d?cQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��dotRL�TLC�Z^�3��T0 k� �`?�d?cQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��doxRL�TLC�Z�3��T0 k� �\@�`@cQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��doxQL�XKC�Z�3��T0 k� �X@�\@cQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do|QL�XKC�Z�3��T0 k� �XA�\AcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do|QL�\KC�Y�3��T0 k� �TA�XAcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do�PL�\KC.�Y�3��T0 k� �TB�XBcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do�PB�`JC.�Y�3��T0 k� �PB�TBcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do�PB�`JC.�Y�3��T0 k� �LC�PCcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do�OB�dJC.�Y�3��T0 k� �LC�PCcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do�OB�hJC.�Y�3��T0 k� �HD�LDcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do�OB�hJ@n�Y�3��T0 k� �DD�HDcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do�OB�lI@n�Y�3��T0 k� �DE�HEcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do�NEpI@n�Y�3��T0 k� �@F�DFcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do�NEtI@n�Y�3��T0 k� �<F�@FcQ�t B(e1't   ��    � �� ��A��N���$$���Y|?��do�NExI@n�Y�3��T0 k� �<G�@GcQ�t B(e1't   ��    � �� ��A��N���($���Y|?��do�ME|IK��Y.�3��T0 k� �8G�<GcQ�t B(e1't   ��    � �� ��A��N���($���Y|?��do�ME�HK��Y.�3��T0 k� �8H�<HcQ�t B(e1't   ��    � �� ��A��N���($���Y|?��do�ME�HK��Y.�3��T0 k� �4H�8HcQ�t B(e1't   ��    � �� ��A��N���($���Y|?��do�ME�HK��Y.�3��T0 k� �0I�4IcQ�t B(e1't   ��    � �� ��A��N���($���Y|?��do�LE��HK��Y.�3��T0 k� �0I�4IcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?��do�LE��HK��Y.�3��T0 k� �,J�0JcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?��do�LE��HK��Y.�3��T0 k� �,J�0JcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?��d_�LE��HK��Y.�3��T0 k� �(K�,KcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d_�KE��HK��Y.�3��T0 k� �$K�(KcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d_�KE��HK��Y.�3��T0 k� �$L�(LcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d_�KE��HK��Y.�3��T0 k� � L�$LcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d_�KE��HK��Y.�3��T0 k� �M� McQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d_�JE��IK��Y.�3��T0 k� �M� McQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d�JE��IK��Y.�3��T0 k� �N�NcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d�JE��IK��Y.�3��T0 k� �N�NcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d�IE��IK��Z.�3��T0 k� �O�OcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d�IE��IK��Z.�3��T0 k� �P�PcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d�IE��IK��Z.�3��T0 k� �P�PcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_do�HE~�IK��Z.�3��T0 k� �Q�QcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_do�HE~�IK��Z.�3��T0 k� �Q�QcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_do�GE~�JK��[.�3��T0 k� �R�RcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_do�GE~�JK��[.�3��T0 k� �R�RcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_do�FE~�JK��[.�3��T0 k� �S�ScQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d_�FI��JK��[.�3��T0 k� � S�ScQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d_�EI��JK��\.�3��T0 k� � T�TcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d_�EI��KK��\.�3��T0 k� ��T� TcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d_�DI��KK��\.�3��T0 k� ��U� UcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_d_�DI� KK��\.�3��T0 k� ��U��UcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_dO�DI�KK��\.�3��T0 k� ��V��VcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_dO�CI�KK��].�3��T0 k� ��V��VcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_dO�CI�KK��].�3��T0 k� ��W��WcQ�t B(e1't   ��    � �� ��A��N���(%���Y|?�_dO�CI�KK��].�3��T0 k� ��W��WcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_dO�CI�KK��].�3��T0 k� ��X��XcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d��CEKK��].�3��T0 k� ��X��XcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d��CEKK��^.�3��T0 k� ��Y��YcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d��CEKK��^.�3��T0 k� ��Y��YcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d��CEKK��^.�3��T0 k� ��Z��ZcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d��CELK��^.�3��T0 k� ��Z��ZcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d��CEo LK��^.�3��T0 k� ��[��[cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d��CEo LK��_.�3��T0 k� ��[��[cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d��CEo$MK��_.�3��T0 k� ��\��\cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d��DEo$MK��_�3��T0 k� ��\��\cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d��DEo$NK��_�3��T0 k� ��]��]cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�|DD?(NK��_�3��T0 k� ��]��]cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�|ED?(OK��_�3��T0 k� ��^��^cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�xED?(PK��_�3��T0 k� ��^��^cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�tED?(PK��_�3��T0 k� ��_��_cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�pFD?(QK��`^�3��T0 k� ��_��_cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�lFD?(QK��`^�3��T0 k� ��`��`cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�hGD?(QK��`^�3��T0 k� ��`��`cQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�dGD?(RK��`^�3��T0 k� ��a��acQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�`HD?(RK��`^�3��T0 k� ��a��acQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�\HD?(RK��`^�3��T0 k� ��b��bcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�\HD?(SK��`^�3��T0 k� ��b��bcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�XHD?$SK��`^�3��T0 k� ��c��ccQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�XHDO$TK��a^�3��T0 k� ��c��ccQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�XHDO$TK��a^�3��T0 k� ��d��dcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�THDO$TK��a^�3��T0 k� ��d��dcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�TIDO$TK��a^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�TIDO$TK��a^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_d�TIDO$TK��a^�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_e�TIDO$TK��a^�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_e�TIDO$T@��a^�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_e�TIDO$T@��a^�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_e�TIDO$T@��a^�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_e�TIDO$T@��a^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_e�TIA�$T@��a^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_e�TIA�$T@��a^�3��T0 k� ��i��icQ�t B(e1't   ��    � �� ��A��N���,&���Y|?�_e�TIA�$T@��a^�3��T0 k� ��i��icQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�TIA�$T@��a^�3��T0 k� ��i��icQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�TIA�$T@��a^�3��T0 k� ��i��icQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�TIA_$T@��a^�3��T0 k� ��i��icQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�TIA_$T@��a^�3��T0 k� ��i��icQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�TIA_ T@��a^�3��T0 k� ��i��icQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�PIA_ T@n�a^�3��T0 k� ��i��icQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�PIA_ T@n�a^�3��T0 k� ��i��icQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�PIA_ T@n�a^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�PIA_ T@n�a^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�PIA_ U@n�a^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���,'���Y|?�e�LIA_ UB��`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�e�LIA_ UB��`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�e�LIA_ UB��`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�e�LIA_ UB��`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/e�LIA_ UB��`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/e�LIA_UB��`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/e�LIA_UB��`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/e�LJA_UB��`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/e�LJA_U@n�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/e�LJA_U@n�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/e�LJA_U@n�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/e�LJA_U@n�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/e�LJA_U@n�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/e�LJA_U@n�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/e�LJA_U@n�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/e�LJA_U@n�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/e�LKA_U@n�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/e�LKA_U@n�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/e�LKMU@�`^�3��T0 k� ��h��hcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/e�LKMU@�`^�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/e�LKMU@�`^�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/f�LKMU@�`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/f�LKMV@�`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/f�LKMVB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/f�LKMVB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�LKMVB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�LKMVB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�LKMVB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�LLM/VB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�LLM/VB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/g�LLM/WB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/g�LLM/WB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/g�LLM/WB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/g�LLM/WB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/g�LLM/WB��`�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/g�LLM/WB��`.�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/g�LLM/W@�`.�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/g�LLMW@�`.�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/h�LLMW@�`.�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/h�LLMW@�`.�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/h�LLMW@�`.�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/h�LLMWBN�`.�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/h�LLMWBN�`.�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/h�LLMWBN�`.�3��T0 k� ��g��gcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�/h�LLMWBN�`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�hLLMWBN�`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���a�?�hLLMWBN�`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�iLLMWBN�`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�iHLMWBN�`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�iHLA_WBN�`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�iHLA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�iHLA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��iHMA_WA��`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��iHMA_WA^�`.�3��T0 k� ��f��fcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��iHMA_WA^�`.�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��hHMA_WA^�`�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��hHMA_WA^�`�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��hHMA_WA^�`�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��gHMA_WA^�`�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��gHMA_WA^�`�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��gHMA_VA^�`�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��gHMA_VA^�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��gHMA_VA^�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��fHMMVA^�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��fHMMVA^�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMMVA^�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMMUA^�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMMUL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�LMMUL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�LMMUL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�LMMUL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�LMMTL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��fLMMTL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��fLMM/TL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��fLMM/TL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��fLMM/TL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��fLMM/TL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�LMM/SL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMM/SL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMM/SL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMM/SL�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMM/SL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMMSL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMMSL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMMSL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMMSL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HMMSL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HNMSL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?��f�HNMSL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f�HNMSL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f�HOMSL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f�HOMSL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f�HOM SL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f�DPM SL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�_f�DPM SL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@QM SL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@QM SL.�`^�3��T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RM SL.�`^�"���T0 k� ��e��ecQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RM SL.�`^�"���T0 k� ��d��dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RM SL.�`^�"���T0 k� ��d��dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RM SL.�`^�"���T0 k� ��d��dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RM SL.�`^�"���T0 k� ��d��dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RM SL.�`^�"���T0 k� ��d��dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RM SL.�`^�"���T0 k� ��d� dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RM SL.�`^�"���T0 k� ��d� dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RM SL.�`^�"���T0 k� ��d� dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RA_ SL.�`^�"���T0 k� ��d� dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RA_ SL.�`^�"���T0 k� ��d� dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�f�@RA_ SL.�`^�3��T0 k� ��d� dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA_ SL.�`^�3��T0 k� ��d� dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA_ SL.�`^�3��T0 k� � d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA_ SL.�`^�3��T0 k� � d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA_ SL.�`^�3��T0 k� � d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA_ SL.�`^�3��T0 k� � d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA_ SL.�`^�3��T0 k� � d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA_ SL.�`^�3��T0 k� � d�dcQ�t B(e1't   ��    � �� ��A��N���0'���Y|?�/f�@RA_ SL.�`^�3��T0 k� � d�dcQ�t B(e1't   ��    � ��                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��. ]�)|){ � ������         ���B�    ������B�                        � =          ^p     ���   0

           ����        � ި    ���� ި                      ���         �     ���   (
           ����   $ $       ��^    ������^           
         ���         �     ���   8
�          '�C    H	     �fV     '�C�fV                       �$          �     ���   (
          ����     	   .�(�    �����(�                     ���H          �     ���   P	B 
         ��a� ��
      B�    ��a��                             ����                 ���    8		 1 	             f�    
	  V��t�     f���t�                      0	 Z��         �     ��@   8
(
          VO�  � �
	  j�ν�     VO�����      ��              	 Z��          �    ��`   @          S��   	    ~����     S������                     	 Z��         �     ��@    

'           a   
	   �����     a����                   .	 Z��         	 �  �  ��@   8
	          ���a    
	   �����    ���a����                     <  Z��         
 &P     ��H  X
         ��<� ��
     � ��W    ��<� ��W                              ���/              y  ��@    0 0                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          du  ��        ��
�H     du�
�      �                   x                j  �   �
   �                          d    ��       ��       d  �           "                                                  �                         �� ����(����������� ����
�         
  	      
     ��x ;�D       �� �t� �� u� � n` �$ n� �D n� �d n� �� o  <�  n@ �� u� � u� �$ v  �D v  �d v@ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0� ���� � � }`���� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �������� �� ?  ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"     "�j��   * �
� �  �  
� ����  ��     ���  �   ��    ��     ���      ����  ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �      �� � ���        � � � ���        �        ��        �        ��        �  
   ��     d, e��        ��                         �w� $ 		�� �                                    �                 ����           �������%��   ����               28 Steve Larmer lny    5:01                                                                        3  3     �B� �/ B� � �C � � C � �k�W k�W �c� � c� � �	k~I � 
k�I �cV\ � c^d �cjK � cr[ � csC � ctF � cuL � cvN �J� � � J� �:"� �: "� �*"� �**� �"� � "� � �� � � 
� �"� � "� � �� � � 
� � � 
� � � 
� �#"� � $"� � �%� � � 
� � � 
� � � 
� � �)"� y � *"� � �+� y � 
� � � 
� � �.� � � 
� � � 
� � �1� � � 
� �X  "K �X  "K �@  "K �X 6"K uX  "K �X  "G wX  "H �8 :"L �P ;"R �X  "K �=*2|7>*:lG  *Gl                                                                                                                                                                                                                         p� P @       �     @ 
             l P E n  ��         
            �������������������������������������� ���������	�
��������                                                                                          ��    ��~!�� ��������������������������������������������������������   �4, @   ��@#� �v��т ��                                                                                                                                                                                                                                                                                                                                           �L                                                                                                                                                                                                                                                   4    7    � �  L�J      �                             ������������������������������������������������������                                                                                                                                     	      �    �              �          ��                 	 	 ��������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� ���������������������                                  -    -    ��  4�J                                     ������������������������������������������������������                                                                                                                                         �  �     �        �          ��               	 
     ������ ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ������           x                                                                                                                                                                                                                                                           
                              	                   �             


           �   }�         ������������   	  '�����������������������������    ��������������������  '}����������������������������                                                       N�                        �ww�ww333wwwwwwww�ww�ww�ww�ww333wwww 0 I =                                 � tLq �\                                                                                                                                                                                                                                                                                    E)h1p  �                             W             m                                          ��                                                                                                                                                                                                                                                                                                                                                                  
 �  � ��  � ��  � 2��  � 2��  � _��  ��H�6���������������������������������G������        <        �w ~           �   & AG� �  k   
              �                                                                                                                                                                                                                                                                                                                                      p I N   �                       !��                                                                                                                                                                                                                            Y��   �� �� ��      �� 4      ��������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� ��������������������������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ������             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    ?   #   D      d                       4     �   �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��     �� p���� ���� p � �N��   `d     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@     B 
df ��  B 
df �$ ^$   2 � ��� �� � ���  � �d �  ��d  �      �  ��   �������2����  g���        f ^�         �� "             ������2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                                    �����   �   �   �   ����                                     	�  		  	 � 	 	 	   	   	   	   	  ��                  ��   	   	   	   	   	   	 	 	 � 		  	�                 �   	    �   	    �   	    �   	   	   �  	   �  	   �  	   �                                                       �����   �   �   �   ����                                     
�  

  
 � 
 
 
   
   
   
   
  ��                  ��   
   
   
   
   
   
 
 
 � 

  
�                 �   
    �   
    �   
    �   
   
   �  
   �  
   �  
   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   """ "!   " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  "!    " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       """ "!   " ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                      �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                             �� ��������p��}`     �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��  ��  ��� �   ��  ���   �                       � ���� ��   � � �                                                                                                                                  �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �   �   "   "   "  !�    ��                              �                        ���� ��� ����            �����                            �   �                        �   ��  �   ��   �       �                                                                                                                                      �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �      �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                     �          ��                                 � ���� ��   � � �           � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         ̰ �� ̻ {�����vz� w��  ��  ��  ̘  	�  
� "��,̻�"�� "#3  34  D  
�  �  " "" """ ! ��  ��                               ˹� �ɩ ��� �͋ ��� ��� ��̀��Ȑ���лܹнȝ0ݙ�@43�PCD�@@E�@ E�@ U�� H�  K�  �   ��    �� "�" ���                          �  �   ��  �  ��                �   �   �   "   "   "  !�    ��                                 �   �                      �������  ���    �    �  �  ��  �   �   �         �       �                        �   ��  ���  � �    �                                                                                                                                       �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                        �   �   �    "�"�����   �� �          ����   �       �                                   �    ���  ��                    ��  ��  ���  �  �  �   �   ��  �                            �   ���                            �   �                                                                                                    �� ̽ �� �� w} 
�� ��� ����̙������ ��� ��� ����̻�������EUUUUEUDUD0�C��� �� �� �� ؠ ۰ ��(� "�����     �   �  �     �  ��  ��  ��� ˸� ��� ����؛� ۻ������ �  �; J�� D�� D�� D;� �۰ ��� ��  ��  ��  �۰ �ً ����"� �   �                    �   �   �   �   �   �  �  "  �         �   �   �   �            � ��  ���  �  � �                     ��� ����                                �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw  ��  �   ��  �                             �  �˰ ��� �wp ���                                                                                                                                                                      �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��                        � ��                  �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  �   �   �   �   �       �     �"  "  �   "                                    �   �   �            �� �� �� g} �� vw                      �          ���� �                                           �   ���                            �   �                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw     �  �  ��  �   �   �                         ���                                                                                                                                                                             �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw    �  �  �� �� �   �                            � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                          �� ̻ ��˛��  �� �˚̻���ۚ����I���䘼�^���^�٘�:�^�� ^�� D�( �) �) �) ��) ˹� ț�+��,��,����  �𫝝 ��� �ɍ ��ݨ��ډ�݊�� ��D@ �D�  J�� ݩ� ��� �ۻ �ک �ڹ�ɻ��̸���������� ����������            �   ��  ��  ��  ��  ��                                          �� ��� ��� ��  �                         �   �                    �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww���������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqB� �/ B� � �C � � C � �k�W k�W �c� � � c� � �	k~I � 
k�I �cV\ � c^d �cjK � cr[ � csC � ctF � cuL � cvN �J� � � J� �:"� �: "� �*"� �**� �"� � "� � �� � � 
� �"� � "� � �� � � 
� � � 
� � � 
� �#"� � $"� � �%� � � 
� � � 
� � � 
� � �)"� y � *"� � �+� y � 
� � � 
� � �.� � � 
� � � 
� � �1� � � 
� �X  "K �X  "K �@  "K �X 6"K uX  "K �X  "G wX  "H �8 :"L �P ;"R �X  "K �=*2|7>*:lG  *Gl3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0�����������������������������������������#��<�Z�K�\�K��6�G�X�S�K�X� � � � � � � � �-�2�3�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������-�2�3� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������,�>�0� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                