GST@�                                                           N}     N�                                               
           � �      ��     � J� 2��������}�����    ����        Ȁ      #    ����                                d8<n    � �     � �  "Df��
���    
  ���D"��   " `  J  jF �   ffffffffff 
ff �   ffffffffff  ff  ��                                                                              ����������������������������������      ��    a bQb  411 c cc cc  	     
    	  
        Gg � (	 (                 pY$ 11"         8:=�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             n�  )!          == �����������������������������������������������������������������������������                                �          �   @  &   �   �                                                                                 'w w  1p1Y"$  )n!�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ��c@�`{D^����sK��SZ3�L0PA�_�@���\D �<�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;��c@�\{D^����sK��SZ3�L0PA�_�@���\D �<�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;��c@�\{D^����sK��SZ3�L0PA�_�@���\D �<�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;��c@�\|D^����sK��Rbs�L0PA�_�@���\D �<�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;��c@�X|D^����sK��Rbs�L0PA�_�@���\D �<�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;��b@�X|D^� ��sK��Rbs�L0PA�_�@���\C �<�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;��b@�X|D^���sK��Rbs�L0PA�c�@���\C �<�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;��b@�X|D^���sK��Rbs�L0PA�c�@���\C �<�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;��b@�T|D^���sK��Rbs�L0PA�c�@���\C �<�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;��b@�T|D^���sK��Rbs�L0PA�c�@���XC �<�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;��b@�T|Dn���sK��Rbs�L0PA�c�@���XC �<�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;��b@�T|Dn�	��sK��Qbs�L0PA�c�@���XC �<�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;��b@�T|Dn���rK��Qbs�L0PA�c�@���XC �<�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;|�b@�P|Dn���rK��Qbs�L0PA�c�@���XC �<�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;|�b@�P|Dn���rL�QZ3�L0PA�c�@���XC �<�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;|�a@�P|Dn���rL�PZ3�L0PA�c�@���XC �<�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;|�a@�P|Dn���qL�PZ3�L0PA�c�@���XC �<�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;|�`@�L}En���qL�PZ3�L0PA�c�@���XB �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�`@�L}En�\�pL�PZ3�L0PA�g�@���XB �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�`@�L}En�\�pL�PZ3�L0PA�g�@���XB �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�`@�L}En�\�pL�OZ3�L0PA�g�@���XB �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�`@�L}En�\�pL�OZ3�L0PA�g�@���XB �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�`@�L}En�\�pL�OZ3�L0PA�g�@���TB �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�_@�H}En�\�oL�OZ3�L0PA�g�@���TB �<#�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�_@�H}En�\�oL�NZ3�L,PA�g�@���TB �<#�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�_@�H}En�!\�oL�Nb��L,PA�g�@���TB �<#�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�_@�H}En�#\�oL�Nb��L,PA�g�@���TB �<#�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�_@�H}E^�%l�oL�Nb��L,OA�g�@���TB �<#�T0 k� ���#�P &�1D"3Q	E1 4#Q ��   � "�;|�_@�D}E^�'l�oL�Nb��L,OA�g�@���TB �<#�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�^@�D}E^�)l�oL�Mb��L,OA�g�@���TB �<'�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�^@�D}E^|*l�oL�Mb��L,OA�g�@���TB �<'�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�^@�D}E^t,l�oL�Mb��L,OA�g�@���TB �<'�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�^@�D}E^p.l�oL�Mb��L,OA�g�@���TA �<'�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�^@�D}E^h/l�nL�Mb��L,OA�g�@���TA �<'�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�^@�@}E^d1l�nL�Lb��L,OA�k�@���TA �<'�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�^@�@}E^\3l�nL�Lb��L,OA�k�@���TA �<'�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�^@�@~E^T4\�nL�LZ3�L,OA�k�@���TA �<+�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�^@�@~C�P6\�nL�LZ3�L,OA�k�@���TA �<+�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�^@�@~C�H7\�nL�LZ3�L,OA�k�@���PA #�<+�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�^@�@~C�@9\�nL�LZ3�L,OA�k�@���PA #�<+�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�^@�@~C�<:\�nL�KZ3�L,OA�k�@���PA #�<+�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��^@�<~C�4<\�nL�KZ3�L,OA�k�@���PA #�<+�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��^K�<~C�,=\�nL�KZ3�L,OA�h @���PA #�<+�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��^K�<~C�$?\�nL�KZ3�L,OA�h @���PA #�<+�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��^K�<~C�@\�nL�KZ3�L,OA�h @���PA #�</�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��^K�<~C�A��nL�KZ3�L,OA�h @���PA #�</�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��^K�<~C�C��nL�JZ3�L,OA�h @���PA #�</�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��^K�<~C�D��nL�JZ3�L,OA�h @���PA #�</�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;��^K�8~C��E��nL�JZ3�L,OA�h @���PA #�</�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;��^K�8~C��G��nL�JZ3�L,OA�h @Û�PA #�</�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;��^K�8~C��H��nL�JZ3�L,OA�h @Ú�PA #�</�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;\�^K�8~C��I��nL�JZ3�L,OA�h @Ú�PA #�</�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;\�^K�8~C��J��nL�JZ3�L,OA�h @Ú�PA #�</�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;\�^K�8~C��L��nL�IZ3�L,OA�l @Ú�PA #�<3�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;\�]K�8~C��M��nL�IZ3�L,OA�l @Ú�P@ #�<3�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;\�]K�8~C��N��nK��IZ3�L,OA�l@Ú�P@ #�<3�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;\�]K�8~C��O��mK��IZ3�L,OA�l@Ǚ�P@ #�<3�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;\�]K�4~C��P��mK��IZ3�L,OA�l@Ǚ�P@ #�<3�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;\�\K�4~C��Q��mK��IZ3�L,OA�l@Ǚ�P@ '�<3�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;\�\K�4~C��S��lK��IZ3�L,OA�l@Ǚ�P@ '�<3�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;\�\K�4D�T��lK��IZ3�L,OA�l@Ǚ�P@ '�<3�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;\�\K�4~D�U��lK��IZ3�L,OA�l@Ǚ�L@ '�<3�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;\�\K�4~D�V��lK��HZ3�L,OA�l@Ǚ�L@ '�<3�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;\�[K�4~D|W��lK��HZ3�L,OA�l@ǘ�L@ '�<3�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;\�[K�4}DtX��lA�HZ3�L,OA�l@ǘ�L@ '�<7�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;l�[K�4}LlY��kA�HZ3�L,OA�l@˘�L@ '�<7�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;l�[K�4}LdZ��kA�HZ3�L,OA�l@˘�L@ '�<7�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;l�ZK�4}L\[��kA�HZ3�L,OA�l@˘�L@ '�<7�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;l�ZK�4|LT\��kA�HZ3�L,OA�l@˘�L@ '�<7�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;l�ZK�4|LL]��kA\�HZ3�L,OA�l@˘�L@ '�<7�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;l�ZK�4|LD^��kA\�HZ3�L,OA�l@˗�L@ '�<7�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;l�YK�4|L<_��kA\�HZ3�L,OA�l@˗�L@ '�<7�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;l�YK�4|L4_��kA\�HZ3�L,OA�l@˗�L@ '�<7�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�YK�4{L,`��kA\�HZ3�L,OA�l@˗�L@ '�<7�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�YK�4{L$a��kA��HZ3�L,OA�l@ϗ�L@ '�<7�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�4{Lb��kA��HZ3�L,OA�l@ϗ�L@ '�<7�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�4{Lb��kA��HZ3�L,OA�l@ϗ�L@ '�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�4zLb��kA��HZ3�L,OA�l@ϗ�L@ '�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�4zLb��kA��HZ3�L,OA�p@ϖ�L@ '�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�4zL-b��kD��IZ3�L,OA�p@ϖ�L@ '�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0zL-c��kD��IZ3�L,OA�p@ϖ�L@ '�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0zL-c��kD��IZ3�L,OA�p@ϖ�L@ '�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0yL-c��kD��IZ3�L,OA�p@ϖ�L@ '�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0yL-c��kD��IZ3�L,OA�p@ϖ�L@ '�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0yL-c��kD��IZ3�L,OA�p@ϖ�L@ '�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0yL-d��jD��IZ3�L,OA�p@Ӗ�L@ +�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0yL-d��jD��JZ3�L,OA�p@Ӗ�L@ +�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0yL-d��jD��JZ3�L,OA�p@ӕ�L@ +�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0xL-d��iD��JZ3�L,OA�p@ӕ�L@ +�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0xL- e��iD��KZ3�L,OA�p@ӕ�L@ +�<;�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0xL- e�hD��KZ3�L,OA�p@ӕ�L@ +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0xL,�e�hD��KZ3�L,OA�p@ӕ�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0xL,�e�gD��KZ3�L,OA�p@ӕ�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0xL,�f�gD��KZ3�L,OA�p@ӕ�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0wL,�f�fD��KZ3�L,OA�p@ӕ�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0wL,�fܴfD��KZ3�L,OA�p@ӕ�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0wL,�fܰfD��KZ3�L,OA�p@ӕ�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0wL,�gܰeA��KZ3�L,OA�p@ו�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0wL,�gܰeA��KZ3�L,OA�p@ו�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0wL,�gܬdA��KZ3�L,OA�p@ה�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0wL,�g�dA��KZ3�L,OA�p@ה�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0vL,�g�cA��KZ3�L,OA�p@ה�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�XK�0vL,�h�cD��KZ3�L,OA�p@ה�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�X@�0vL,�h�cD� KZ3�L,OA�p@ה�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�X@�0vL,�h�cD� KZ3�L,OA�p@ה�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;l�X@�0vL,�h��bD� KZ3�L,OA�p@ה�L? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;\�X@�0vL,�i��bD� KZ3�L,OA�p@ה�H? +�<?�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;\�X@�0vL,�i��bD� KZ3�L,OA�p@ה�H? +�<?�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;\�X@�0uL,�i��bD� KZ3�L,OA�p@ה�H? +�<C�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;\�X@�0uL,�i��bD� KZ3�L,OA�p@ה�H? +�<C�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;\�X@�0uL,�i��bD� KZ3�L,OA�p@ה�H? +�<C�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;\�X@�0uL,�j��aD�KZ3�L,OA�p@ה�H? +�<C�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;\�X@�0uL,�j��aD�LZ3�L,OA�p@۔�H? +�<C�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;\�X@�0uL,�j��aD�LZ3�L,OA�p@ۓ�H? +�<C�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;\�X@�0uL,�j��`D�LZ3�L,OA�t@ۓ�H? +�<C�T0 k� ���#KP &�1D"3Q	E1 4#Q ��   � "�;\�X@�0uL,�j��`D�LZ3�L,OA�t@ۓ�H? +�<C�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;��X@�0uL,�j��`D�LZ3�L,OA�t@ۓ�H? +�<C�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;��X@�0tL,�k��_D�LZ3�L,OA�t@ۓ�H? +�<C�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;��X@�0tL,�k��_D�LZ3�L,OA�t@ۓ�H? +�<C�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;��X@�0tL,�k��_D�LZ3�L,OA�t@ۓ�H? +�<C�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;��X@�0tL�k��^D�LZ3�L,OA�t@ۓ�H? +�<C�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;��X@�0tL�k��^D�LZ3�L,OA�t@ۓ�H? +�<C�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;��X@�0tL�k��^A�LZ3�L,OA�t@ۓ�H? +�<C�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;��X@�0tL�l��]A�LZ3�L,OA�t@ۓ�H? +�<C�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;��X@�0tL�l��]A�LZ3�L,OA�t@ۓ�H? /�<C�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;��X@�0tL�l��]A�LZ3�L,OA�t@ۓ�H? /�<C�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;��X@�0tE\�l��]A�LZ3�L,OA�t@ۓ�H? /�<C�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;��X@�0sE\�l��\D�LZ3�L,OA�t@ۓ�H? /�<C�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sE\�l��\D�LZ3�L,OA�t@ۓ�H? /�<C�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sE\�l��\D�LZ3�L,OA�t@ۓ�H? /�<C�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sE\�m��\D�LZ3�L,OA�t@ۓ�H? /�<C�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sEL�m��[D�LZ3�L,OA�t@ۓ�H? /�<C�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sEL�m��[D�MZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sEL�m��[D�MZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sEL�m��[D�MZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sEL�m��ZD�MZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sEL�m��ZD�NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sE<�l��ZD�NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0sE<�l��ZD�NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��X@�0rE<�l��YD�NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�X@�0rE<�k��YD�NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�X@�0rE<�k��YD�NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�X@�0rE<�k��YL]NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�X@�0rE,�j��YL]NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�X@�0rE,�i��YL]NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�X@�0rE,�i��YL]NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�X@�0rE,�i��YL]NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�X@�0rE,�i��YL]NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�X@�0rB��i��YL]NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��   � "�;<�X@�0rB��i��YL]NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�X@�0rB��i��YL]NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�Y@�0rB��i��YL]NZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�Y@�0rB��i��XLmNZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;<�Y@�0rE,�i̜XLmNZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�Y@�0rE,�i̠XLmNZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�Y@�0qE,�i̠WLmOZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�Y@�0qE,�h̤WLmOZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�Y@�0qE,�h̤VLmOZ3�L,OA�t@ߒ�H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�Z@�0qK��g̤VLmOZ3�L,OA�t@��H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�Z@�0qK��g̨VLmOZ3�L,OA�t@��H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�Z@�0qK��g̨ULm OZ3�L,OA�t@��H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��   � "�;L�Z@�0qK��f̬ULm OZ3�L,OA�t@��H? /�<G�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;L�Z@�0qK��f̬ULm PZ3�L,OA�t@��H? /�<G�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;L�Z@�0qK��e̬TLm PZ3�L,OA�t@��H? /�<G�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;L�[@�0qK��eܰTLm$PZ3�L,OA�t@��H? /�<G�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;L�[@�0qK��eܰTLm$PZ3�L,OA�t@��H? /�<K�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;L�[@�0qK��dܰTLm$PZ3�L,OA�t@��H? /�"|K�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;L�[@�0qK��dܴTLm$PZ3�L,OA�t@��H? /�"|K�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;L�[@�0qK��dܴTLm(PZ3�L,OA�t@��H? /�"|K�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;L�[@�0qK��dܴTLm(QZ3�L,OA�t@��H? /�"|K�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;L�[@�0qK��dܴTLm(QZ3�L,OA�t@��H? /�"|K�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;L�\@�0qK��dܴSLm(QZ3�L,OA�t@��H? /�"|K�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;L�\@�0qK��d �SLm,QZ3�L,OA�t@��H? /�"|K�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;L�\@�0qK��d �SLm,QZ3�L,OA�t@��H? /�"|K�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;L�\@�0qK��c �SLm,QZ3�L,OA�t@��H? /�"|K�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;L�\@�0qK��c �SLm,QZ3�L,OA�t@��H? /�"|K�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;L�\@�0qK��c �SLm0QZ3�L,OA�t@��H? /�"|K�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;L�]@�0pK��c��SLm0QZ3�L,OA�t@��H? /�<K�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;L�]@�0pK��c��SLm0QZ3�L,OA�t@��H? /�<K�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;L�]@�0pK��c��SLm0QZ3�L,OA�t@��H? /�<K�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;M ]@�0pK��c��SLm4RZ3�L,OA�x@��H? /�<K�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;M ]@�0pK��c��SLm4RZ3�L,OA�x@��H? /�<K�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;M ]@�0pK��c��SLm4RZ3�L,OA�x@��H? /�<K�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;M ]@�0pK��c��SLm4RZ3�L,OA�x@��H? /�<K�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;M^@�0pK��c��SLm8RZ3�L,OA�x@��H? /�<K�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;M^@�0pK��d��SLm8RZ3�L,OA�x@��H? /�<K�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;M^@�0pK��d��SLm8RZ3�L,OA�x@��H? /�<K�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;M^@�0pK��d��SLm8RZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M^@�0pK��d��SLm8RZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M^@�0pK��d�SLm<RZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M^@�0pK��d�SLm<RZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M^@�0pK��d�SLm<RZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M_@�0pK��d�SLm<RZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M_@�0pK��d�SL]<SZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M_@�0pK��d l�SL]@SZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=_@�0pK��d l�SL]@SZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=_@�0pK��d l�SL]@SZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=_@�0pK��d l�SL]@SZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=_@�0pK��d l�SL]@SZ3�L,OA�x@��H? /�"�K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=_@�0pK��d ��SL]@SZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=_@�0pK��d ��SL]@SZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=`@�0pK��d ��SL]@SZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=`@�0pK��d ��SL]DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=`@�0pK��d ��SL]DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=`@�0pK��d ��SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=`@�0pK��d ��SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;=`@�0pK��d ��SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��d ��SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��d�SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��d�SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��d�SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��d�SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��d�SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��d�SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��d�SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��e�SA�DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��e�SA]DSZ3�L,OA�x@��H? /�<K�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0pK��e�SA]@SZ3�L,OA�x@��H? /�<O�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e�SA]@SZ3�L,OA�x@��H? /�<O�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e�SA]@SZ3�L,OA�x@��H? /�<O�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e\�SA]@SZ3�L,OA�x@��H? /�<O�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e\�SC�@SZ3�L,OA�x@��H? /�<O�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e\�SC�<SZ3�L,OA�x@��H? /�<O�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e\�SC�<SZ3�L,OA�x@��H? /�<O�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e\�SC�<SZ3�L,OA�x@��H? /�<O�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e�SC�<SZ3�L,OA�x@��H? /�<O�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e�SC�<SZ3�L,OA�x@��H? /�<O�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e�SC�<SZ3�L,OA�x@��H? /�<O�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e�SC�<RZ3�L,OA�x@��H? /�<O�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e�SC�8RZ3�L,OA�x@��H? /�<O�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e�SC�4RZ3�L,OA�x@��H? /�<O�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e�SC�4RZ3�L,OA�x@��H? /�<O�T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e�SC�4RZ3�L,OA�x@��H? /�<O�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e,�SC�0QZ3�L,OA�x@��H? /�<O�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;�`K�0oB��e,�SE�0QZ3�L,OA�x@��H? /�<O�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@l�e,�SE�,QZ3�L,OA�x@��H? /�<O�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@l�e,�SE�,QZ3�L,OA�x@��H? /�<O�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@l�e,�SE�,QZ3�L,OA�x@��H? /�<O�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@l�e,�SE�,QZ3�L,OA�x@��H? /�<O�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@l�e,�SE�(QZ3�L,OA�x@��H? /�<O�T0 k� ���#{P &�1D"3Q	E1 4#Q �    � "�;�`K�0o@��e,�SE�$PZ3�L,OA�x@��H? /�<O�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@��e,�SE�$PZ3�L,OA�x@��H? /�<O�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@��e�SE� PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@��e�SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@��e�SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@��e�SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@��e�SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��   � "�;�`K�0o@��e�SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@��e�SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@��e�SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@��e�SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0o@��e��SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��   � "�;�`K�0oA�e��SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SE�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SA�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SA�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SA�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SA�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SA�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SA�PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`K�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��   � "�;�`@�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SA]PZ3�L,OA�x@��H? /�<O�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SAPZ3�L,OA�x@��H? /�<O�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;�`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#KP &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e��SAPb��L,OA�x@��H? /�<O�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;=`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�eL�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�eL�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�eL�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�eL�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�eL�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�eL�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�eL�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�eL�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�eL�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�e<�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�e<�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�e<�SAPbs�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;M`@�0oA�e<�SAPZ3�L,OA�x@��H? /�<O�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��hE|�vB���M_�En��Z3��@^E�S�� 4|0q	M���T0 k� �P?�T?&�1D"3Q	E1 4#Q ��?    � (�8��hE|�uB���M_�En��Z3��@`E�S��5|4q	M���T0 k� �\=�`=&�1D"3Q	E1 4#Q ��    � (�8��jE��uB���M[�En��Z3��@`E�K~�6|8s	M���T0 k� �t8�x8&�1D"3Q	E1 4#Q ��    � (�9��jE��uB���MW�En��Z3�	|@aE�K~� 6|<s	M#�";�T0 k� ��6��6&�1D"3Q	E1 4#Q ��    � (�:��kE� tB���MT En� Z3�	|@aE�G�(6�@s'�"< T0 k� ��4��4&�1D"3Q	E1 4#Q ��    � (�;	�kE�tB���=TEn�Z3�	|@bE�G�07�Hs+�"< T0 k� ��1��1&�1D"3Q	E1 4#Q ��    � (�<	 lE�tB���=PEn�Z3�	|DcE�C��@7�Ps3�"<T0 k� ��-��-&�1D"3Q	E1 4#Q  ��    � (�=	mE�sB���=LE^�Z3�	|DcE�?��L7�Ps7�"T0 k� ��*��*&�1D"3Q	E1 4#Q  ��    � (�>	mE�sB���=LE^�Z3�	�DcE�?��T7�Ts;�"T0 k� ��(��(&�1D"3Q	E1 4#Q  ��    � (�?	nE�sB���-H	E^�Z3�	�DcE�;�~\7�Xt?�"T0 k� ��&��&&�1D"3Q	E1 4#Q  ��    � (�@	nE�$rB���-DE^xZ3�	�DdE�7�~l7�\tG�"T0 k� ��!��!&�1D"3Q	E1 4#Q  /�    � (�A	oE}$rB���-DE^pZ3�	�DdE�3�~t7�`tK�"T0 k� ��� &�1D"3Q	E1 4#Q  ��    � (�B	oE}(rB���-DC�l	Z3�	|DdE�3�~|7�`tO��T0 k� ��&�1D"3Q	E1 4#Q  ��    � (�D	pE},rB���-@C�d
Z3�	|DdE�/�~�7�dtW��T0 k� ��&�1D"3Q	E1 4#Q  ��    � (�F	qE}4qB��-<C�TZ3�	|DdE�+�~�6�ht-_��T0 k� �0�4&�1D"3Q	E1 4#Q  ��    � (�H	qE}8qB��-<C�PZ3�	|DdE�+�~�6�ht-c��T0 k� �<�@&�1D"3Q	E1 4#Q  ��    � (�J	rE}<qB��-8C�HZ3�	�DdE�'�~�6�ht-g�|T0 k� �H�L&�1D"3Q	E1 4#Q  �    � (�H	rEm<pB��-8C�@Z3�	�DdF'�~�5�ht-k�|T0 k� �0�4&�1D"3Q	E1 4#Q  ��    � (�G	 sEmDpB�/�-4C�0Z3�	�DdF#�~�4�lt-o�| 
T0 k� ��&�1D"3Q	E1 4#Q ��    � (�F	$sEmHpB�7�-4C�(Z3�	�DdF#�~�3�ls-s�| 	T0 k� ��	��	&�1D"3Q	E1 4#Q ��    � (�E	$tEmHpB�?�-0C�$Z3��DdF�~�3�ls-w�| T0 k� ����&�1D"3Q	E1 4#Q ��    � (�D	$tEmLpB�G�-0C�Z3��DdD����2�ps{�!� T0 k� ����&�1D"3Q	E1 4#Q ��    � (�C�(tEmLpB�O�-0C�Z3��DdD����1�pr�!� T0 k� ����&�1D"3Q	E1 4#Q ��    � (�B�,uEmPpB�c�-, C�Z3��DdD����/�pq��!� T0 k� �� �� &�1D"3Q	E1 4#Q ��    � (�A�0uEmPpB�k�-(!C� Z3��DdD����.�tq��!� T0 k� �w��{�&�1D"3Q	E1 4#Q ��    � '�@�0uEmPpB�s�-("C��Z3��DdD����-�tp��� T0 k� �_��c�&�1D"3Q	E1 4#Q ��   � &�?�4uEmTpI{� ($E��Z3��DdD����,�to��� T0 k� �K��O�&�1D"3Q	E1 4#Q ��    � %�>|8vEmTqI�� $&E��Z3��DdE���*�to��� T0 k� �#��'�&�1D"3Q	E1 4#Q ��    � $�=|8vD=TqI�� $'E��Z3��DdE���)�xn��� T0 k� ����&�1D"3Q	E1 4#Q ��   � #�<|8vD=TqI�� $(E��Z3��DdE�#��(�xm��� T0 k� ������&�1D"3Q	E1 4#Q ��    � "�;|<vD=TrI���$)E��Z3�L@dE�#��'�xm��� T0 k� ���#;P &�1D"3Q	E1 4#Q  �    � "�;|@vD=TsI,���$+E�Z3�L@cE|#��$$�|k��� T0 k� ���#;P &�1D"3Q	E1 4#Q�    � "�;�DuEmTtI,���$-E�Z3�L@cE|#��0!��i ���T0 k� ���#;P &�1D"3Q	E1 4#Q��    � "�;�HtEmPtI,���$/E�Z3�L@bE|#��8 ��i ��� T0 k� ���#KP &�1D"3Q	E1 4#Q��    � "�;�HtEmPuI,���$0E�Z3�L@bE|'��<��h ��� T0 k� ���#KP &�1D"3Q	E1 4#Q��    � "�;�LsEmPuE���$1E� Z3�L@bA�'��@��g ��� T0 k� ���#KP &�1D"3Q	E1 4#Q��    � "�;�LsEmLvE���$2E�!Z3�L@bA�'��H��f ����T0 k� ���#KP &�1D"3Q	E1 4#Q��    � "�;PrE]LvE���(4E��!Z3�L@bA�'��L��f ����T0 k� ���#KP &�1D"3Q	E1 4#Q��    � "�;PrE]HwE���(5E��"Z3�L@aA�'��T��e ����T0 k� ���#[P &�1D"3Q	E1 4#Q��   � "�;PrE]HwE���(6E��#Z3�L@aA�'��X��d ����T0 k� ���#[P &�1D"3Q	E1 4#Q��    � "�;TqE]DwE��,7E�x%Z3�L@`A�'��\��d ����T0 k� ���#[P &�1D"3Q	E1 4#Q��    � "�;XpE]@xE���,9E�p&Z3�L@`A�'��d��c ����T0 k� ���#[P &�1D"3Q	E1 4#Q��    � "�;\pEM@xE���,:E�l'Z3�L@`A�'��h��b ����T0 k� ���#[P &�1D"3Q	E1 4#Q��    � "�;\oEM<xE���0;D�d(Z3�L@`A�+��l��a ����T0 k� ���#kP &�1D"3Q	E1 4#Q��    � "�;`nEM8xE�'��0=D�`)Z3�L@_A�+��p��a ����T0 k� ���#kP &�1D"3Q	E1 4#Q��    � "�;`nEM4yE�3��0>D�X*Z3�L@_A�+��t��` ����T0 k� ���#kP &�1D"3Q	E1 4#Q��    � "�;dnEM4yE�;��4@D�P,Z3�L@_A�+��|
��_ ����T0 k� ���#kP &�1D"3Q	E1 4#Q��    � "�;dmE=0yE�C��4AD�L-Z3�L<^A�+��	��^ ����T0 k� ���#kP &�1D"3Q	E1 4#Q��    � "�;�hlE=,yE�K��4CD�D.Z3�L<^A�+����^ ����T0 k� ���#{P &�1D"3Q	E1 4#Q��    � "�;�llE=(xE�W��8ED�@0Z3�L<^A�+����] ����T0 k� ���#{P &�1D"3Q	E1 4#Q��    � "�;�pkE=(xL}_��8FD�<1Z3�L<]A�+����\ ����T0 k� ���#{P &�1D"3Q	E1 4#Q��    � "�;�tkE=$xL}g��8HD�42Z3�L<]A�+����[ ����T0 k� ���#{P &�1D"3Q	E1 4#Q��    � "�;�xjE- xL}o��<JD�04Z3�L<]A�+�� ��Z ����T0 k� ���#{P &�1D"3Q	E1 4#Q��    � "�;�|iE- wL}{��<KD�(5Z3�L<]A�/�����Z ����T0 k� ���#�P &�1D"3Q	E1 4#Q��    � "�;��iE-wL}���<MD�$7Z3�L<\A�/�����Y ��|�T0 k� ���#�P &�1D"3Q	E1 4#Q��    � "�;��hE-wL}���<OD� 8Z3�L<\A�/�����X ��|�T0 k� ���#�P &�1D"3Q	E1 4#Q��    � "�;��hE-vL}���<PD�:Z3�L<\A�/�O����X ��|�T0 k� ���#�P &�1D"3Q	E1 4#Q��    � "�;��hK�vL}���<RD�;Z3�L<\A�/�O����W ��|�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��hK�vL}���<TD�=Z3�L<[A�/�O����V ��|�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��gK�uL}���<VD�>Z3�L<[A�/�O����U ��|�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��gK�uL}���<WD�@Z3�L<[A�/�O����U ��|�T0 k� ���#�P &�1D"3Q	E1 4#Q .�   � "�;��fK�uL}���<YD� AZ3�L<[A�/�O����T ��|�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��fK�tL}���<[D��CZ3�L<ZA�/�O����S ��|�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��eK�tL}���<]D��EZ3�L<ZA�/�O����S ��|�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��eK�tL����<^D��FZ3�L<ZA�/�O����R ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��dK�tL����8`D��HZ3�L8ZA�3�O����Q ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��dK�sL����8bE��IZ3�L8YA�3�O����Q ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��dK�sL����8cE��IZ3�L8YA�3�O����P ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��cK� sL����4eE��JZ3�L8YA�3�O����P ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	�cK� sL����4gE��KZ3�L8YA�3�O����P ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	�cK��rL����0hE��LZ3�L8YA�3�O����O ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	�cK��rL����0hE��MZ3�L8XA�3�O����O ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	�cK��rL���0iE��NZ3�L8XA�3�O����O ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	�bK��rL���,jF�OZ3�L8XA�3�O����O ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	,�bK��rL���,kF�PZ3�L8XA�3�O����N ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	,�bK��rL���,lF�QZ3�L8XA�3�O����N ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	,�bK��rL���(mF�RZ3�L8WA�3�@���N ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	,�bK��rL�#��(nF�RZ3�L8WA�3�@���N ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	,�bK��rL�+��(oI��RZ3�L8WA�3�@���N ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	�bK��sL�/��$pI��SZ3�L8WA�7�@���M ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	�bK��sL�3��$qI��SZ3�L8WA�7�@���M ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	�cK��sL�;�� rI��SZ3�L8VA�7�@���M ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	�cK��sL�?�� rI��SZ3�L8VA�7�@���M ����T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;	�cK��sL�G��sI��SZ3�L8VA�7�@���L ����T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;	,�cK��tL�K��sJ�SZ3�L8VA�;�@���L ����T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;	,�cK��tL�O��tJ�SZ3�L8VA�;�@���L ����T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;	,�cK��tL�S��tJ�SZ3�L8VA�;�@#���L ����T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;	,�cK��tL�[��uJ�SZ3�L8UA�;�@#���L ����T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;	,�cK��tL�_��uJ�SZ3�L8UA�;�@'���L ����T0 k� ���#;P &�1D"3Q	E1 4#Q ��   � "�;	�cK��tL�c��uBL�SZ3�L8UA�?�@+���K ����T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;	�cK��uL�g��uBL�SZ3�L8UA�?�@/���K ����T0 k� ���#;P &�1D"3Q	E1 4#Q ��   � "�;	�cK��uL�o��vBL�SZ3�L8UA�?�@/���K ����T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;	�cK�uL�s��vBL�SZ3�L8UA�?�@3���K ����T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;	�cK�uL�w��vBL�SZ3�L8UA�C�@7���K ����T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�; �cK�uL�{��vA��SZ3�L4TA�C�@7���J ����T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�; �cK�uL���vA��SZ3�L4TA�C�@;���J ����T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�; �cK�vL����uA��SZ3�L4TA�C�@?���J ����T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�; �cK�vL����uA��SZ3�L4TA�C�@?���J ����T0 k� ���#[P &�1D"3Q	E1 4#Q ��    � "�; �cK�vL���� uA��SZ3�L4TA�G�@C��|J ����T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�; �cK�vL���� uA��SZ3�L4TA�G�@C��|J ����T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�; �cK�vL���� tA��SZ3�L4TA�G�@G��|I ��,l�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�; �cK�vL�����tA��SZ3�L4TA�G�@K��|I ��,l�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;L�cK�wL�����tA��SZ3�L4SA�G�@K��xI ��,l�T0 k� ���#kP &�1D"3Q	E1 4#Q ��    � "�;L�cK�wL�����sA��SZ3�L4SA�G�@O��xI ��,l�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;L�cK�wL�����sA��SZ3�L4SA�K�@O��xI ��,l�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;L�cK�wL~����sA��SZ3�L4SA�K�@S��xI �,l�T0 k� ���#{P &�1D"3Q	E1 4#Q ��   � "�;L�cK�wL~����sA��SZ3�L4SA�K�@W��tI �,|�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;|�cK�wL~����sA��SZ3�L4SA�K�@W��tH �,|�T0 k� ���#{P &�1D"3Q	E1 4#Q ��    � "�;|�cK�wL~����sA��SZ3�L4SA�K�@[��tH �,|�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�cK�xL~��\�sA��SZ3�L4SA�K�@[��tH �,|�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�cK�xL~��\�sA��SZ3�L4RA�O�@_��pH �,|�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�cKܐxE���\�sA��SZ3�L4RA�O�@c��pH �,|�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�cK܌xE���\�sA��SZ3�L4RA�O�@c��pH �,��T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�cK܌xE���\�sA��SZ3�L4RA�O�@g��lG �,��T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�cK܌xE���\�sA��SZ3�L4RA�O�@g��lG �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�cK܈xE���\�sA��SZ3�L4RA�O�@k��lG �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;|�c@��yE~��\�sA��SZ3�L4RA�S�@k��lG �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@��yE~��l�sA��SZ3�L4RA�S�@o��hG �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@��yE~��l�sA��SZ3�L4RA�S�@o��hG �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@��yE~��l�sA��SZ3�L4RA�S�@s��hG �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@��yE~��l�sA��SZ3�L4QA�S�@s��hG �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@��yD>��l�sA��SZ3�L4QA�S�@s��hG �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��   � "�;��c@�|yD>��l�sA��SZ3�L4QA�S�@w��dF �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�|yD>��l�sA��SZ3�L4QA�W�@w��dF �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�xyD>��l�sA��SZ3�L4QA�W�@{��dF �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�xzD>��l�sA\�SZ3�L4QA�W�@{��dF �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�xzD>��\�sA\�SZ3�L4QA�W�@��dF �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�tzD>��\�sA\�SZ3�L4QA�W�@��dF �,���T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�tzD>��\�sA\�SZ3�L4QA�W�@��dF �,��T0 k� ���#�P &�1D"3Q	E1 4#Q ��   � "�;��c@�tzD>��\�sA\�SZ3�L4QA�W�@���dF �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�pzD>��\�sA\�SZ3�L4QA�W�@���dF �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�pzD>��\�sA\�SZ3�L4QA�[�@���dE �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�lzD>��\�sA\�SZ3�L4QA�[�@���dE �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�lzDN��\�sA\�SZ3�L4QA�[�@���dE �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�lzDN��\�sA\�SZ3�L4QA�[�@���dE �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�lzDN����sA\�SZ3�L4PA�[�@���`E �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�h{DN����sA\�SZ3�L4PA�[�@���`E �<�T0 k� ���#�P &�1D"3Q	E1 4#Q ��    � "�;��c@�h{DN����sA�SZ3�L0PA�[�@���`E �<�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;��c@�h{DN����sA�SZ3�L0PA�[�@���`E �<�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;��c@�d{DN����sA�SZ3�L0PA�[�@���`E �<�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;��c@�d{DN����sA�SZ3�L0PA�_�@���`D �<�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;��c@�d{DN����sA�SZ3�L0PA�_�@���`D �<�T0 k� ���$P &�1D"3Q	E1 4#Q ��    � "�;��c@�`{DN����sA�SZ3�L0PA�_�@���`D �<�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;��c@�`{DN����sA�SZ3�L0PA�_�@���`D �<�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;��c@�`{D^����sA�SZ3�L0PA�_�@���\D �<�T0 k� ���#;P &�1D"3Q	E1 4#Q ��    � "�;                                                                                                                                                                            � � �  �  �  d A�  �K���� ' �     6 \��wp ]�

 � � `�o   � �	    ��D��     `�o�D��           	            	 Z�;          P�    ��    0	&
          o��      ��9     o���9                         Z�;         ��     ��   (	           e8�         �2��     e8��2��                      
	 Z�;         �     ��    0
           S#�   � �
    �/��     S#��/��                      *	 Z�;          ��    ��    H	$
          P�*    	    /�E��     P�*�E��           	            
	 Z�;          3P     ��    03            l� ��
	      C �;     l� �;                             ���k              �  ��    P		 5              Ow�  $ $      W�G1     Ow��G1                              ��        .�     ���   (
	          Ju      k��     Ju��                         � �         Y`     ���   
		          ���  $ I      :	K    ��� :	K                       	    �         .      ���   8	           ?q�          ����     ?q����                            �$         	 '0     ���   0
3         ��          ���۱    ����۱                           �$         
  0�     ���   H

         �� ��     ��L�    ���L�                             ���              }  ���    		 5 	                 ��      �                                                                           �                               ��        ���          ��                                                                 �                         ���E  ��        ���z    ���E��z         "                  x                j  �   �    �                             � <<       ���       ��   �    T�                                      . $       �                          ` o e S P  O �� ?����    ��         
    	      
  �   f �� .b�D       ��  }� �� }� � @c` �� `c� �D d� �d d� V� d� �  _� �D ` ���X � �d \� �D d� �d  d� �d b  Є b@ Ф b`���J ����X � J g@ J$ g` 
�\ W� 
�< W� 
� X  
� W� 
�\ X  �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  � }����� ����� � ބ �[� "� �`� #� a� �� �o� ��  p� �� 0q  �D q� S �j� T  k� TD l  Td l@���� � %� p� �� �e� �� @f� 
�< W� 
�� W� 
�| X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �����;�� "      �� �  "Df�
��� �  
   ���D"� �  " `   J jF  �  ffffffffff
 ff  �  ffffffffff  ff �  �  
�  e    ��     ���  �    o    ��     ��      ��    ��     � :          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �         �� � � ���        � � � ��        �        ��        �        ��        �   >�    ��������        ��                         ���    �                                     �                 ����             d��  �%�$�&��$   "�;��                 18/37 (48%) e o y      6:51                                                                       1  48     � �"% � �"	 � �"# �" �*%8 �*5P � "P c_	J�@ 
J�8c� c� c� �c� �c� � c� � �kk � ks � �C �C& � C%. � C& � C' �K; �K+ �B�8 � B�> �B�1 �B�9 � B�A �K/& � K7 �!c� �*""�A* #"�S$"�=%*�L s &*K~ � '*P~ � (*L~ � )*C~ � **K~; +*JfK ,*QV[ -*IV[  *Hv[ /*Lv[  *LV[ 1*Lv[  *LV[ 3*Lv[  *LV[  *LV[  *LV`  *LP]  *LP8 9*E`P :*ShX ;*LpX  *LP �  "F p#>*;3  *H                                                                                                                                                                                                                         G �   �        C 
     %d �     P P E _  ��                    ������������������������������������� ���������	�
���������                        �                                                                ��    �|� � 
������������ �!�"�#�$�k�l�'�(�)�*�+�m�n�o�/�0�1�2�p�q�r�6�7�1�2�N�s�O�;�<�1�2�=�a�?�2�@�A�B�C�t�E�B�F ��o ?   ����� �Q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     4       ��J     �]                              ������������������������������������������������������                                                                                                                                            ����  ��                                             �� ����� � �������  �� �������������������������� ������� �������������� �  ���� ������������������ �� ��� ������� ��� ��� ��� ���� ���� ���  ���������������������������  ������������������  ������� �������������������� ����������� ���                                   �     %    �� 
ĳJ      	�  	                           ������������������������������������������������������                                                                                                                                              ����  �  �                                           ������ � ������������� ����� ���������� �� �� ������������������ ������������������������������ ����� ������  �������� ������� ������� ������������� �������������� ����� ���� ��������������������  �� �������������� �����                                                                                                                                                                                                                                                                                                 	           
                   �              


           �   }�       ���������������������������������������������˾ܽ������˽��۾������������ܽ��ݼ�����������ܽ��ݼݼ�����������ܽ��ݼ�����������������ܿ��ݼ�����������ݽ��˼�޼�ݼ���˼�������������������������ݼ�����������������������������������������������������ܻ�ܻ����� : D 7                                  � ��� �G                                                                                                                                                                                                                                                                                         1p1Y"$  )n!�              l            k         W       m                                                                                                                                                                                                                                                                                                                                                                                                                � � �  � q��  � #��  � #��  � #��  � ��  �����&�����������h����������\����������h�����#                 u � :�� {       $   �   &  QW  �   y                    �                                                                                                                                                                                                                                                                                                                                      0 K K            (             !��                                                                                                                                                                                                                            Z   �� �~ �       �� e      �� ����� � �������  �� �������������������������� ������� �������������� �  ���� ������������������ �� ��� ������� ��� ��� ��� ���� ���� ���  ���������������������������  ������������������  ������� �������������������� ����������� ��������� � ������������� ����� ���������� �� �� ������������������ ������������������������������ ����� ������  �������� ������� ������� ������������� �������������� ����� ���� ��������������������  �� �������������� �����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     =   !   5   "� ��                       e     �   �����J���J'      ��     *   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ��  � ��     � ��   	 ��   p �� �� ��   ��   ��   ��     ��    �� �� �z ��   � ��    �� �� �z    P� �$  ��    ��   � �� �� �z   � �   �$ ^$      �    ��  � ��     ��  x x  0         �  0         �   ����2����  @ �J �            �     �     ��    � �J���2������}����     ��  ~�  }dQ   yL      ����������������������������������ܻ�ܻ�ܻ�ݻ��������������ݻ�������������������������������������������������������������������������������������ܻ�ܻ�ܻ��������������ܻ�ݻ�����������������������������������������������������������������������������������۽�������ݻ���ܻ��ܻ�ܻ�ܻ����������������������������������������ܻ�ݻ��ݼ�����������������ݽ��ͽ�������������ݼ����޻�����ܼ�ܻ�ݻ��ݽ�����������ܽ��ݼ�������������������ܻ�����������������ܼ�ܻ�ݻ������������������ݻ�����������������������������������������������������������ܻ����������������������������������ܼ���˽�������ݻ�������������������������������ݼ���ۼ�����������������������������������������ۻ�������������������������ۼ������������ܽ��ݼ�����ݼ���۽���������������������������������������ܽ��ݼ����������ܼ�ܻ�ܻ�ݻ�������������������������������������������������������������������������������������������ܻ�����������ܻ�����������������������ݻ�����������������������������������������������������ܻ�ܻ�ܻ��������������ܻ�ݻ����������������������������������������ܽ��ݼ�����������ܻ�������ͻ�ܽ��ݼ���˾�ܽ��������������������������������������ܽ˾ݼ���������������������������������������ݽ��ݽ��������������������������������������������������������������������������������������������������ݼ���۽�������ݻ���ܼ�������������������������������ݽ�������ݻ�ݻ���������������������������������������������������������������������ܻ�ܻ�ܻ�ݻ���������������������������������������ܼ�����������ݻ��ݽ���˼�����������ܽ�ݻ���������ܽ��ݽ��ܽ�����ܼ���˼���������������������������������������������������ܽ��ݼ��ܼ��������˼�˼�˼�����������������������������������������������������������������������������������ܼ���۽�����������������������������������ݻ���ܼ���۽�������ݻ����������������������ݻ��������������ܻ�ܻ�ܻ�ݻ��������������ݻ������������������������������������������˾ܽ������˽��۾������������ܽ��ݼ�����������ܽ��ݼݼ�����������ܽ��ݼ�����������������ܿ��ݼ�����������ݽ��˼�޼�ݼ���˼�������������������������ݼ�����������������������������������������������������ܻ�ܻ��������������������������������������"�"���-��-��-"-�-�������������-���������������-��������������!���!�!!"�!�����"����������������!!-!!-!!��---������!�-�!-!!"�!��!���-����������������"�--��-����-��-��-���-�����-���-����-�"-������-���������������������-���-����������"""�"���""-���--�!-�"��-�"�--���-����-���-��-��������������������������!""��-���-���-�������-���-��"�-��"���-�������������"�-"��-��"����������-���"-�-���-������������������������������������������������""-������������������������������������������������-��-�"��-�"��-��������"!-�-�-�-��"�""-���������������������"-��"!�-���"�"-"-��"""��"!����"��!���"�""-����-�-"-�""����"""""��"!������"�""-��""-���"!-��"�""-"!�-"��-�"��-����""���"!-��""!-��"�""-��"!-���"!���"�""-�������������������������������������������"�������������������"""��������������������������""���""�����������"���-�-�"���-������-�����!���-�!!-�-�""�����"����������-"!-��-�"��!���"�!��"�""-��"!-�"-��-��-��"�""-��!��������"�""-�"������"����"""�"������"�������"-���"!-�"--�-��"�""-��-�-�"!-�-��-�"����-����������������"-����"��-��-�---�-�""���"�-�"�������"�"���-�������������"""��!!-!-�-��-�"����!�---��-�"��!���"�"-������"-���"!-�-�!�-���""-��!���"�!����"�"��"!-�"���"!���"�""-!!����������������"-�������������"��"-��-��-�"�-�-�-����"���-�-�!�"��-�"��-��"�-��"�-��-�"��-����"��-�������"-"!��"��-�"��-�"""�����-��-��""�-���-���-������������!"��-��"���-���������������������������"""�����������"��-"-��"""���-���"�-----�""�����������"�-�--��-�""������-�-"-----��"""����������"!�-""-���""-���"�������-�������"-����������""--�-�"-�-���-���"�------�-�-�����-�����-��-��-����""�������-�����-��-��-�-�-���-��-�!-"�!�-��-�-����-��-��-��-��-����""����������!!!!�-"�����������!�������"�"����������"�----�-�""����������"�---""�-�����������""--�-�"-��-�����������"�"��-����""�����������""-���"�-�""�����������"-�-��-������"-����������------��"""����������----�-�"���-����������!!!�!��"�-�����������"�-��"��-�"����������----�-�"-�-����������!-�"��-���""-���������-��-�������-�����������������-����������-��-�����wwwwwwww33333333333333333333wwwvwwwv33363336333633363336FdffFdffAC333C333C333C333C333��������33333333333333333333�f�f�fFf�33�333�333�333�333�3�fff�fff33333333333333333333ffffffff33333333333333333333333d333d333d333d333d3333����wwww333333333333333333333333����wwww333633363336333633363333����wwwwC333C333C333C333C3333333����wwww33�333�333�333�333�33333����wwww�����<��5UUU5UUSU553SS2#33"532 5�����<��5UUU5UUUU555SSSS33333��������UUUUUUUU5555SSSS3333��������UUU�UU_�55=�SS]�33;������l���eUUUUUUSU552SS2#S3"3S2 0�����<��5UUU5UUSU552SS2#33"332 0����ȩ��S�UUU��US:�U59��38��009������<��UUUUUUUU5555SSSS33333������ÓUUX�UUS�SSX�553�338�003�����3���UUUU5UUUU555SSSS33333�����̚�Ue�5UX�U5Y�5X��S9��3����������UUUUUUUSU5523S2#"302 0�����<��5UUU5UUSU552SS2#33"302 0�����<��5UUV5UUUU555SSSU33353��������UUUUUUUUU5553SSS33330����l���eUUSUUU3SSS%U3"5S2#3S" "#  %                     200            "          "                         0;�  ��  �� ��  ۰  ۰  ��  ��                          #                         P"R                         "#                       "#  "                    0"                                                    �  9                     �#�� ��� ��� ��  �       02(�" �  � ��0(�������� �����   �                    "                         205            "         R 20R                                                                                    ��  ��  �� �� �  �  �  �   �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��  �S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                                                  U  T   T   T     T UDUDDUDDDDDDDDDDDDDDDP   E�  DU� DDU�DDDUDDDDDDDDDDDD                UP  E�  E   E                                           ���U�UTD�DDDDDDTDD TDD   �   U_ DEU�DDDUDDDDD��DZT�DDDDDDDDDDDDTDDDDDDDDUTU�����DDDDDDDDDDDEDDDEDDDDTUTU�Ԫ���Z_   P   � �U�UTDUDDDDUTD�DT��D        U_��DEU_DDD_DDDPDDE�DDE  �DD DD DD �DD �UD  �U       DZTDEDDDDE�DDE�DDE�TDDT�DE�TE���DDTU�ZD���������DDTDD��ZT�T���ZTDDE��D��T�T��DUTTT��Z��TQTDDUTD�DDDTDDD�DDDDDDE�DD_TDE�DD_ DDP DDP DD_ DU_ U�  �                                       TE�DDD�UUU                    ���DDDUUUTD  D  D  D  D  U��D�TDDDDEUUDP  DP  DP  DP  UP  TDE�DDDPUUU_                                                    wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwtwwwCwwt1wwCwt1wC�t1��C1����������""""���������������!���""!����,���ww��7����������������wwwwwwwwwwwwwwwwwwww7wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwws��w1wt1�wC�t1��s��s��s������"$��Gw�!������������L���q��"r��������!�����!ww�r�w�ww!�wwrwwwwwwqwwwrwwww�7ww�ww�ww��7w��w���G��'!wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����   �   �   �   ����                                     	�  		  	 � 	 	 	   	   	   	   	  ��                  ��   	   	   	   	   	   	 	 	 � 		  	�                 �   	    �   	    �   	    �   	   	   �  	   �  	   �  	   �                      �   �   
                                       
   �  
   �  
   
   
    �   
�            ����        �   
    �   
    �  
   �  
   �      
   �  
   �  
   �  
   �                   ����   
   
   
   
   
   
   
   
   
   
�  

  
 � 
 
 
  �
  

   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         "!  "" "  """ ""   "! " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  "! ""! " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """ "!    " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                          �  �� �� wȠb���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 " "" "  �   �   �           �   �   �           �  "�  "                   �     �                                                                                                                                                                                                  �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��r`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   �". ". ����                /���"/�  ��                    �                                                                            �               �     "   "               !��� �                                                                                                                                                                                                       �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp��& ��vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �" �"" �"   �                    .   .   �    �   �".  .                            �   �    �   �       �   �   �                .      ���.�                         ��   �  ��  �  �  �         � ".��".��/����  �                                                                                                                                                                              " �"  �      �    "" ""  "!� !������������ ����  ��  "  ""  "!  "���                     
         �  � "��""- �"- "   � "� ""� ""$ "$  C  3  �  �  �   �   +w{� &'� vv� �w� ��� ɪ������˹��̻����̰݊� �ɨ �˅@̻�@�D�@4U�@4U� 4U� 4U� 3UXP�EX��U����  ��                    �  ��� ݼ� �    �    �   �                     �         "   "   �                                     �  ��� ݼ� w{� &'� vw�                    �   ���                            �   "                                                                                                                 �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp��& ��vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �" �"" �"   �                    .   .   �                   �   ��  �ڛ�}ک�"   "   "  �� ��                   �".��".���                                  "  .���"    �     �                                                                                                                                                                                           �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ����))������؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� ����"  �". �.  �                                        �� ��                  �          �         �   �  �  �   �               �   �                  �   � �                   �         �  "� "  �  ��                                                                                                                                            �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   �   " � ��      �    �       �   ��  �   �    �  ��   �"" �"  �                        .   .   �                              �".��".���                   �  �  �  �               ���                                                                                                                                                                                            �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���        T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ��"� �"� ����                                                                                                                                                                                                                                        b}z�gg��j�� 
�� 	�� �� �� 
�� �� ��̻�"+��" 4"  4   D   H   H   �  +  ""    ��       ��  �٠ �ڛ ̸� ̻� �̽ �̀ �ɀ ��0 ��C 4�T H�T H�D �T@ �T  �C  �0  ɚ  ��� ��� �" �"  �"�                 �� �� �� {�             �   �  " � "�� � �  ��                                        �   �   �   "   "   "  !�    ��                              �                        ��"� �"� ����                            �   ���                                                                                                                                                                                                     �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���                        �   �   �   "   "   "  !�    ��              "   "   "  �� ��                   �".��".���                          .  ". ""  "    � ���                                                        ���                          ����                  �   �� �       �  �  "�  "   "                                             �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �               �   �       �       Ț  ��  ��" �"��"/��"���  �             "   "      �  �                         �  ���               �".��".  ���    �       �  �  �  �               ���                                                                                                                                                                                                                     �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ���������""��""��""�����        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  "   "                                                                              2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ DD D@  �D�JJN�I��I��I��I��JJD�N�                    �   �        �� ���ɑ��� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ����������������""��#3��#w��#w������������""""3333wwwwwwww�������������""9�34y�w4y�w4y���#w��#w��#w��#w��#w��#w��#w��#wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4y�w4y�w4y�w4y�w4y�w4y�w4y�w4y���#w��#w��#3��$D��7w������������wwwwwwww3333DDDDwwww������������w4y�w4y�34y�DDy�wwy�������������                                ""     "                                      !  ! !!"!   "             !! !! !!         ! ! !!"! !                "                              "                                     """" ""     !  "   "                                      !""                   "   "                " "    "             "                                                 ""                                                  "   "         "!    " ""                "  "!  "" "  """ "!  " ! " ""      " ""   """"" "!   " ""  ""   "! " "" "! "   "      ""  "! ""! " ""  "!  "! " ""                                         "              """                         ""  ""          "      "            !  !!  ""    "         "!   " !"!"""  "!  "       " ""  !""" "  "  """"  "     "   "!  "   " ""    "!    "               "    "            "" " "   " "           """ !! !    " !     " !""     "   "!  !  ""  !"!" " "!  "  "! " "" !!          "  " "    "       "    !"  "  "   "   "     "       " "!  "   "  """        ""                 !"   "                              """          "  "  """       "      ""          "       ""        "      """         "!  ""   ""   "           "          ""    "         "                            ""                              ! " !                        ""          !!!! "         ! " "         "       ""          "    ""            ""    "             " "      ""          ""   "  ""          "           "                  """                "            !!!! "           "   "  "                "            !  "    ""                                               wwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD������������������=�J�V�Y�L����������������������������������������������������������������������������������������������������������������������������=�O�V�[�Z�����������!��������������������������������������������������������������������������������������������������������������=�O�V�V�[�P�U�N��:�J�[������ ����������������������������������������������������������������������������������������������������������������-�Y�L�H�R�H�^�H�`�Z��������� ���������������������������������������������������������������������������������������������������������������U�L��>�P�T�L�Y�Z���������!������������������������������������������������������������������������������������������������������������:�L�U�H�S�[�`��=�O�V�[�Z��������������������������������������������������������������������������������������������������������������!�������1�H�J�L�V�M�M�Z��A�V�U���������������������������������������������������������������������������������������������������������������������-�V�K�`��.�O�L�J�R�Z���������%��������������������������������������������������������������������������������������������������������������:�L�U�H�S�[�P�L�Z���������������������������������������������������������������������������������������������������������������"�&�!������,�[�[�H�J�R��D�V�U�L������� �&�� �������������������������������������������������������������������������������������������������$���#��b� �$��c����:�H�Z�Z�P�U�N������ ��!���b� �"��c����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������LDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDD    "% � �"	 � �"# �" �*%8 �*5P � "P c_	J�@ 
J�8c� c� c� �c� �c� � c� � �kk � ks � �C �C& � C%. � C& � C' �K; �K+ �B�8 � B�> �B�1 �B�9 � B�A �K/& � K7 �!c� �*""�A* #"�S$"�=%*�L s &*K~ � '*P~ � (*L~ � )*C~ � **K~; +*JfK ,*QV[ -*IV[  *Hv[ /*Lv[  *LV[ 1*Lv[  *LV[ 3*Lv[  *LV[  *LV[  *LV`  *LP]  *LP8 9*E`P :*ShX ;*LpX  *LPqqDqwqwwDwtwwww3333DDDDAqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD���������������������������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD������� �!�"��� ����n�o�}�~�d�e�w�x����������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ���#�$�k�l�'�(�)��� ����������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ���*�+�m�n�o�/�0��� �� ��8�H�U�Z�V�U��b��c�������""""UUUUUQQADAQQ""""UUUUUUUAUQEE���1�2�p�q�r�6�7��� ���,�Z�Z�P�Z�[��I�`�&��������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD���1�2�N�s�O�;�<��� ��"��<�L�P�J�O�L�S��b��c������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD���1�2�=�a�?�2�@��� ��$��=�H�]�H�Y�K��b��c�������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD���A�B�C�t�E�B�F�����������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD��������������������������������""""-���-���-���-���-���-���""""�����������������������������������������������������""""�������A��A�A""""�������A��A�A��������������������������������""""������MDDMA��M""""��������������������������������������������������������������������������������3333DDDD�DD�H�H����3333DDDD���������������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��������������������������������������������������������3333DDDD���4���4���4���4���4���43334DDDD��������������������������������""""������A�D��I��""""�������D����������������������������������""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��>�%�$�&��$���������������� �8�>�7������A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �>��<�����""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,�����������DDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II����������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	���������������������������������������� ����������������������������������	�	�	�*����������������������������� ���	�
��������������������������������������6�	�	�7�������������������������+��,�-� ����������������������������������	�	�������������������������8�9�:�;� ��n�o�d�e�y�z�l�m�x�x���������d�e�����r���������r�h�i����������	�������������������������
���� ������������������x�x�ŤƤǤȤ����ǤȤ��ŤƤǤȤ������ŤƤ��!�"�#�$�������������������������������������������������������������0�1�2�%��4�U�Z�[�H�U�[��<�L�W�S�H�`����������	�%����� ���������-�.�/�0�1�2�%����3�4�5������������?�	�@����0�K�P�[��7�P�U�L�Z��������������	�
����������;�<�=�>�?�	�@����������������������������	�A�������������������������         	 	 
     	 	 	 	       	    	     	 	 	 	 	 ������������������������      	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *������������������������        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7������������������������ +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	������������������������ 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	������������������������ 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                