GST@�                                                           @^�                                                        �   ��             	      ��������	 J�����������X���z���        �h     #    z���                                d8<n    �  ?     B����  �
fD�
�L���"����D"� j   " B   J  jF�"    "�j* ,  �����
�"     �j@ �    ��
  )�                                                                              ����������������������������������      ��    bb QQb  114 44c c   c      		 

       	   
       ��G �   ( (                 nhp ))1         888�����������������������������������������������������������������������������������������������������������������������������?=  00  54  81                        
     
                ��  4�  �  ��                  Yn  	          : �����������������������������������������������������������������������������                                �]  ]   �  ��   @  #   �   �                                                                                'w w  )n)h1p  Y	n    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E ) �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������     ��P��D���� r�M|,SQ�E�S�  ���4=�T0 k� �D$�H$!Q8D"%d1O   ��   � 0 � ��P��D���� r�M|,SQ�E�O�  ���4<�T0 k� �D#�H#!Q8D"%d1O   ��   � 0 � ��P��D���� r�M|,SQ�E�K�  ���0;�T0 k� �@#�D#!Q8D"%d1O    ��  � 0 � ��P��D���� r�M|,SQ�E�G�  ���0:�T0 k� �@"�D"!Q8D"%d1O    ��   � 0 � ��P��D���� r�M|,SQ�D2C�  ���,9�T0 k� �<!�@!!Q8D"%d1O    ��   � 0 ��P��D���� r�M|,SQ�D2?�  � �,8�T0 k� �< �@ !Q8D"%d1O    /�   � 0 ��Q�
D����r�N|,Sa�D27�  ��(7�T0 k� �8�<!Q8D"%d1O    ��   � 0 ��Q�D����r�N|,Sa�D23�  �s(6�T0 k� �8�<!Q8D"%d1O    ��   � 0 ��Q�D����r�N|,Sa�D2/�  �s$5�T0 k� �4�8!Q8D"%d1O    ��   � 0 ��Q�D����r�N|,Sb D2'�  �s$4�T0 k� �4�8!Q8D"%d1O    ��   � 0 ��Q�D����r�N|,Sb D2#�  �s$3�T0 k� �0�4!Q8D"%d1O    ��   � 0 �Q�Q�D����r�N|,SbD2�  �s 2�T0 k� �0�4!Q8D"%d1O    ��   � 0 �Q�Q�D{���r�N|,SrD2�  �c 1�T0 k� � �$!Q8D"%d1O    ��   � 0 �Q�Q�Dw���r�N|,SrDB�  �c/�T0 k� ��!Q8D"%d1O    ��   � 0 �Q�P��Do���r�N|,SrDB�  �c.�T0 k� ��!Q8D"%d1O    ��   � 0 ���P��C�_���r�N|,SrDB�  �c,�T0 k� ��� !Q8D"%d1O    ��   � 0 ��{�P��C�W���r�N|,SrDB�  �c+�T0 k� ����!Q8D"%d1O    ��   � 0 ��{�P��C�O���r�N|,SrDA�   �c)�T0 k� ����!Q8D"%d1O    ��   � 0 ��{�E��C�G���r�N|,SrDA�   �c(3�T0 k� ����!Q8D"%d1O    ��   � 0 ��w�E��C�?���r�N|,SrDA�   �c'3�T0 k� ����!Q8D"%d1O    ��   � 0 ��w�E��C�7���r�N|,Sr DA�  �c%3�T0 k� ����!Q8D"%d1O    ��   � 0 ��s�E��C�/���r�N|,Sr$DA�  �c%3�T0 k� ����!Q8D"%d1O    �   � 0 ��o�E��C����r�O|,Sr(DA�  �S$3�T0 k� ����!Q8D"%d1O    ��   � 0 ��k�E��C����r�O|,Sr,DQ�  �S$3�T0 k� ����!Q8D"%d1O    ��   � 0 ��g�A��C����r�O|,Sr,DQ�  �S$3�
T0 k� �� �� !Q8D"%d1O    ��  � 0 ��g�A��C����r�O|,Sr0DQ�  �S$3�
T0 k� ��#��#!Q8D"%d1O    ��   � 0 ��c�A��C���� r�O|,Sr0DQ�  �S $3�
T0 k� ��%��%!Q8D"%d1O    �   � 0 ��[�A��C���rr�O|,Sr8DQ�  �b�$3�	T0 k� "�&��&!Q8D"%d1O   ��   � 0 ��W�A��C���rr�O|,Sr8DQ�  �b�$3�	T0 k� "�'��'!Q8D"%d1O   ��   � 0 ��S�A��C���rr�O|,Sr<DQ�  Cb�$3�	T0 k� "�'��'!Q8D"%d1O   ��   � 0 ��O�A��C���rr�O|,Sr<E�  Cb�$3�	T0 k� "�(��(!Q8D"%d1O   ��   � 0 ��K�A��C���rr�O|,Sr@E�	  Cb�$3�	T0 k� "�)��)!Q8D"%d1O   ��   � 0 ��G�A��C���rr�O|,SrDE�
  C��$�
T0 k� "�)��)!Q8D"%d1O   ��   � 0 �C�A��C��br�O|,SrDE�
  C��$�
T0 k� ��*��*!Q8D"%d1O   ��   � 0 �;�Eb�C��br�O|,SrHE�  3��$�
T0 k� ��*��*!Q8D"%d1O   ��   � 0 �7�Eb�C��br�O|,SrLE�  3��%�
T0 k� ��+��+!Q8D"%d1O   ��   � 0 �3�Eb�Eҧ�br�O|,SrPE�|  3��%�
T0 k� ��,��,!Q8D"%d1O   ��   � 0 �/�Eb�Eҟ�br�O|,SrPE�x  3��%�
T0 k� ��,��,!Q8D"%d1O   ��   � 0 �'�Eb�Eҗ�"r�O|,SrTE�p  3��%�
T0 k� 2�-��-!Q8D"%d1O   ��   � 0 �#�ER�Eҏ�" r�O|,SrTE�l  ��%�
T0 k� 2�.��.!Q8D"%d1O   ��   � 0 ��ER�E҇�!�r�O|,SrXE�d  ��%�
T0 k� 2�.��.!Q8D"%d1O   ��   � 0 ��ER�E��!�r�O|,Sr\E�\  ��%�
T0 k� 2�/��/!Q8D"%d1O   ��   � 0 ��ER�E�w�!�r�O|,Sr\E�X  ��%�
T0 k� 2�0��0!Q8D"%d1O   ��   � 0 ��ER�E�o�!�	r�O|,Sr`E�P  ��%�
T0 k� ��0��0!Q8D"%d1O   ��   � 0 ���ER�E�_�!�r�P|,SrdE�D  
���%�
T0 k� ��2��2!Q8D"%d1O   ��  � 0 ���ER�D2W�!�r�P|,SrhE�@  
��%�
T0 k� ��2��2!Q8D"%d1O   ��   � 0 ��ER�D2O�!�r�P|,SrhE�8  
��%�
T0 k� ��3��3!Q8D"%d1O   ��  � 0 ��ER�D2G�!�r�P|,SrlE�4  
�R�%�
T0 k� "�4��4!Q8D"%d1O   ��   � 0 ��EB�D2?�!�r�P|,SrlE�0  
� R�%�
T0 k� "�4��4!Q8D"%d1O   ��   � 0 �߽EB�D27�!� r�P|,Srp
E�(  
� R�%�
T0 k� "�5��5!Q8D"%d1O   ��   � 0 �׽EB�D2/�!��r�P|,Srp
F$  
� R�%�
T0 k� "�6��6!Q8D"%d1O   ��   � 0 �ϽEB�D2'�!��r�P|,Srt
F    
�$R�%�
T0 k� "�6��6!Q8D"%d1O   ��   � 0 �˽EB�D2�!��r�P|,Srt	F!  
�$R�%�
T0 k� �7��7!Q8D"%d1O   ��   � 0 �ýC��D2�!��r�P|,Srt	F#  
�(R�&�
T0 k� �8��8!Q8D"%d1O   ��   � 0 �໽C��D2�!��r�P|,SrtF$  
�(R�&�
T0 k� �8��8!Q8D"%d1O   ��   � 0 �೽C��D2�!��r�P|,SrtF&  
�,R|&�
T0 k� �9��9!Q8D"%d1O   ��   � 0 �૽C��D1��!��r�P|,SrtF'  
�0Bx&�
T0 k� �:��:!Q8D"%d1O   ��  � 0 ����EҔDA��!��r�P|,SrtF *  
�4Bh&�
T0 k� B�;��;!Q8D"%d1O   ��   � 0 ����EҔDA��	�����P|,SrtF �,  
�8B`&�
T0 k� B�<��<!Q8D"%d1O   ��   � 0 ����EҌDA��	�����P|,SrtF �-  
�8BX&�
T0 k� B�<��<!Q8D"%d1O   ��   � 0 ����EҀDA��	�����P|,SrtF �/  
�<�T&�
T0 k� B�=��=!Q8D"%d1O   ��   � 0 ��{�E�xDA��	�����P|,SrtE��0  
�@�L&�
T0 k� B�>��>!Q8D"%d1O   ��   � 0 ��s�NRpDA��	�����P|,SrtE��1  
�D�D&�
T0 k� �>��>!Q8D"%d1O   ��   � 0 ��k�NRhDA��	�����P|,SrtE��3  
�H�<'�
T0 k� �?��?!Q8D"%d1O   ��   � 0 ��g�NR`DA��	�����P|,SrtE��4  
�L�4'�
T0 k� �@��@!Q8D"%d1O   ��   � 0 ��_�NRTDA��	�����P|,SrtE��6  
�PB,'�
T0 k� �@��@!Q8D"%d1O    ��   � 0 �W�NRLDA��	�����P|,Srt E��7  
�PB$'�
T0 k� �A��A!Q8D"%d1O    ��   � 0 ~�O�NRDDQ��	���"�P|,Srw�E��8  
�TB'�
T0 k� "�B��B!Q8D"%d1O    -�   � 0 }�G�NR<DQ��	���"�P|,Srw�E��:  
�XB(�
T0 k� "�B��B!Q8D"%d1O    ��   � 0 |�7�NR,DQ��a��"�P|,Srw�B��<  
�\B(�
T0 k� "|C��C!Q8D"%d1O    ��   � 0 {�/�NR$DQ��a��"�P|,Srw�B��=  
�\A�)�
T0 k� "|D��D!Q8D"%d1O    ��   � 0 z�'�NRDQ�a��"�P|,Srw�B��?  
�`A�)�
T0 k� �xE�|E!Q8D"%d1O   ��   � 0 y��NRDQw�a��"�Q|,Srw�B��@  
�`A�*�
T0 k� �xE�|E!Q8D"%d1O   ��   � 0 x��NRDQo�a��"�Q|,Srw�B��A  
�`A�*�
T0 k� �tF�xF!Q8D"%d1O   ��   � 0 w��NRDQg�Q��"�Q|,Srw�E��B  
�dA�+�
T0 k� �tG�xG!Q8D"%d1O   ��   � 0 w �NR DQ_�Q�� ��Q|,Srw�E��C  
�dA�+�
T0 k� �pG�tG!Q8D"%d1O   ��   � 0 v��NQ�DQW�Q�� ��Q|,Srw�E��E  
�dA�,�
T0 k� 2pH�tH!Q8D"%d1O   ��   � 0 v��NQ�DaO�Q�� ��Q|,Srw�E��F  
�h1�,�
T0 k� 2lI�pI!Q8D"%d1O   ��   � 0 u�NQ�DaG�Q�� ��Q|,Srw�E��G  
�h1�-�
T0 k� 2lI�pI!Q8D"%d1O   ��   � 0 u�NQ�DaC��� ��Q|,Srw�E��H  
�h1�.�
T0 k� 2hJ�lJ!Q8D"%d1O   ��   � 0 to߽NQ�Da;��� ��R|,Srw�E��I  
�h1�/�
T0 k� 2hK�lK!Q8D"%d1O   ��   � 0 to۽NQ�Da3���R|,Srw�E��J  
�h1�/�
T0 k� �dK�hK!Q8D"%d1O   ��   � 0 soӽNQ�Da+���R|,Srw�E��K  
�h1�0�
T0 k� �dL�hL!Q8D"%d1O   ��   � 0 soϾNQ�Da#���S|,Srw�E��L  
�h1�1�
T0 k� �`M�dM!Q8D"%d1O    ��   � 0 roǾE��Da���S|,Srw�E��M  
�h1�2�
T0 k� �`M�dM!Q8D"%d1O    ��   � 0 roþEѼDa���T!�,Srw�E��M  
�h1�3�T0 k� �\N�`N!Q8D"%d1O    ��   � 0 q��EѴDa���T!�,Srw�E��N  
�h1|4�T0 k� "XO�\O!Q8D"%d1O    ��   � 0 p��EѰDa���ҔU!�,Srw�E��O  
�h!x5�T0 k� "XO�\O!Q8D"%d1O    ��  � 0 p��EѨD0����ҐU!�,Srw�E��O  
�h!p6�T0 k� "\P�`P!Q8D"%d1O    /�D   � 0 p��I��D0����ҌV!�,Srw�E��P  
�h!d9�T0 k� "\Q�`Q!Q8D"%d1O    ��D   � 0 p��I��D0����ҌW!�,Srw�E��Q  
�h!\:�T0 k� �`R�dR!Q8D"%d1O    ��D   � 0 q��I��D0����B�W!�,Srw�E��Q  
�h!X;�T0 k� �hU�lU!Q8D"%d1O    �D   � 0 u��I��E���Q{�B�X!�,Srw�C@�R  
�h�P<�T0 k� �pX�tX!Q8D"%d1O   ��O  � 0 x���I��E���Qw�B�X!�,Srw�CA R  
�h�L=�T0 k� �t[�x[!Q8D"%d1O   ��O   � 1 {���I�|E���Qo�B�Y!�,Srw�CA R  h�H?�T0 k� �|^��^!Q8D"%d1O   ��O   � 2 ~���I�xE���Qk�B�Y|,Srw�CAR  h�D@�T0 k� ��a��a!Q8D"%d1O   ��O   � 3 ����I�pE��Qg�b�Z|,Srw�CAR  h�@A�T0 k� ��d��d!Q8D"%d1O   ��O   � 4 ���I�lE��Q_�b|Z|,Srw�CAR  h!<C�T0 k� ��g��g!Q8D"%d1O   ��O   � 5 �s�I�dE��QW�bx[|,Srw�CAR  Ch!4E�T0 k� ��m��m!Q8D"%d1O   ��O   � 6 �o�E�`E��QO�bt\|,Srw�CAR  Ch!4E�T0 k� ��p��p!Q8D"%d1O   ��O   � 7 �k�E�XE���QK�Rt\|,Srw�CAS  Ch!4F�T0 k� ��s��s!Q8D"%d1O   ��O   � 8 �g�E�TE��AC�Rt]|,Srw�CAS  Ch14F�T0 k� ��v��v!Q8D"%d1O   ��O   � 9 �c�E�PE���A?�Rp]|,Srw�CQT  Ch14G�T0 k� ��y��y!Q8D"%d1O   ��O   � : �c�E�HE�� A7�Rp^|,Srw�CQT  Ch14G�T0 k� ��|��|!Q8D"%d1O   ��O   � ; �_�E�DE��A3�Rl^|,Srw�CQT  Ch14G�T0 k� ����!Q8D"%d1O   ��O   � < ��[�E�<E�xA+�Bl_!�,S�{�CQU  Ch14G�T0 k� �؂�܂!Q8D"%d1O   ��O   � < ��W�E�8E�tA#�Bh_!�,S�{�CQU  ChA0H�T0 k� �����!Q8D"%d1O  	 )�O   � < ��W�E�0E�lA�Bh_!�,S�{�CQU  ChA0H�T0 k� ����!Q8D"%d1O  	 ��O   � < ��S�E�,E�hA�Bd`!�,S�{�CQU  ChA0H�T0 k� �����!Q8D"%d1O  	 ��O   � < ��S�E�$E�`A�Bd`!�,S�{�CQV  ChA0I�T0 k� �����!Q8D"%d1O   ��O   � < ��S�E� E�\	A�B`a!�,S�{�CQV  ShA0I�T0 k� ���� �!Q8D"%d1O   ��O   � < ��O�E�D�T
A�B`a!�,S�{�CQV  ShA0I�T0 k� ����!Q8D"%d1O   ��O   � < ��O�E�D�P0��B`b!�,S�{�CQV  ShA0I�T0 k� ����!Q8D"%d1O   ��O   � < ��O�E�D�H0��B\b!�,S�{�CaV  Sh	10I�T0 k� ����!Q8D"%d1O   ��O   � < ��O�E�D�D0��B\b!�,U"{�CaV  Sh	10I�T0 k� ��!Q8D"%d1O   ��O   � < ��K�E� D�@0��BXc!�,U"{�CaV  Sh
10J�T0 k� � ~�$~!Q8D"%d1O   ��O   � < ��K�E��E�80��BXc|,U"{�CaV  Sh10J�T0 k� �(~�,~!Q8D"%d1O   ��O   � < ��K�E��E�40��BXc|,U"{�CaV  Sh10J��T0 k� �0}�4}!Q8D"%d1O   ��O   � < ��K�E��E�00��BTd|,U"{�CaV  Sh a0J��T0 k� �8|�<|!Q8D"%d1O   ��O   � < ��O�E��E�(0��BTd|,U"{�Ca V  Sh a,J��T0 k� �<{�@{!Q8D"%d1O   ��O   � < ��O�E��E�$@��BTd|,U"{�Ca V  Sh a,J��T0 k� �D{�H{!Q8D"%d1O   ��O   � < ��O�E�� E� @��BPe|,U"{�Ca V  ch a,J��T0 k� �Lz�Pz!Q8D"%d1O   ��O   � < ��O�E��!E�@��BPe|,U"{�Ca V  ch a,J��T0 k� �Ty�Xy!Q8D"%d1O   ��O   � < ��S�E��!E�@��BPe|,@�{�C`�V  ch�,J��T0 k� �\x�`x!Q8D"%d1O   ��O   � < ��S�E��"E�@��BLf|,@�{�Cp�V  ch�0J��T0 k� �`x�dx!Q8D"%d1O   ��O   � < ��S�F �#F  @��BLf|,@�{�Cp�U  ch�0J��T0 k� �hw�lw!Q8D"%d1O   ��O   � < ��W�F �$F "@��BLf|,@�{�Cp�U  ch�0J��T0 k� �pv�tv!Q8D"%d1O   ��O   � < ��W�F �%F #@��BLf|,@�{�Cp�T  ch�0J��T0 k� �xu�|u!Q8D"%d1O   ��O   � < ��[�F �&F  %@��BLf|,E�{�Cp�T  ch�0J��T0 k� �u��u!Q8D"%d1O   ��O   � < ��[�F �'F�'@��BLf|,E�w�E �S  ch�4J��T0 k� �t��t!Q8D"%d1O    ��O  � < ��_�F �)F�(@��BLf|,E�w�E �S  ch�4J��T0 k� �s��s!Q8D"%d1O    ,�O   � < ��c�F �*F�*@��BLf|,E�w�E �R  ch�8J��T0 k� �r��r!Q8D"%d1O    ��O   � < ��g�F �+F�,P��RLf|,E�w�E �R  3h�8K��T0 k� �r��r!Q8D"%d1O    ��O   � < ��g�F �,F�-P��RLf|,E�w�E �Q  3h�8K��T0 k� Ӥq��q!Q8D"%d1O    ��O   � < ��k�F �-F�/P��RLf|,E�w�E �Q  3h �<K��T0 k� Ӭp��p!Q8D"%d1O   �O    � < ��o�F �.F�1P�RLf|,E�s�E �P  3h"�@L��T0 k� Ӱp��p!Q8D"%d1O   �O    � < ��s�E��0F�3P{�RLf|,E�s�E �O  3h#@L��T0 k� Ӹo��o!Q8D"%d1O   ��O    � < ��w�E��1E��40w��Lf|,E�s�E �O  3h$DL��T0 k� ��n��n!Q8D"%d1O   ��O    � < ��{�E��2E��60s��Lf|,As�@`�N  3h&DM��T0 k� �m��m!Q8D"%d1O   ��O   � < ���E��3E��80o��Lf|,As�@`�M  3h'HM��T0 k� �m��m!Q8D"%d1O   ��O    � < ����E��4E��:0k��Lf|,Ao�@`�M  3h(LM��T0 k� �l��l!Q8D"%d1O   ��O    � < ����B��5E��;0g��Lf|,Ao�@`�L  3h*PN��T0 k� �k��k!Q8D"%d1O   ��O    � < ����B��6E��=�c��Lf|,Ao�@`�L   �h+TN��T0 k� �j��j!Q8D"%d1O   ��O    � < ����B��8E��>�_��Lf|,Ao�@`�K   �h,XN��T0 k� ��j��j!Q8D"%d1O   ��O    � < ����B��9E��@�[��Lf|,Ao�@`�K   �h-XN��T0 k� ��i��i!Q8D"%d1O   ��O    � < ����B��:B��A�W��Lf|,Ak�@`�J   �h.\O��T0 k� ��h� h!Q8D"%d1O   ��O    � < ����B��;B��C�S��Lf|,Ak�@`�I   �h0 `O��T0 k� � g�g!Q8D"%d1O   ��O    � < ����B��<B��D�O�BLf|,Ak�@`�I  3h1 dO��T0 k� �g�g!Q8D"%d1O   ��O    � < ����B��=B��F�K�BLf|,Ak�@`�H  3h2 hP��T0 k� �f�f!Q8D"%d1O   ��O    � < ����B��>B��G�G�BLf|,Ak�@`�H  3h3 lP��T0 k� �e�e!Q8D"%d1O   ��O    � < ����B��?B��I�C�BLf|,Ak�@`�G  3h5 pP��T0 k� � d�$d!Q8D"%d1O   ��O    � < ����B��@B��J�?�BLf|,Ag�@`�G  3h6 tP��T0 k� �$d�(d!Q8D"%d1O   ��O    � < ����B��AB��L�;�BLf|,Ag�@`�F  3h7 xQ��T0 k� �,c�0c!Q8D"%d1O   ��O    � < ����B��AB��M�;�BLf|,Ag�@`�F  3h9 |Q��T0 k� �4b�8b!Q8D"%d1O    ��O    � < ����B��BB��N�7�BLf|,Ag�@`�E  #h: �Q��T0 k� �<a�@a!Q8D"%d1O    ��O    � < ����B��CB��P�3�BLf|,Ag�@`�E  #h< �Q��T0 k� �Da�Ha!Q8D"%d1O    ��O    � < ����B��DB��Q�/�BLf|,Ag�@`�E  #h= �R��T0 k� �H`�L`!Q8D"%d1O    /�O    � < ���B��EB��R�+�BLf|,Ac�@`�D  #h> �R��T0 k� �P_�T_!Q8D"%d1O    ��O    � < ���B��FB��S�+�BLf|,Ac�@`�D  #h@ �R� T0 k� �X_�\_!Q8D"%d1O    ��O    � < ���B��GB��U�'�BLf|,Ac�@`�C  #lA �R� T0 k� �`^�d^!Q8D"%d1O    ��O    � < ���B��GB��V�#�BLf|,Ac�@`�C  #lC �S� T0 k� �h]�l]!Q8D"%d1O    ��O    � < ���B��HB��W��BLf|,Ac�@`�B  #lD �S� T0 k� �l\�p\!Q8D"%d1O    ��O    � < ���B��IB��X��BLf|,Ac�@`�B  #lF �S� T0 k� �t\�x\!Q8D"%d1O    ��O    � < ���B��JB��Y��BLf|,Ac�@`�B  #pG �S� T0 k� �|[��[!Q8D"%d1O    ��O    � < ���B��KB� Z��BLf|,A_�@`�A  pI �S� T0 k� �Z��Z!Q8D"%d1O    *�O    � < � �B��KB�\��BLf|,A_�@`�A  tJ �T� T0 k� �Y��Y!Q8D"%d1O    .�O    � < � �B��LB�]��BLf|,A_�@`�@  tL �T� T0 k� �X��X!Q8D"%d1O    ��O    � < � �B��MB�^��BLf|,A_�@`�@  tM �T� T0 k� �V��V!Q8D"%d1O    ��O    � < ��B��NB�_��BLf|,A_�@`�@  xO �T� T0 k� �U��U!Q8D"%d1O    ��O    � < ��B��NB�`��BLf|,A_�@`�?   xP �T� T0 k� �T��T!Q8D"%d1O    ��O    � < �'�B��OB�a��BLf|,A_�@`�?   |Q �U�T0 k� �R��R!Q8D"%d1O    ��O    � < �+�B��PB�b��BLf|,A[�@`�?   |S �U�T0 k� �Q��Q!Q8D"%d1O    ��O    � < �3�B��PB� c��BLf|,A[�@`�>   |T �U�T0 k� �P��P!Q8D"%d1O    ��O    � < �;�B��QB�$d���BLf|,A[�@`�>   �U �U�T0 k� ��N��N!Q8D"%d1O   ��O    � < �?�B��RB�,e���BLf|,A[�@`�=   �V �U�T0 k� ��M��M!Q8D"%d1O   ��O    � < �G�B��RB�0f�� BLf|,A[�@`�=   �X �V�T0 k� ��L��L!Q8D"%d1O   ��O    � < �O�B��SB�4g�� BLf|,A[�@`�=   �Y �V�T0 k� ��J��J!Q8D"%d1O    ��O    � < �S�B� TB�8h��BLf|,A[�@`�<   �Z �V�T0 k� ��I��I!Q8D"%d1O    ��O    � < �[�L�TB�@i��BLf|,A[�@`�<   �[ �V�T0 k� ��H��H!Q8D"%d1O    ��O    � < � c�L�UB�Dj��BLf|,A[�@`�<   �] �V�T0 k� ��G��G!Q8D"%d1O    ��O    � < � g�L�VB�Lj��rLf|,AW�@`�<   �^ �V�T0 k� ��E��E!Q8D"%d1O    ��O    � < � o�L�VB�Pk��rLf|,AW�@`�;   �_ �W�T0 k� ��D��D!Q8D"%d1O    ��O   � < � w�L�WB�Tl��rLf|,AW�@`�;   �` �W�T0 k� ��C��C!Q8D"%d1O    ��O    � < � {�L� WB�\m��rLf|,AW�@`�;   �a �W�T0 k� ��A��A!Q8D"%d1O    ��O    � < � ��L�(XB�`n��rLf|,AW�@`�:   �b �W�T0 k� ��@��@!Q8D"%d1O    ��O    � < � ��L�,XK�ho��rLf|,AW�@`�:   �c �W�T0 k� ��?��?!Q8D"%d1O    ��O    � < � ��L�0YK�lp��rLf|,AW�@`�:   �d �W�T0 k� ��>��>!Q8D"%d1O    ��O    � < � ��L�4ZK�tp��rLf|,AW�@`�:   �e �X�T0 k� ��<��<!Q8D"%d1O    ��O    � < � ��L�<ZK�xq��rLf|,AW�@`�9   �f �X�T0 k� ��;��;!Q8D"%d1O    ��O    � < � ��L�@[K��r��rLf|,AW�@`�9   �g �X�T0 k� ��:��:!Q8D"%d1O    ��O    � < ���L�D[K��s��rLf|,AS�@`�9   �h �X�T0 k� ��8��8!Q8D"%d1O    ��O    � < ���L�H\K��s��rLf|,AS�@`�8   �i �X�T0 k� ��7��7!Q8D"%d1O    ��O    � < ���L�L\K��t��	rLf|,AS�@`�8   �j �X�T0 k� ��6��6!Q8D"%d1O    ��O    � < ���L�P]K��u��	rLf|,AS�@`�8   �k �X�T0 k� ��5��5!Q8D"%d1O    ��O    � < ����L�X]K��v��
�Lf|,AS�@`�8   �l �Y�T0 k� ��3��3!Q8D"%d1O    ��O    � < ����L�\^K��v��
�Lf|,AS�@`�7   �m �Y�T0 k� ��2��2!Q8D"%d1O    ��O    � < ����L�`^K��w���Lf|,AS�@`�7   �n �Y�T0 k� ��1��1!Q8D"%d1O    ��O    � < ����L�d_K��x���Lf|,AS�@`�7   �o �Y�T0 k� ��0��0!Q8D"%d1O    ��O    � < ����L�h_K��x���Lf|,AS�@`�7   �p �Y�T0 k� ��/��/!Q8D"%d1O    ��O    � < ����L�l_K��y?��Lf|,AS�@`�7   �q �Y�T0 k� ��-��-!Q8D"%d1O    ��O    � < ����L�p`K��z?��Lf|,AS�@`�6   �q �Y�T0 k� ��,��,!Q8D"%d1O    ��O    � < ����L�t`K��z?��Lf|,AS�@`�6   �r �Z�T0 k� ��+��+!Q8D"%d1O    ��O    � < ����L�xaK��{?��Lf|,AS�@`�6   �s �Z�T0 k� ��*��*!Q8D"%d1O    ��O    � < ����L�|aK��{?��Lf|,AO�@`�6   �t �Z�T0 k� ��(��(!Q8D"%d1O    ��O    � < ����L��bK��|/��Lf|,AO�@`�5   �u �Z�T0 k� ��'��'!Q8D"%d1O    ��O    � < ����B��bK��}/��Lf|,AO�@`�5   �u �Z�T0 k� ��&��&!Q8D"%d1O    ��O    � < ���B��bK��}/��Lf|,AO�@`�5   �v �Z�T0 k� ��%��%!Q8D"%d1O    ��O    � < ���B��cK��~/��Lf|,AO�@`�5   �w �Z�T0 k� ��$��$!Q8D"%d1O    ��O    � < ���B��cK��~/��Lf|,AO�@`�5   �x �Z�T0 k� ��"��"!Q8D"%d1O    ��O    � < ���B��dK��/��Lf|,AO�@`�4   �x  Z�T0 k� ��!��!!Q8D"%d1O    ��O    � < ���B��dK��/��Lf|,AO�@`�4   �y  [�T0 k� �� �� !Q8D"%d1O    ��O    � < ���B��dK��/��Lf|,AO�@`�4   �z  [�T0 k� ����!Q8D"%d1O    ��O    � < ���B��eK��/��Lf|,AO�@`�4   �{ [�T0 k� ����!Q8D"%d1O    ��O    � < ��'�B��eK��/��Lf|,AO�@`�4   �{ [�T0 k� ����!Q8D"%d1O    ��O    � < ��+�B��eK����Lf|,AO�@`�3   �| [�T0 k� ����!Q8D"%d1O    ��O    � < ��/�B��fK��~��Lf|,AO�@`�3   �} [�T0 k� ����!Q8D"%d1O    ��O    � < ��0 B��fK��~��Lf|,AO�@`�3   �} [�T0 k� ����!Q8D"%d1O    ��O    � < ��4B��fK��~��Lf|,AO�@`�3   �~ [�T0 k� ����!Q8D"%d1O    ��O    � < ��8B��gK� ~��Lf|,AO�@`�3   � [�T0 k� ����!Q8D"%d1O    ��O    � < ��<B��gK�}���Lf|,AK�@`�3   � [�T0 k� ����!Q8D"%d1O    ��O    � < ��@B��gK�}���Lf|,AK�@`�2   �� \�T0 k� ����!Q8D"%d1O    ��O    � < ��DB��hK�}���Lf|,AK�@`�2   �� \�T0 k� ����!Q8D"%d1O    ��O    � < ��HB��hK�}���Lf|,AK�@`�2   � \�T0 k� ����!Q8D"%d1O    ��O    � < ��LB��hK�}���Lf|,AK�@`�2   � \�T0 k� ����!Q8D"%d1O    ��O    � < ��PB��iK�|���Lf|,AK�@`�2   � [�T0 k� ����!Q8D"%d1O    ��O    � < ��TB��jK�|�� �Lf|,AK�@`�2   � [�T0 k� ����!Q8D"%d1O    ��O    � < ��XB��jK�|��!�Lf|,AK�@`�2   �~ [�T0 k� ����!Q8D"%d1O    ��O    � < ��\B��kK� |��"�Lf|,AK�@`�1   �~ [�T0 k� ����!Q8D"%d1O    ��O    � < ��`B��kK�$|��"�Lf|,AK�@`�1   �~ [�T0 k� ����!Q8D"%d1O    ��O    � < ��`	B�lK�${��#�Lf|,AK�@`�1   �~ [�T0 k� ��
��
!Q8D"%d1O    ��O    � < ��d	B�lK�({��$�Lf|,AK�@`�1   �}  Z�T0 k� ��	��	!Q8D"%d1O    ��O    � < ��h
B�mK�,{��$�Lf|,AK�@`�1   �}  Z�T0 k� ����!Q8D"%d1O    ��O    � < ��l
B�mK�,{��%�Lf|,AK�@`�1   �}  Z�T0 k� ����!Q8D"%d1O    ��O    � < ��pB�nK�0{��&�Pf|,AK�@`�1   �}  Z�T0 k� ����!Q8D"%d1O    ��O   � < ��tB�oK�4z��&�Pf|,AK�@`�0   �}  Z�T0 k� ����!Q8D"%d1O    ��O    � < ��tB�oK�8z��'rTe|,AK�@`�0   �| $Z�T0 k� ����!Q8D"%d1O    ��O    � < ��xB�pK�8z��(rTe|,AK�@`�0   �| $Z�T0 k� ����!Q8D"%d1O    ��O    � < ��|B�$qK�<z��(rXe|,AK�@`�0   �| (Y�T0 k� ����!Q8D"%d1O    ��O    � < ���B�(qK�@z��)rXe|,AK�@`�0   �| (Y�T0 k� �� �� !Q8D"%d1O    ��O   � < ���B�,rK�@z��)r\d|,AK�@`�0   �{ ,Y�T0 k� ������!Q8D"%d1O    ��O    � < ���B�0sK�Dy��*r\d|,AK�@`�0   �{ ,Y�T0 k� ������!Q8D"%d1O    ��O    � < ���B�8sK�Dy��+B`d|,AG�@`�0   �{ ,Y�T0 k� ������!Q8D"%d1O    ��O    � < ���B�<tK�Hy��+B`d|,AG�@`�0   �{ 0Y�T0 k� ������!Q8D"%d1O    ��O    � < ���B�DtK�Ly��,Bdd|,AG�@`�/   �{ 0X�T0 k� ������!Q8D"%d1O    ��O    � < ���B�HuK�Ly��,Bdc|,AG�@`�/   �{ 0X�T0 k� ������!Q8D"%d1O    ��O    � < ���B�PuK�Py��-Bdc|,AG�@`�/   �z 4X�T0 k� ������!Q8D"%d1O    ��O    � < ���B�TvB�Py��-Bhc|,AG�@`�/   �z 4X�T0 k� ������!Q8D"%d1O    ��O    � < ���E�\wB�Tx��.Bhc|,AG�@`�/   �z 4X�T0 k� ������!Q8D"%d1O    ��O    � < ���E�`wB�Xx��.Blc|,AG�@`�/   �z 8X�T0 k� ������!Q8D"%d1O    ��O    � < ���E�hxB�\x��/Blb|,AG�@`�/   �z 8X�T0 k� ������!Q8D"%d1O    ��O    � < ���E�pxB�\x��/Bpb|,AG�@`�/   �z 8W�T0 k� ������!Q8D"%d1O    ��O    � < ���E�tyB�`x��0Bpb|,AG�@`�/   �y <W�T0 k� ������!Q8D"%d1O    ��O    � < ��E�|yB�dx��0Bpb|,AG�@`�/   �y <W�T0 k� ������!Q8D"%d1O    ��O    � < ��E��zB�hx��1Btb|,AG�@`�.   �y <W�T0 k� ������!Q8D"%d1O    ��O    � < ��E��zB�lx��1Bta|,AG�@`�.   �y @W�T0 k� ������!Q8D"%d1O    ��O    � < ��E��{B�pw��2Bta|,AG�@`�.   �y @W�T0 k� ������!Q8D"%d1O    ��O    � < ��E��{B�tw��2Bxa|,AG�@`�.   �y @W�T0 k� ������!Q8D"%d1O    ��O    � < ��E��|B�xw��3Bxa|,AG�@`�.   �x DW�T0 k� ������!Q8D"%d1O    ��O    � < ��E��|B�|w��3B|a|,AG�@`�.   �x DW� T0 k� ������!Q8D"%d1O    ��O    � < ��E��|B��w��4B|a|,AG�@`�.   �x DV� T0 k� ������!Q8D"%d1O    ��O    � < ��E��}B��w��4B|`|,AG�@`�.   �x DV� T0 k� ������!Q8D"%d1O    ��O    � < ���E��}B��w��4B�`|,AG�@`�.   �x HV� T0 k� ������!Q8D"%d1O    ��O    � < ���L��}B��w��5B�`|,AG�@`�.   �x HV� T0 k� ������!Q8D"%d1O    ��O    � < ���L��}B��v��5B�`|,AG�@`�.   �x HV� T0 k� ������!Q8D"%d1O    ��O    � < ��L��~B��v��6B�`|,AG�@`�-   �w LV� T0 k� ������!Q8D"%d1O    ��O    � < ��L��~B��v��6B�`|,AG�@`�-   �w LV� T0 k� ������!Q8D"%d1O    ��O    � < ��L��~B��v��6B�_|,AG�@`�-   �w LV� T0 k� ������!Q8D"%d1O    ��O    � < ��L��~B��v��7B�_|,AG�@`�-   �w LV� T0 k� ������!Q8D"%d1O    ��O    � < ��L��B��v��7B�_|,AG�@`�-   �w PV� T0 k� ������!Q8D"%d1O    ��O    � < �� L��B��v��8B�_|,AG�@`�-   �w PU� T0 k� ������!Q8D"%d1O    ��O    � < ��!L� B��v��8B�_|,AG�@`�-   �w PU� T0 k� ������!Q8D"%d1O    ��O    � < ��"L�B��v��8B�_|,AG�@`�-   �w PU� T0 k� ������!Q8D"%d1O    ��O    � < ��#L��B��v��9B�_|,AG�@`�-   �v TU� T0 k� ������!Q8D"%d1O    ��O    � < ��$L�B��u��9B�^|,AG�@`�-   �v TU� T0 k� ������!Q8D"%d1O    ��O    � < ��%L�B��u��9B�^|,AG�@`�-   �v TU� T0 k� ������!Q8D"%d1O    ��O    � < ��&L� B��u��:B�^|,AG�@`�-   �v TU� T0 k� ������!Q8D"%d1O    ��O    � < � 'L�$B��u��:B�^|,AG�@`�-   �v TU� T0 k� ������!Q8D"%d1O    ��O    � < �)L�,~B��u��:B�^|,AG�@`�-   �v XU� T0 k� ������!Q8D"%d1O    ��O    � < �*L�0~B��u��;B�^|,AG�@`�-   �v XU� T0 k� ������!Q8D"%d1O    ��O    � < �+L�4~B��u��;B�^|,AG�@`�,   �v XU� T0 k� ������!Q8D"%d1O    ��O    � < �"-L�@}B�u��<B�]|,AG�@`�,   �v \T� T0 k� ������!Q8D"%d1O    ��O    � < �" .L�H}B�u��<B�]|,AG�@`�,   �u \T� T0 k� ������!Q8D"%d1O    ��O    � < �"$/L�L}B�u��<B�]|,AC�@`�,   �u \T� T0 k� ������!Q8D"%d1O    ��O    � < �",1L�P}B�u��=B�]|,AC�@`�,   �u \T� T0 k� ������!Q8D"%d1O    ��O    � < �"02L�X|B�$u��=B�]|,AC�@`�,   �u \T� T0 k� ������!Q8D"%d1O    ��O    � < �83L�\|B�,t��=B�]|,AC�@`�,   �u `T� T0 k� ������!Q8D"%d1O    ��O    � < �<4L�`|B�4t��>B�]|,AC�@`�,   �u `T� T0 k� ������!Q8D"%d1O    ��O    � < �D5L�h|B�<t��>B�]|,AC�@`�,   �u `T� T0 k� ������!Q8D"%d1O    ��O   � < �L6E�l|B�Dt��>B�]|,AC�@`�,   �u `T� T0 k� ������!Q8D"%d1O    ��O    � < �P7E�p{B�Lt��>B�]|,AC�@`�,   �u `T� T0 k� ������!Q8D"%d1O    ��O    � < ��X8E�t{B�Tt��?B�\|,AC�@`�,   �u `T� T0 k� ������!Q8D"%d1O    ��O    � < ��`9E�|{B�\t��?B�\|,AC�@`�,   �u dT� T0 k� ������!Q8D"%d1O    ��O    � < ��d:E��zB�dt��?B�\|,AC�@`�,   �t dT�!T0 k� ������!Q8D"%d1O    ��O    � < ��l;E��zB�lt��?B�\|,AC�@`�,   �t dT�!T0 k� ������!Q8D"%d1O    ��O    � < ��t<E��zB�tt��@B�\|,AC�@`�,   �t dS�!T0 k� ������!Q8D"%d1O    ��O    � < ��|=E��yE�|t��@B�\|,AC�@`�,   �t dS�!T0 k� ������!Q8D"%d1O    ��O    � < ���=E��yE��t� @B�\|,AC�@`�,   �s dS�!T0 k� ������!Q8D"%d1O    ��O    � < ���>E��yE��t� @B�\|,AC�@`�,   �s hS�!T0 k� ������!Q8D"%d1O    ��O    � < ���?E��yE��t�AB�\|,AC�@`�+   �s hS�!T0 k� ������!Q8D"%d1O    ��O    � < ���@E��yE��t�AB�\|,AC�@`�+   �r hS�!T0 k� ������!Q8D"%d1O    ��O    � < ���ALӐxE��s�AB�\|,AC�@`�+   �r hS�!T0 k� ������!Q8D"%d1O    ��O    � < ���BLӔxE��s�AB�[|,AC�@`�+   �r hS�!T0 k� ������!Q8D"%d1O    ��O    � < ���CLӔxE��s�BB�[|,AC�@`�+   �q hS�!T0 k� ������!Q8D"%d1O    ��O    � < ���CLӘxE��s�BB�[|,AC�@`�+   �q lS�!T0 k� ������!Q8D"%d1O    ��O    � < ���DLӘxE��s�BB�[|,AC�@`�+   �q lS�!T0 k� ������!Q8D"%d1O    ��O    � < ���ELӜwB��s�BB�[|,AC�@`�+   �q lS�!T0 k� ������!Q8D"%d1O    ��O    � < ���FL�wB��r�CB�[|,AC�@`�+   �p lS�!T0 k� ������!Q8D"%d1O    ��O    � < ���GL�wB��r�CB�[|,AC�@`�+   �p lS�!T0 k� ������!Q8D"%d1O    ��O   � < ���HL�wB��r�CB�[|,AC�@`�+   �p lS�!T0 k� ������!Q8D"%d1O    ��O    � < ���IL�wB��r�Cr�[|,AC�@`�+   �p lS�!T0 k� ������!Q8D"%d1O    ��O    � < ���IL�wB��q�Cr�[|,AC�@`�+   �o pS�!T0 k� ������!Q8D"%d1O    ��O    � < ���JL�vB��q�Dr�[|,AC�@`�+   �o pS�!T0 k� ������!Q8D"%d1O    ��O    � < ���KL�vB�q�Dr�[|,AC�@`�+   �o pS�!T0 k� ������!Q8D"%d1O    ��O    � < ���LL�vCp�Dr�[|,AC�@`�+   �o pS�!T0 k� ������!Q8D"%d1O    ��O    � < �� ML�vCp� Dr�Z|,AC�@`�+   �o pR�!T0 k� ������!Q8D"%d1O    ��O    � < ��NLӰvCo� Dr�Z|,AC�@`�+   �n pR�!T0 k� ������!Q8D"%d1O    ��O    � < ��OLӰvC$o�$Dr�Z|,AC�@`�+   �n pR�!T0 k� ������!Q8D"%d1O    ��O    � < ��PLӴuC,n�$Er�Z|,AC�@`�+   �n pR"!T0 k� ������!Q8D"%d1O    ��O    � < �	3PLӴuE�4n�$Er�Z|,AC�@`�+   �n tR"!T0 k� ������!Q8D"%d1O    ��O    � < �	3 QLӸuE�<m�(Er�Z|,AC�@`�+   �m tR"!T0 k� ������!Q8D"%d1O    ��O    � < �	3$RLӸuE�Dm�(Er�Z|,AC�@`�+   �m tR"!T0 k� ������!Q8D"%d1O    ��O    � < �	3,RLӼuE�Hl�(Er�Z|,AC�@`�+   �m tR"!T0 k� ������!Q8D"%d1O    ��O    � < �	30SLӼuE�Pl�,Fr�Z|,AC�@`�+   �m tR"!T0 k� ������!Q8D"%d1O    ��O    � < �	C4SL��uE�Xk�,F��Z|,AC�@`�+   �m tR"!T0 k� ������!Q8D"%d1O    ��O    � < �	C8TCC�tE�`k�,F��Z|,AC�@`�+   �l tR"!T0 k� ������!Q8D"%d1O    ��O    � < �	C<TCC�tE�hj�0F��Z|,AC�@`�+    l tR"!T0 k� ������!Q8D"%d1O    ��O    � < �	C@TCC�tE�pi�0F��Z|,AC�@`�+    l tR"!T0 k� ������!Q8D"%d1O    ��O    � < �	CDUCC�sE�xi�0F��Z|,AC�@`�+    l xR"!T0 k� ������!Q8D"%d1O    ��O    � < �	3HUCC�sE��h�4F��Z|,AC�@`�+   l xR�!T0 k� ������!Q8D"%d1O    ��O    � < �	3LUE��sE��g�4G��Z|,AC�@`�+   k xR�!T0 k� �����!Q8D"%d1O    ��O    � < �	3PUE��rE��f�4G��Z|,AC�@`�*   k xR�!T0 k� �����!Q8D"%d1O    ��O    � < �	3TVE��rE��e�8G��Z|,AC�@`�*   k xR�!T0 k� �����!Q8D"%d1O    ��O    � < �	3XVE��qE��d�8G��Y|,AC�@`�*   k xR�!T0 k� �{���!Q8D"%d1O    ��O    � < ��XVE��pKӠc�8G��Y|,AC�@`�*   k xR�!T0 k� �{���!Q8D"%d1O    ��O    � < ��\VE��pKӠc�8G��Y|,AC�@`�*   j xR�!T0 k� �w��{�!Q8D"%d1O    ��O    � < ��`VE��pKӤa�<H��Y|,AC�@`�*   j xR�!T0 k� �w��{�!Q8D"%d1O    ��O    � < ��dVE��pKӨ`�<H��Y|,AC�@`�*   j xR�!T0 k� �w��{�!Q8D"%d1O    ��O    � < ��dWE��pKӰ_�<H��Y|,AC�@`�*   j xR�!T0 k� �s��w�!Q8D"%d1O    ��O    � < ��hWE��oKӴ^�@H��Y|,AC�@`�*   j |R�!T0 k� �s��w�!Q8D"%d1O    ��O    � < ��lWE��oKӸ]�@H��Y|,AC�@`�*   j |R"$!T0 k� �o��s�!Q8D"%d1O    ��O    � < ��lWE��nKӼ\�@H��Y|,AC�@`�*   i |R"$!T0 k� �o��s�!Q8D"%d1O    ��O    � < ��pWE��nK��[�@H��Y|,AC�@`�*   i |R"$!T0 k� �o��s�!Q8D"%d1O    ��O    � < ��tWE��mK��Z�DH��Y|,AC�@`�*   i |R"$!T0 k� �k��o�!Q8D"%d1O    ��O    � < ��xXE��lK��Y�DI��Y|,AC�@`�*   i |R"$!T0 k� �k��o�!Q8D"%d1O    ��O    � < ��xXE��lK��X�DI��Y|,AC�@`�*   i |R"$!T0 k� �g��k�!Q8D"%d1O    ��O   � < ��|XE��kK��V�DI��Y|,AC�@`�*   i |R"$!T0 k� �g��k�!Q8D"%d1O    ��O    � < ��|XE��kK��V�HI��Y|,AC�@`�*   h |Q"$!T0 k� �c��g�!Q8D"%d1O    ��O    � < �ÀXE��jK��U�HI��Y|,AC�@`�*   h |Q"$!T0 k� �c��g�!Q8D"%d1O    ��O    � < �ÄXC��jK��T�HI��Y|,AC�@`�*    h |Q"$!T0 k� �c��g�!Q8D"%d1O    ��O    � < �ÄXC��iK��S�LI��Y|,AC�@`�*    h |Q"$!T0 k� �_��c�!Q8D"%d1O    ��O    � < �ÈYC��iK��R�LI��Y|,AC�@`�*    h �Q�!T0 k� �_��c�!Q8D"%d1O    ��O    � < �ÈYC��hK��Q�PI��Y|,AC�@`�*   $h �Q�!T0 k� �[��_�!Q8D"%d1O    ��O    � < �ÌYC��hK��P�PJ��Y|,AC�@`�*   $g �Q�!T0 k� �[��_�!Q8D"%d1O    ��O    � < �ÐYC��gK��O�TJ��Y|,AC�@`�*   $g �Q�!T0 k� �W��[�!Q8D"%d1O    ��O    � < �ÐYC�gK��N�TJ��Y|,AC�@`�*   (g �Q�!T0 k� �W��[�!Q8D"%d1O    ��O    � < �ÔYC�gK��M�XJ��Y|,AC�@`�*   (g �Q�!T0 k� �S��W�!Q8D"%d1O    ��O    � < �ÔYC�gK� L�\J��Y!�,AC�@`�*   (g �Q�!T0 k� �S��W�!Q8D"%d1O    ��O    � < �ÔXC�gK�L�\J��Y!�,AC�@`�*   (g �Q�"T0 k� �S��W�!Q8D"%d1O    ��O    � < �ÔXC�gK�K�`J��Y!�,AC�@`�*   ,g �Q�"T0 k� �O��S�!Q8D"%d1O    ��O    � < �ØXC�gK�J�dJ��X!�,AC�@`�*   ,g �Q�"T0 k� �O��S�!Q8D"%d1O    ��O    � < �ØWC�gK�I�hJ��X!�,AC�@`�*   ,f �Q�"T0 k� �K��O�!Q8D"%d1O    ��O    � < �ØWC�gK�H�lJ��X!�,AC�@`�*   ,f �Q�"T0 k� �K��O�!Q8D"%d1O    ��O    � < �ØWC�gK�H�lK��X!�,AC�@`�*   0f �Q�"T0 k� �G��K�!Q8D"%d1O    ��O    � < �ØWC�gK�G�pK��X!�,AC�@`�*   0f �Q�"T0 k� �G��K�!Q8D"%d1O    ��O    � < �ÜVC�gK�F�tKr�X!�,AC�@`�*   0f �Q�"T0 k� �C��G�!Q8D"%d1O    ��O    � < �ÜVEC�gK�E�xKr�X!�,AC�@`�*   0f �Q�"T0 k� �C��G�!Q8D"%d1O    ��O    � < �ÜVEC�gK� E�xKr�X!�,AC�@`�*   4f �Q�"T0 k� �?��C�!Q8D"%d1O    ��O    � < � �BrdE_�1+��I!�,E��E�  B��%��H"s�T0 k� ����!Q8D"%d1O    �� 
  � 6 � �BrdEg�1'��I!�,E��E�  %r��%��H"s�T0 k� ����!Q8D"%d1O    �� 
  � 6 � �BrdE�o�1��I!�,E��E�  %r��%��H"s�T0 k� ����!Q8D"%d1O    �� 
  � 6 � �BrdE�w�1��I!�,E��E�  %r��%��H"s�T0 k� ����!Q8D"%d1O    �� 
  � 6 � �H�dE�{�1��I|,E���E�  %r��%��H3�T0 k� ����!Q8D"%d1O    ��   � 6 � �H�dE���1��I|,E���E�  %r��%��H3�T0 k� ����!Q8D"%d1O    ��   � 6 � �H�hE���1��J|,E���E�  %r��%��H3�T0 k� �|��!Q8D"%d1O    ��   � 5 � �H�hE���!��J|,E���E�  %r��%��I3�T0 k� �x�|!Q8D"%d1O    ��   � 5 � �H�hE���!��J|,E���E�  %r��%��I3�T0 k� �x�|!Q8D"%d1O    ��   � 5 � �H�hE��� ���J|,E���E�  %r��%��I3�T0 k� �x�|!Q8D"%d1O    ��   � 5 � a�H�lE��� ���J|,E���@��  %r��%��I3�T0 k� �x�|!Q8D"%d1O    ��   � 5 � a�H�lE��� ���J|,E���@��  %r��%��I3�T0 k� �|��!Q8D"%d1O    ��   � 5 � a�H�lEs�� ���J|,E���@��  %r��%��I3�T0 k� �|��!Q8D"%d1O    ��   � 5 � a�H�pEs�� ���J|,E���@��  %r��%��I3�T0 k� �|��!Q8D"%d1O    ��   � 5 � a�H�pEs������J|,E���@��  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 5 � a�H�pEs������J|,D���A�  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 4 � a�H�tEs������J|,D���A�  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 4 � a�H�tEs������J|,D���A�  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 4 � a�H�tEs������J|,D���A�  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 4 � a�H�tEs������J|,D���A�  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 4 � a�H�xEs������J|,D���C��  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 4 � a�H�xEs�� ���J|,D���C��  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 4 � a�H�xEs�� ���J|,D���C��  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 3 � a�H�xEc�� ���J|,D���C��  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 3 � a�H�|Ed� ���J|,D���C��  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 3 � a�H�|Ed� ���J|,D���A�  %r��%��I3�T0 k� ����!Q8D"%d1O    $�   � 3 � a�H�|Ed� ���J|,D���A�  %r��%��I3�T0 k� 2���!Q8D"%d1O    ��   � 3 � a�H�|Ed� ���J|,D���A�  %r��%��I3�T0 k� 2���!Q8D"%d1O    ��   � 3 � a�H�|
Ed�� �J|,D���A�  %r��%��I3�T0 k� 2���!Q8D"%d1O    ��   � 2 � a�HҀ
Ed���J|,D���A�  %r��%��I3�T0 k� 2���!Q8D"%d1O    ��   � 2 � a�HҀ
Ed#���J|,D���E2�  %r��%��I3�T0 k� 2���!Q8D"%d1O    ��   � 2 � a�HҀ	Ed'���J|,D���E2�  %r��%��I3�T0 k� ����!Q8D"%d1O    ��   � 1 � a�HҀ	Ed+���|J|,E��E2�  C�%��I3�T0 k� ����!Q8D"%d1O    ��   � 1 � a�HҀ	ET/����|J|,E��E2�  C�%��I3�T0 k� ����!Q8D"%d1O    ��   � 1 � a�H�	ET3����|J|,E��E2�  C�%��I3�T0 k� ����!Q8D"%d1O    ��   � 1 � a�H�ET7����|J|,E��E2�  C�%��I3�T0 k� ����!Q8D"%d1O    ��   � 0 � a�H�ET7����|J|,E��E2�  C�%��I3�T0 k� ����!Q8D"%d1O    �   � 0 � a�H�ET;���	�|J|,E��E2�  3���I3�T0 k� ����!Q8D"%d1O   ��   � 0 � a�H�ET?���
�|J|,F��E2�  3���I3�T0 k� ����!Q8D"%d1O   ��   � 0 � a�H�ET?����|J|,F��E2�  3��I3�T0 k� ����!Q8D"%d1O   ��   � 0 � a�H�ETC����|J|,F��E2�  3��I3�T0 k� ��!Q8D"%d1O   �   � 0 � a�H�C�C���SxJ|,F��E2|  3��I3�T0 k� �� !Q8D"%d1O   ��   � 0 � a�H�C�G���StJ|,F��E2|  C�S�I3�T0 k� �4�8!Q8D"%d1O   ��   � 0 � a�H�C�G���SpJ|,Dџ�E2|  C�S�I)��T0 k� �L�P!Q8D"%d1O   ��   � 0 � a�I�C�G���SpJ|,Dџ�CB|  C�S�I)��T0 k� �d�h!Q8D"%d1O   ��   � 0 � a�I�C�G���SlJ|,Dћ�CB|  C�S�I)��T0 k� �|��!Q8D"%d1O   ��   � 0 � a�I�C�G���ShJ|,Dћ�CBx  C�S�I)��T0 k� ����!Q8D"%d1O   ��   � 0 � a�I�E�G���SdJ|,Dћ�CBx   ��S�I)��T0 k� ����!Q8D"%d1O  	 $�   � 0 � a�I�E�G���SdK|,Dћ�CBx   ��S�I)��T0 k� ì��!Q8D"%d1O  	 ��   � 0 � a�I�E�G���c`K|,Dћ�CBx   ��S�I)��T0 k� è��!Q8D"%d1O  	 ��   � 0 � a�I�E�G���c\K|,Dћ�CBx   ��S�I)��T0 k� è��!Q8D"%d1O   ��   � 0 � a�I�E�G���c\K|,Dћ�CBx   ��S�I)��T0 k� è��!Q8D"%d1O   ��   � 0 � a�I�A�G�� cXK|,Dћ�CBx  #�S�I)��T0 k� è��!Q8D"%d1O   ��   � 0 � a�I�A�G��cTK|,Dџ�CBx  #�S�I)��T0 k� è��!Q8D"%d1O   ��   � 0 � a�I�A�G��cTK|,D��CBx  #�S�I)��T0 k� Ӥ��!Q8D"%d1O   ��   � 0 � a�I� A�G��cPK|,D��@�x  #�S�I)��T0 k� Ӥ��!Q8D"%d1O   ��   � 0 � a�I� A�G��sLK|,D��@�x  #�S�I)��T0 k� Ӥ��!Q8D"%d1O   ��  � 0 � a�I��A�G��sLK|,D��@�x  ��S�I)��T0 k� Ӥ��!Q8D"%d1O   ��   � 0 � a�I��A�G��sHK|,D��@�x  ��S�I)��T0 k� Ӥ��!Q8D"%d1O   ��   � 0 � a�I��A�G� sHK|,F��@�x  ��S�I)��T0 k� ���!Q8D"%d1O   ��   � 0 � a�I��A�C�$sDK|,F��E"x  ��S�I)��T0 k� ���!Q8D"%d1O   ��   � 0 � a�I��A�C�,s@K|,F��E"x  ��S�I)��T0 k� ���!Q8D"%d1O   ��   � 0 � a�I��A�C�0s@K|,F��E"|  ��S�H)��T0 k� ���!Q8D"%d1O   ��   � 0 � a�Dҗ�ATC�4s<K|,F��E"|  ��S�H)��T0 k� ���!Q8D"%d1O   ��   � 0 � a�Dҗ�AT?�<s<K|,F��E"|  �#�S|H)��	T0 k� ���!Q8D"%d1O   ��   � 0 � a�Dҗ�AT?�@s8K|,F��E�|  �#�SxH)��	T0 k� � �� !Q8D"%d1O   ��   � 0 � a�Dҗ�AT?�Hs8K|,E���E�|  �#�SxH)��	T0 k� �!��!!Q8D"%d1O   ��   � 0 � a�Dқ�AT;��Ls4K|,E���E�|  �'��tH)��	T0 k� �"��"!Q8D"%d1O   ��   � 0 � a�Dқ�C�;��Ts0K|,E��E�|  �'��tH)��	T0 k� �"��"!Q8D"%d1O   ��   � 0 � a�Dқ�C�7��Xs0L|,E��E�|  �'��pH)��	T0 k� �#��#!Q8D"%d1O   ��   � 0 � a�Dҟ�C�3��` s,L|,E��E�|  �'��lH)��	T0 k� �$��$!Q8D"%d1O   ��   � 0 � a�Dң�C�3��d s,L|,I�E�|  �'��lH)��	T0 k� �%��%!Q8D"%d1O   ��   � 0 � a�Dң�C�/�	�h s(L|,I�E�|
  �'��lH)��	T0 k� �&��&!Q8D"%d1O    ��   � 0 � a�Dҧ�C�+�	�l!s(L|,I�E�|
  �'��hH)��	T0 k� �&��&!Q8D"%d1O    ,�   � 0  a�Dҧ�C�'�	�t!s$L|,I�E�|	  �'��dH)��	T0 k� Ә'��'!Q8D"%d1O    ��   � 0  a�D��C�'�	�x!s$L|,I�	E�|  �'��dH)��	T0 k� Ӕ(��(!Q8D"%d1O    ��   � 0  a�D��C�#�	�|!s L|,I!�
E�x  �'��`G)��	T0 k� Ӕ)��)!Q8D"%d1O    ��   � 0  a�D��C��
�!sL|,I!�E�x  �'��\G3�	T0 k� Ӕ*��*!Q8D"%d1O   ��   � 0  a�D��C��
�!sL|,I!�E�x  �'��\G3�	T0 k� Ӕ*��*!Q8D"%d1O   ��   � 0  a�D��C��
�!sL|,I!�E�t  �'��XF3�	T0 k� �+��+!Q8D"%d1O   ��   � 0  a�D��C��
�!sL|,I!�E�t  �'��XF3�	T0 k� �,��,!Q8D"%d1O   ��   � 0  a�D��C��
�!sL|,B��E�p  �'��TE3�
T0 k� �-��-!Q8D"%d1O   ��   � 0 � a�D���C��	�!sL|,B��E�p  �#��PE�
T0 k� �-��-!Q8D"%d1O   ��   � 0 � a�D���C��	�!sM|,B��E�l  �#�sLC�
T0 k� t+�x+!Q8D"%d1O   ��   � 0 � a�D���C���	�!sM|,B��E�h  ��sHC�T0 k� �h*�l*!Q8D"%d1O   ��   � 0 � a�D���C���	�!sM|,E��E�d  ��sDB�T0 k� �`*�d*!Q8D"%d1O   ��   � 0 � a�D���D��
�!sM|,E��E�d  ��sDA�T0 k� �\)�`)!Q8D"%d1O   ��   � 0 � a�D�� D��
�!sM|,E��E�`  ��s@@�T0 k� �T(�X(!Q8D"%d1O   ��   � 0 � a�D�� D��
�!sM|,E��E�\  ��s<@�T0 k� �L'�P'!Q8D"%d1O   ��   � 0 � a�D��D��
�!s M|,SQ�E�X   ��s8>�T0 k� �H&�L&!Q8D"%d1O   �   � 0 � a�D��D����!r�M|,SQ�E�T   ��s8=�T0 k� �H%�L%!Q8D"%d1O   ��   � 0 �                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��� ]�+V+U � �� VR   � �
	  � �~�     Vil �N�    ���            l	 Z �          ��    ���  H
!
          gi�  T T    � �b�     g�� �+�    ���   	           Z �         b     ��� 8�           E�  � �	   �v     Eؘ�    ��          E Z �         H`�    ���  	@	           Kn�   � 4      ��     KX- ?�    UM            Z  Z �           �@�     ���  H$
          X��   � �    . �fj     X�U �S�    ��   
          H  Z �         n�    ���  (

          �  
     B�V[     ��V[                  	         �����         �    
  ���      0            ����        V ��    ���� ��    ��                   )��                ��@   0	%           *u       j >��     *w� >��    ��                   ?��          �  �  ��@   8
          �T�      ~  ��    �T�  ��               ��       	 � !         �       ��F   0
 
          f+g           �	�     fH���    �Hy                	    �         	  ��     ��H   P
           Q�,          � �!     Q�� ��    �� �                  �         
  �p     ��B   P	          "� ��      �l�     "�l�                             ���3             �  ��@    P                   ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��4#  ��        ��    ����$�    �{��                  x                j  �   �   �                         ��    ��       �      ��             "                                                 �                          � �  �� � >   ���  	          
     
  d  �  ���K       ;� `^@ <� _  <� _  <�  _@ ��  a� �� ]`��� ����  ����. ����< ����J ����X � �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0� ���� � 
�\ U� 
� V  
�| V  
�\ W� 
�� W� 
�\ W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���� �  <���)  ������  
�fD
��L���"����D" � j  "  B   J jF�"    "�j * , ����
��"     �j @�    �
� �  �  
�  W    ��     � �  �    X    ��     � �       f��  ��     �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �O      ��+T ���        �T ���        �        ��        �        ��        �    ��    ��  ��        ��                         襩 4 � ���                                     �                 ����            W ����%��   < ��� 7 w           �EDM Verbeek son     0:00                                                                        2  2      �kV t7k^ dc� �C. �C6	 C9 �C: � �B� � 	B� � 
B�  �B�  � B� � B� �J� � J� � J� �J�* � c� � �c� � � c� � �K �K	  � K �K  �K � �c�# �	� � �	� � �� � �� � "�   "�"!"�"*� �#"� � $"�, �%� �&
�)  '*QL  ()�T )*\ � **RT �+*&\ �,*6d �-* l � .*Od � /*Kd � 0*Jt �1)�d �2* |3)�tO 4*KdO 5*Jt_ )�dO  *Et_  *AdO 9*Et_  *Ad[ )�wT *2�G )�pI )�p;  *J� � 
�                                                                                                                                                                                                                 �� P        �     @ 
              h P E h  ���� F   	            	�������������������������������������� ���������	�
��������                                                                                          ��    �g�� ��������������������������������������������������������   �4, =� * �� ���	�@����0���[	�                                                                                                                                                                                                                                                                                                                                 M @����                                                                                                                                                                                                                                  -        �	�  H�J      �j                             �������������������������������������������������������                                                                                                                                   o       d              �     � l          
 	  
	 
 	 	 ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ���         	   �              c    1    � �  D�J    	  6�  	                           ������������������������������������������������������                                                                                                                                        �             ^        �        x      �    	  
 	 
 	 	 ���������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������           #                                                                                                                                                                                                                                      
                                                                        �             


           �   }�                                       O	                           +                     ����������������  '{������������  +'����������������    ��������������������  '{�������������������������ww�ww333wwwwwwww�ww�ww�ww�ww333wwww A C 6                	                 � ���F �^@       |3b�T�q�$Hb2�                                                                                                                                                                                                                                                           )n)h1p  Y	n                                                    m           ��                                                                                                                                                                                                                                                                                                                                                                                                    � � �  � ��  � ��  � <��  �  ��  EZmX  �N \�����i�����F�����������������'����������X^          <   4 
 ����          	�   & AG� �  s   
           �2�                                                                                                                                                                                                                                                                                                                                     p C B   �     p   !             !��                                                                                                                                                                                                                            Y   �� �~ ��      �� ?      ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ������������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������   �� @     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    7      ;      ��                       X     �  �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��  p���� �$ ^h  ��     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@     | 
hv ��  | 
hv �$ ^$   l ^@ ;� �� ^@ ;� �$  �  ��  �      �      &�����������J   g���         f ^�         �� � <      &      ���~�������J���J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �   3       �  �3 3�=������<��̼��� �3 33==ƙ�<ə�ƙ�3ƙ��ƙ���i� 3= ��3=�l�ә��<��l<��l<��l<���<    �   3=  �30 ��� ���=��������                        +   3     0  �<  3� 3� =� =� 0� 0������������������3�33033�0�3�0��;f��;��̽�������3��3��<���<�f���̳=�=�������3303<�<00�<30�3����������������=��=��3�3�=�3�0  �=  �3  �3� ��0 ̳0 �0 �0  0� =� =� 3�  3�  �<  0  33�0�3�0�3�0�3303�303�303�303303��<���0<��0<033<033003300330033030�30�<00�<0330333033303330333033�0��<���0�03303303=03=03��0 ̳0 ��0 �3� �3� �=  0  3�     �                           <�03=��3=�� 3��  �=  �        033003300330�330��303= ��33    330333033303330333<��333ݰ    0=�0<3���;�3 �=  3�             �                           wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           " """ "!   " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             " """ "!   " ""  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                            " ""   "" !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                       "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ���"�!/"�  �                                                                                                                                                                                   �� ���
�������˽������̽�]��+I۲"T�""T32.T33>@4C CDT �E@ ��  ʐ  �       "   "�� � ��� �wp ��� �vz �w� �����˻���˰�̰� ��  ��  ��� � �+ �+ �  .   "�   �   �   �    � ��  �                     �  �˰ ���                 ��  ��  ���           U   U  U  U  	T  ,� ,� "  " "  ��  �              �   � � �  ��� ��  �      �   �  �  �  �   �  �  �   �  �                                                �          �       �                        �   ��  ���  � �    �                                                                                                                                                     � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �         ��                                 � ���� ��   � � �                            ����                  �   �� �       �  �  ��  �   �   �   �                                                    � ̻ �ۼͺ�	ۚ����C�˽T;��UJ��ET�35J�D3T�  ̰ ̻	�̻���w������wv��wpʨ� ��� ��� ��  "�� .� "�� ��0 "          �  �  ��  �   �         �  �� ʝ ,��+� "" "��CEJ�D5J� J�  �� 
�� �  �� �+� �"" """����    �        �   �   � ���� �� ����                    �� ��������p��}`     �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��  ��  ���                        "  "  "                                                                                                                                                                  �� ̽ ̽��۽ }�  wz  � ��������ɜ���̚��̸ ��  ��  �  �  T�  T�  H� �E �E �D�[ ˻  ˸  ��  
� ,"�"" �"  �"              "   *�  ��� ��� �ة��ڋ�̽� ��  ��  ̻� ̻� ��� ��@ ��@ DD0 T30 B3� ��  ��  ��  
� +� �"" �"� �" ��� ����  ��          ���    �                       
 "� ""� ""� "                       �                             ���                         �  ��                    �����                                             ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �      �  �                                             �  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �        ��  ̽  ��  }�  ��  ��� ̼� �ܚ��٩�����̽�̽��˹�.��""��"�3��33� 33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �                          �     �     �   �   �   �   �   �                      	   	   	   	�" �!  �  �� �   �                �  �� Ș ��  ��  �                        �   �   ��  ���   ˰  ̹  ��@ ��UP�EEXDTD�    �   ��  ���  � �    �                                                                                                                                                     �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �     �   �     �   �        �                       �  �   ��  �   ��  �  �   �  �  �  �  �   �   �   �  �  �  �  �   �  �  �   �   ��  �                            �   ���                            �   �    �                                                                                                                   	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                      �   �                              �   �                      �������  ���    �        � ��                    ���� �                           �   ��  ���  � �    �                                                                                                                                       ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r`ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                       ���� ��� ����                            �    � �  ��                  ���                              �   ���                            �   �                                                                                                    �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �   �   �   ˰  ˙  ɪ  ��� ټ� �̰ �̰ ��� ��  ��                              ��          �  ��� ̻� ��� rbp wgz�               �������  ���    �                    ��  ��  ���   ���� �                                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �   �   �   ˰  ˙  ɪ  ��� ټ� �̰ �̰ ��� ��  ��  �   �   �                                       �                        ���� ��� ����                            �    � �  ��                  ���                                                                                                                                                                                           �  ��� ܽи�؀  � ˚ �̹�̹�˹�˻ܻ��ܘ��܉���D���U�D�J�N T�� D�  T�  �  ��  �� �� ,ث"���"��� ���۝� {�� ��  ��� ��(�������� ˸� ɀ  ��  ��� �̀ �̈ �� ���虎�(���"��� ��� � �/�����              �   �   �   �   �   �� (���+�����"/  ��                    �� ��� ��� ��  �                         �   �                    �          �         �   �  �  �   �               �   �                     �                             �   �   �   �   �   �                                                                                                                                                �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������    <     = 8 0 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>108(=((( (<���������������� L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L����������������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7����������������  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqkV t7k^ dc� �C. �C6	 C9 �C: � �B� � 	B� � 
B�  �B�  � B� � B� �J� � J� � J� �J�* � c� � �c� � � c� � �K �K	  � K �K  �K � �c�# �	� � �	� � �� � �� � "�   "�"!"�"*� �#"� � $"�, �%� �&
�)  '*QL  ()�T )*\ � **RT �+*&\ �,*6d �-* l � .*Od � /*Kd � 0*Jt �1)�d �2* |3)�tO 4*KdO 5*Jt_ )�dO  *Et_  *AdO 9*Et_  *Ad[ )�wT *2�G )�pI )�p;  *J�3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������#� ��9�K�Z�X��5�R�O�S�G� � � � � � � � � � �/�.�7����������������������������������������� ��5�K�\�O�T��=�U�J�J� � � � � � � � � � �/�.�7�����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������2�0�.� ���������������������������������������/�.�7�	�
�������������������� � � � � � �����������������������������������������%��������������������/�.�7� �� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�A�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                