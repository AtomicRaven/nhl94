GST@�                                                            \     �                                               6���      �  �            ����e ����J�����������x�������        �g      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"     �j�
�   ��
  3�                                                                              ����������������������������������       ��    =b? 0Q0 45 118  4             	 

    
               ��� �4 �  ��                 nY 
)         8:�����������������������������������������������������������������������������������������������������������������������������o=  0  o4   1  +      '           �                    	�  7�  V�  	�                    
          : �����������������������������������������������������������������������������                                ��  �   �  ��   @  #   �   �                                                                                '    
)nY  
    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E k �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    K�kCSHd30U��<��P|,  �@8( b E pA� f3�T0 k� �K��O�T2e   2$    ��&    �  �K�kCSHd30U��<��P|,  �@8( b E pA� f3�T0 k� �O��S�T2e   2$    ��&    �  �K�kCSHd34U��<��P|,  �@8( bE pA� f3�T0 k� �O��S�T2e   2$    ��&    �  �L�kCSHd34U��<��P|,  �@8( bE pA� f3�T0 k� �S��W�T2e   2$    ��&    �  �L�kCSHd38T��<��P|,  �@8( bE pA� f3�T0 k� �S��W�T2e   2$    ��&    �  �L�k@�Hd38T��<��P|,  �@8( bF pA� f3�T0 k� �W��[�T2e   2$    ��&    �  �L�k@�Hd3<T��<� P|,  �@8( bF pA� f3�T0 k� �W��[�T2e   2$    ��&    �  �L�j@�HdC@T��<� P|,  �@8( bF pA� f3�T0 k� �[��_�T2e   2$    ��&    �  �L�j@�HdC@T��<� P|,  �@8( bF oA� f3�T0 k� �[��_�T2e   2$    ��&    �  �L�j@�HdCDT��<� P|,  �@8( bF oA� f3�T0 k� �_��c�T2e   2$    ��&    �  �L�j@�HdCDS��<� P|,  �@8( bF oA� e3�T0 k� �_��c�T2e   2$    ��&    �  �L�j@�HdCHS��<� P|,  �@8( bF oA� e3�T0 k� �c��g�T2e   2$    ��&    �  �L�j@�HdCHS��<� P|,  �@8( bFoA� e3�T0 k� �c��g�T2e   2$    ��&    �  �L�j@�HdCLS��<  P|,  �@<( bGoA� e3�T0 k� �g��k�T2e   2$    ��&    �  �L�j@�HdCLS��<  P|,  �@<( bGoA� e3�T0 k� �g��k�T2e   2$    ��&    �  �L�j@�HdCPS��<  P|,  �@<( bGoA� e3�T0 k� �g��k�T2e   2$    ��&    �  �L�j@�Hd3PR��<  P|,  #�@<( bGoA� e3�T0 k� �k��o�T2e   2$    ��&    �  �L�j@�Hd3TR��<  P|,  #�@<( b GoA� e3�T0 k� �k��o�T2e   2$    ��&    �  �L�j@�Hd3TR��<  P|,  '�@<( b GoA� e3�T0 k� �o��s�T2e   2$    ��&    �  �L�j@�Hd3XR��<  P|,  '�@<( b GnA� e3�T0 k� �o��s�T2e   2$    ��&    �  �L�j@�Hd3XR��<  P|,  '�@<( b$GnA� e3�T0 k� �o��s�T2e   2$    ��&    �  �L�j@�Hd3\R��< c P|,  +�@<( b$GnA� e3�T0 k� �s��w�T2e   2$    ��&    �  �L�j@�Hd3\R��< c P|,  +�@<( b$GnA� e3�T0 k� �s��w�T2e   2$    ��&    �  �L�j@�Hd3`R��< c P|,  /�@<( b(GnA� e3�T0 k� �w��{�T2e   2$    ��&    �  �L�j@�Hd3`Q��< c P|,  /�@<( b(HnA� e3�T0 k� �w��{�T2e   2$    ��&    �  �L�j@�Hd�dQ��< c Q|,  /�@<( b,HnA� e3�T0 k� �w��{�T2e   2$    ��&    �  �L�j@�Hd�dQ��<�Q|,  3�@<( b,HnA� e3�T0 k� �{���T2e   2$    ��&    �  �L�j@�Hd�hQ��<�Q|,  3�@<( b,HnA� e3�T0 k� �{���T2e   2$    ��&    �  �L�j@�Hd�hQ��<�Q|,  3�@@( b0HnA� e3�T0 k� �{���T2e   2$    ��&    �  �L�j@�Hd�hQ��<�R|,  7�@@( b0HnA� e3�T0 k� �����T2e   2$    ��&    �  �L�j@�Hd�lQ� <�R|,  7�@@( b0HnA� e3�T0 k� �����T2e   2$    ��&    �  �L�j@�Hd�lQ� <�R|,  7�@@( b4HnA� d3�T0 k� �����T2e   2$    ��&    �  �L�j@�Hd�pP�<�S!�,  ;�@@( b4HmA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�pP�<�S!�,  ;�@@( b4HmA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�pP�<S!�,  ;�@@( b4HmA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�tP�<T!�,  ;�@@( b8ImA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�tP�<T!�,  ?�@@( b8ImA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�tP�<T!�,  ?�@@( b8ImA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�xP�<T!�,  ?�@@( b<ImA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�xP�<�T!�,  C�@@( b<ImA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�xP�<�U!�,  C�@@( b<ImA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�|P�<�U!�,  C�@@( b@ImA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�|O�<�U!�,  C�@@( b@ImA� d3�T0 k� ������T2e   2$    ��&    �  �L�j@�Hd�|O�<�U|,  G�@@( b@JmA� d3�T0 k� ������T2e   2$    ��&    �  �K�j@�Hd��O�<�U|,  G�@@( bDJmA� d3�T0 k� ������T2e   2$    ��&    �  �K�j@�Hd��O�<�U|,  G�@@( bDJmA� d3�T0 k� ������T2e   2$    ��&    �  �K�j@�Hd��O�<�U|,  K�@D( bDJmA� d3�T0 k� ������T2e   2$    ��&    �  �K�j@�Hd��O� <�U|,  K�@D( bHJmA� d3�T0 k� ������T2e   2$    ��&    �  �E.  I�˩	�`QM8*]ü#3��[�C�D}� OA�+C�Dl"s�T0 k� ������T2e   2$    ��D    ����;E.�I�é	�XQM4(]��#3��S�C�<}��MA|+C�@k"s�T0 k� ������T2e   2$    ��D    ����;E-��I���	�PQM,%]���3��C�C�(}�JAp*C�0j"s�T0 k� �s��w�T2e   2$    ��D    ����;E��I���	�LPM$#]���3�M;�C� }�HAh*C�,i"s�T0 k� �k��o�T2e   2$    ��D    ����;E��I���	�DPM "]���3�M/�C�}�FQ`)C�$i3�T0 k� �c��g�T2e   2$    ��D    ����;E��I���	�@PM ]���3�M'�C�}�EQX)C�h3�T0 k� �_��c�T2e   2$    ��D    ����;E��I���	�<PM]���3�M�C�}�CQT(C�g3�T0 k� �W��[�T2e   2$    ��D    ����;E��I���	�8P]]���3�M�C��}�AQL'C�f3�T0 k� �O��S�T2e   2$    ��D    ����;E��I���	�4P]]��3�M�C��}�?QD'C�e3�T0 k� �G��K�T2e   2$    ��D    ����;E��I���	�4P]]{��3�M�C��}�>Q<&C� e3�T0 k� �C��G�T2e   2$    ��D    ����;E��I���	�0P]]s��3�L��C��}�<Q4%C��d3�T0 k� �;��?�T2e   2$    ��D    ����;E��I���	�(P\��g��3�L��D�}�8Q$$C��b3�T0 k� �3��7�T2e   2$    ��D    ����;E��I���	�(P\��_��3�<��D�}��7Q#C��a3�T0 k� �/��3�T2e   2$    ��D    ����;E��I���	�$P	���W��3�<��D�}��5Q"C��`3�T0 k� �+��/�T2e   2$    ��D    ����;E���I���	� P	���S��3�<��D�}��3a"C��_"��T0 k� �'��+�T2e   2$    ��D    ����;E���I���	� P	���K��3�<��D�}��2a!C��^"��T0 k� �#��'�T2e   2$    ��D    ����;E���I���	�P	���C��/�<��D�~��0a  C��]"��T0 k� ���#�T2e   2$    ��D    ����;E���I���	�P	���;��/�<��D�~��.`�C��\"��T0 k� ����T2e   2$    ��D    ����;E���I���	�P	���3��/�<��D�~��-`�C��["��T0 k� ����T2e   2$    ��D    ����;D���I���	�P	��
�#��/�<��D�~��*`�C��X"��T0 k� �����T2e   2$    ��D    ����;D��I���	�P	��	���/�<��Dt~��(`�C��W"��T0 k� ������T2e   2$    ��D    ����;D��I���	�P	�����/�<��Dl~��&`�C��V"��T0 k� ����T2e   2$    ��D    ����;D��I���	�P	�����/�<��Dd~��%`�C��U"��T0 k� ����T2e   2$    ��D    ����;D��I���	�P	�����/�,{�D\~��#`�C��T"��T0 k� �ߵ��T2e   2$    ��D    ����;D��I���	�P	������/�,s�DP~��"0�C��S3�T0 k� �׳�۳T2e   2$    ��D    ����;D��I���	�P	������/�,k�DH~��!0�C�xQ3�T0 k� �ϱ�ӱT2e   2$    ��D    ����:D��I���	�P	������/�,c�D@~��0�C�pP3�T0 k� �ǰ�˰T2e   2$    ��D    ����9D��I���	�P	������+�,_�D8~��0�C�lO3�T0 k� ����ïT2e   2$    ��D    ����8D��I���	�P	������+�,W�D,~��0�E@dN3�T0 k� ������T2e   2$    ��D    ����8D��A���	�P	������+�,G�D~����E@TK3�T0 k� ������T2e   2$    ��D    ����8D��A���	�P	�����+�,?�C�~����E@LJ3�T0 k� ������T2e   2$    ��D    ����8D��A���	�P	̼����'�,;�C�~����E@DI3�T0 k� ������T2e   2$    ��D    ����8D�#�A���	�P	̼����'�\3�C� ~���xE@<H3�T0 k� ������T2e   2$    �D    ����8D�'�A���	�P	̼ ����#�\3�C��~���pE@4G3�T0 k� ������T2e   2$    ��D    ����8D�'�BN���P	�� ����#�\+�C��~���lE@0E3�T0 k� ������T2e   2$    ��D    ����8D�+�BN���P	�� �����\'�C��~���dE@(D3�T0 k� ������T2e   2$    ��D    ����8D�/�BN���P	��������\#�C��~���\E@ C3�T0 k� ������T2e   2$    ��D    ����8D�3�BN���P	��������\�C��~���T
E0A3�T0 k� ������T2e   2$    ��D    ����8D�7�BN���P	��������\�C��~���P	E0@3�T0 k� ������T2e   2$    �D    ����@D�?�@��NP	̿��s���\�EM�~���@E0=3�T0 k� ����îT2e   2$   ��O    ����HD�C�@��NP	̿��k���l�EM�~���8E?�<3�T0 k� �˯�ϯT2e   2$   ��O    ����OD�G�@��NP	̿��c���l�EM�~��
�4E?�;3�T0 k� �۰�߰T2e   2$   ��O    ����VD�K�@��NP	̿��[���k��EM�~��	�,E?�93�T0 k� ����T2e   2$   ��O    ����]D�O�@��NP	̿��W���k��EM�~� �$E?�83�T0 k� ������T2e   2$   ��O    ����dD�S�B����P����O���k��EM�~�� E?�63�T0 k� ����T2e   2$   ��O    ����jD�W�B����P����G���k��EM�~�� E?�53�T0 k� ����T2e   2$   ��O    ����pD�[�B����P����C���k��EMx}���E?�33�T0 k� �#��'�T2e   2$   ��O    ����vE[�B����P����;���{��EMp}���E?�23�T0 k� �/��3�T2e   2$   ��O    ����|E_�B����P����3���{��EMh}���E/�03�T0 k� �?��C�T2e   2$   ��O    �����Ec�B����P����/���{��C�`|� �E/�/3�T0 k� �K��O�T2e   2$   ��O    �����Eg�B����P����'���{��C�T|�$��E/�-3�T0 k� �[��_�T2e   2$   ��O    �����Ek�B����P����#���{��C�L|�( ��E/�,3�T0 k� �g��k�T2e   2$   ��O    �����Eo�B���� P�������{��C�D{�/���E/�*3�T0 k� �w��{�T2e   2$   ��O    �����Es�B���� P�������{��C�<{�7���E/�(3�T0 k� ������T2e   2$   ��O    �����Ew�B����$PL������{��EM0{�;���E/�'3�T0 k� ������T2e   2$   ��O    �����E{�B����(PL������{��EM(z�C���E/�%3�T0 k� ������T2e   2$   ��O    �����E�B����,PL������{��EM z�G���E/�#3�T0 k� ������T2e   2$   ��O    �����E��B����0PL�������{��EMy�O���E/�"3�T0 k� ������T2e   2$   ��O    �����E��B����0PL�������{��EMy�W���E/� 3�T0 k� ������T2e   2$   ��O    �����E��B����4P�������{��EMx�[���E�3�T0 k� ������T2e   2$   ��O    �����E��B����8P�������{��E<�w�c����E�3�T0 k� ������T2e   2$   ��O    �����E��B����<P�����|�{��E<�w�k����E�3�T0 k� ������T2e   2$   ��O    �����E��B����@P�����|�{��E<�v�o����E�3�T0 k� ����T2e   2$   ��O    �����E��B�ǩ�HP����ߵ|�{��E<�u�w����E�3�T0 k� ����T2e   2$    ��O    �����E��B�˩�LP����۵|�{��E<�u�����E�3�T0 k� ���#�T2e   2$    ��O    �����E��B�ϩ�PP����״|�{��E<�t������E�3�T0 k� �+��/�T2e   2$    ��O    �����E��B�ө�TP����Ӵ|�{��E<�s������B��3�T0 k� �;��?�T2e   2$    /�O    �����E��B�ש�XP����˴|#�{��E<�r������B��3�T0 k� �G��K�T2e   2$    ��O    �����E��B�ߩ�`P����ǳ|#�{��E<�q������B��3�T0 k� �W��[�T2e   2$    ��O    �����E��B���dP����ó|#�{��E<�p������B��3�T0 k� �c��g�T2e   2$    ��O    �����E��B���hP������|#�{��E<�o������B��3�T0 k� �o��s�T2e   2$    ��O    �����E��B���pP������|#�{��E,�n������B��3�T0 k� �����T2e   2$    ��O    �����E��B���tP������|'�{��E,�m������B��3�T0 k� ������T2e   2$    ��O    �����E��B����|P������|'�{��E,�l������B��
3�T0 k� ������T2e   2$    ��O    �����E��B���΀P������|'�{��E,�k������B��	3�T0 k� ������T2e   2$    ��O    �����E��B��ΈP������|'�{��E,�j������B��3�T0 k� ������T2e   2$    ��O    �����E��B��ސP�����|'�{��E,�h������B��3�T0 k� ������T2e   2$    ��     �����B^��B��ޔP�����|'�{��E,�g������B��3�T0 k� ������T2e   2$    ��     �����B^��B��ޜP�����|+�{��E,|f������B��3�T0 k� ������T2e   2$    ��     �����B^��B��ޤP�����|+�{��E,xe������B��3�T0 k� ������T2e   2$    ��     �����B^��B�'�ިP�����|+�{��E,td�����B��3�T0 k� ������T2e   2$    ��     �����B^��B�/�ްP�����|+�{��Epb����B�� 3�T0 k� ������T2e   2$    ��     �����B^��B�3�޸P�����|+�{��Ela����B���3�T0 k� ������T2e   2$    ��     �����B^��B�;���P�����|+�{��Eh`����B���3�T0 k� ������T2e   2$    ��     �����B^��B�C���P������|+�{��Ed_����B���3�T0 k� ������T2e   2$    ��     �����B^��B�K���P������|+�{��E`^�'����B���3�T0 k� ������T2e   2$    ��     �����B^��B�S���P������|+�{��E\\�/����E��3�T0 k� �����T2e   2$    ��     �����B^��B�_���P������|+�{��EXZ�?����E��3�T0 k� ����T2e   2$    ��     ���  Bn��B�g���P������|+�{��ETY�G����E��3�T0 k� ����T2e   2$    ��     ��� Bn��B�o���P������|+�{��B�TX�O����E��3�T0 k� ����T2e   2$    ��     ��� Bo�B�w���P������|+�{��B�TW�W����E��3�T0 k� ����T2e   2$    ��     ��� Bo�B���P������|+�{��B�PV�_����E��3�T0 k� ����T2e   2$    ��     ��� Bo�B����P������|+�{��B�PU�g����E��3�T0 k� ���#�T2e   2$    ��     ��� E��B����P������|+�{��B�PT�o����E��3�T0 k� �'��+�T2e   2$    ��     ��� E��B���� P������|+�{��B�PS�w���E��3�T0 k� �+��/�T2e   2$    ��     ��� E��B����(P������|+�{��B�LR���E���3�T0 k� �/��3�T2e   2$    ��  
   ��� E�#�B����0P�����|+�{��B�LQ��
@�E���3�T0 k� �7��;�T2e   2$    ��  
   ��� 	E�'�B����<P�����|+�{��B�LP��
@�E���3�T0 k� �;��?�T2e   2$    ��  
   ��� 
E�/�B����DP�����|+�{��B�LO��
@�E���3�T0 k� �?��C�T2e   2$    ��  
   ��� E�3�B����LP�����|+�{��B�PN��
@�E���3�T0 k� �G��K�T2e   2$    ��  
   ��� E7�B�ǩ�TP�����|+�{��B�PM��
@�E���3�T0 k� �G��K�T2e   2$    ��  
   ��� EC�B�ө�hP�����|+�{��B�PK�� #�E���3�T0 k� �S��W�T2e   2$    ��  
   ��� EG�B�۩�pP�����|+�{��B�TJ�� '�E���3�T0 k� �W��[�T2e   2$    ��  
   ��� EO�B���xP�����|/�{��B�TJ�� +�E���3�T0 k� �[��_�T2e   2$    ��  
   ��� FS�B����P�����|/�{��B�TI�� +�E���3�T0 k� �g��k�T2e   2$    ��  
   ��� FW�B����P�����|/�{��B�XH�� /�E���3�T0 k� �w��{�T2e   2$    ��  
   ��� F[�B����P�����|/�{��B�XGo��03�B���3�T0 k� �����T2e   2$    ��  
   ��� Fc�B�����P�����|/�{��B�\Fo��0;�B���3�T0 k� ������T2e   2$    ��  
   ��� Fg�B�����P�����|/�{��B�`Eo��0?�B���3�T0 k� ������T2e   2$    ��  
   ��� Ek�B����P�����|/�{��B�`Eo��0C�B���3�T0 k� ������T2e   2$    ��  
   ��� Es�B����P ����|/�{��B�dDo��0K�B��3�T0 k� �� �� T2e   2$    ��  
   ��� Ew�B����P ����|/�|�B�hCo��0O�B��3�T0 k� ����T2e   2$    ��  
   ��� E{�B����P ����|/�|�B�lBo��0S�B��3�T0 k� ����T2e   2$    �  
   ��� H��B����P ��ǜ|/�|�B�pA`�0_�B��3�T0 k� ��
��
T2e   2$    �� 
   ���  H��E����P ��˜|/�|�B�t@`�0c�B�'�3�T0 k� ����T2e   2$    �� 
   ��� $H��E����P ��Ϝ|/�|�B�x?`�0g�B�/�3�T0 k� ����T2e   2$    �� 
   ��� (H��E����P ��Ӝ|/�|�B�|?`�0o�B�7�3�T0 k� ����T2e   2$   �� 
   ��� ,H��E�#���P ��۝|/�|�B̄>P�@s�B�;�3�T0 k� ����T2e   2$   �� 
   ��� 0H��E�'��P ��ߝ|/�|�B̈=P�@w�B�C�3�T0 k� ����T2e   2$   �� 	   ��� 4H���E�/��P ���|/�|�B̌=P�@�B�K�3�T0 k� ����T2e   2$   �� 	   ��� 8H���E�3��P m���|/�|�B̐<P�@��B�S�3�T0 k� � �T2e   2$   �� 	   ��� <H���E�7��P m���|/�|�Bܔ;P#�@��B�[�3�T0 k� � � T2e   2$   �� 	   ��� @H���E�?��$P m���|/�|�Bܜ;P#�@��E�_�3�T0 k� �#�#T2e   2$   �� 	   ��� DH���E�C��,P m���|, |�Bܠ:P'�@��E�g�3�T0 k� � &�$&T2e   2$   ��/ 	   ��� HI��D�G��8P m���|, |�Bܤ9P'�@��E�o�3�T0 k� �,)�0)T2e   2$   ��/ 	   ��� KI��D�O��@P ���|, |�Bܬ9P+�@��E�w�3�T0 k� �8+�<+T2e   2$    ��/ 	   ��� NI��D�S��HP ���|, |�Bܰ8P+�@��E��3�T0 k� �D.�H.T2e   2$    ��/ 	   ��� QI� D�[��PP ���|, |�Bܸ7@+�@��E���3�T0 k� �L1�P1T2e   2$    ��/ 	   ��� TI�D�_��XP ���|, |�Bܼ7@/�P��E���3�T0 k� �X4�\4T2e   2$    ��/ 	   ��� WI�D�g��dP ���|, |�B��6@/�P��DЗ�3�T0 k� �d6�h6T2e   2$    ��/ 	   ��� ZI�D�k�lPM #�|, |�B��6@/�P��DЛ�3�T0 k� �p9�t9T2e   2$    ��/ 	   ��� ]I�D�w�|PM /�|, |�B��5@/�PˏDЫ�3�T0 k� ��?��?T2e   2$    ��/ 	   ��� _I�D���PM3�|, |�B��4@3�PӎDг�3�T0 k� ��C��CT2e   2$    ��" 	   ��� aI�DЃ��PM;�|, |�B��4@3�PیDл�3�T0 k� ��D��DT2e   2$    ��" 	   ��� cI�DЋ��PM?�|, |�B��3@3�PߋD���3�T0 k� ��E��ET2e   2$    ��"    ��� eI�D����PMG�|, |�B��203�P�D���3�T0 k� ��F��FT2e   2$    ��"    ��� gI�	D����PMO�|, |�B��203�P�D���3�T0 k� ��G��GT2e   2$    ��"    �  iI�	D����P]S�|, |�B� 103�P�D���3�T0 k� ��G��GT2e   2$    ��"    �  kI�
Dࣥ�P]�[�|, |�B�103�`��D���3�T0 k� ��G��GT2e   2$    ��"    �  mI�D৥�P]�c�|, |�B�003�a�D���3�T0 k� ��G��GT2e   2$    ��"    �  oI�I���P]�g�|, |�B�0@/�a�D���3�T0 k� ��C��CT2e   2$    ��"    � 	 qI�I���P]�o�|, |�B� 0@/�a�D���3�T0 k� ��@��@T2e   2$    ��"    � 
 sI�I���P]�w�|, |�B�(/@/�a�D��3�T0 k� ��>��>T2e   2$    ��"    �  uI�I���P]�{�|, |�B�0/@/�a�D��3�T0 k� ��=��=T2e   2$    ��"    �  wF J Ǧ��O]���|, ��B�@.@/�+�D��3�T0 k� �<�<T2e   2$    ��"    �  zF J ˦� O]���|, ��B�H-@/�3�D�#�3�T0 k� �;�;T2e   2$    ��"    �  |F J Ϧ�O]���|, ��B�P-@/�;�D�+�3�T0 k� �9� 9T2e   2$    ��"    �  ~F J Ӧ�Om���|, ��B�X,P/�C�D�3�3�T0 k� �$9�(9T2e   2$    ��"    �  �F J ӦQOm	���|, �#�B�d,P/�K�D�;�3�T0 k� �0:�4:T2e   2$    ��"    �  �F I�צQ$Nm	���|, �#�B�l,P/�S�D�G�3�T0 k� �8;�<;T2e   2$    ��"    �  �F I�ۦQ,Nm	���|, �#�B�t+P/�[�D�O�3�T0 k� �@;�D;T2e   2$    ��"    �  �F I�ߦQ4Nm
���|, �#�B�|+P/�c�D�W�3�T0 k� �H<�L<T2e   2$    ��"    �  �E� I��Q<Mm
���|, ,#�B��*P/�k�D�_�3�T0 k� �P;�T;T2e   2$    ��"    �  �E�$I���DMm���|, ,'�B��*P/�s�D�g�3�T0 k� �\:�`:T2e   2$    ��"    �  �E�(J ��LLm�ó|, ,'�B͘*P/�{�D�o�3�T0 k� �d9�h9T2e   2$    ��"    �  �E�,J ��XLm�˳|, ,'�B͠)P/���E�w�3�T0 k� �l7�p7T2e   2$    ��"    �  �E�4J ��`Km�ϴ|, ,'�Bͨ)P/���E��3�T0 k� �t6�x6T2e   2$    ��"    �  �E�8J ��hKm�ӵ|, ,'�Bʹ(P/���E���3�T0 k� �|5��5T2e   2$    ��"    �  �E�<J ��pJ-,۵|, ,+�Bͼ(`/���E���3�T0 k� ��4��4T2e   2$    ��"    �  �E�@I���xJ-,߶|, ,+�B��(`/���E���3�T0 k� ��3��3T2e   2$    ��"    �  �E�HI����I-,�|, ,+�B��'`/���E���3�T0 k� ��3��3T2e   2$    ��"    �  �E�LI����I-,�|, ,+�B��'`/���E���3�T0 k� ��2��2T2e   2$    ��"    �  �E�XI���q�H-,��|, /�B��&`/���E���3�T0 k� ��0��0T2e   2$    ��"    �  �E�\ E���q�G-,��|, /�B��&`/�ǘEq��3�T0 k� ��/��/T2e   2$    ��"    �  �E�d E���q�F�|, 3�B��&0/�Q˙Eq��3�T0 k� ��.��.T2e   2$    ��"    �  �E�h!E���q�E�|, 3�B�%0/�QӚEq��3�T0 k� ��-��-T2e   2$    ��"    �  �E�p"E��q�D�|, 7�B�%0/�QۛEq��3�T0 k� ��,��,T2e   2$    ��"    �  �E�t#E��q�C�|, 7�B�%0/�QߛEq��3�T0 k� ��+��+T2e   2$    ��"    �  �E�|#E��q�B�|, ;�B�$0/�Q�Eq��3�T0 k� ��*��*T2e   2$    ��"    �  �E��$B��q�A��#�|, ?�B�($0/�Q�Eq��3�T0 k� ��)��)T2e   2$    ��"    �  �E�%B��q�@��'�|, ?�B�0$ /�Q�Eq��3�T0 k� ��(��(T2e   2$    ��"    �  �E�&B��q�>�$�7�|, G�B�@# 3�Q��Er�3�T0 k� ��%��%T2e   2$    ��"    �  �E�&B���=�(�?�|, �K�B�H# 3�Q��D��3�T0 k� ��%��%T2e   2$    ��"    �  �E�'B���<�(�C�|, �O�B�T# 3�R�D��3�T0 k� ��%��%T2e   2$    ��"    �  �E�(B�#��;�,�K�|, �S�B�\"�3�B�D��3�T0 k� ��$� $T2e   2$    ��"    �  �B��(B�'� :�0�S�|, �W�B�d"�3�B�D��3�T0 k� ��#� #T2e   2$    ��"    �  �B��)B�/�9�4�[�|, �[�B�l"�7�B�D�'�3�T0 k� �"�"T2e   2$    ��"    �  �B��)B�3��7�8�c�|, �_�B�x"�7�B�D�+�3�T0 k� �!�!T2e   2$    ��"    �  �B��*B�7��6�<�k�|, �g�B��!�7�B�D�0 3�T0 k� �!�!T2e   2$    ��"    �  �B��+B�;��5�@�s�|, �k�B��!�;�B�D�83�T0 k� �!�!T2e   2$    ��"    �  �B��,B�G��(3�H���|, �w�B��!�?�B�D�D3�T0 k� ��T2e   2$    ��"    �  �B��,B�K�r02�L���|, �{�B�� �?�B�D�H3�T0 k� ��T2e   2$    ��"    �  �B��-B�S�r41�T���|, ���B�� �C�B�D�P3�T0 k� ��T2e   2$    ��"    �  �B��-B�W�r<0�X���|, ���B�� �C�2�D�T
3�T0 k� � �$T2e   2$    ��"    �  �B��.B�_�r@/�\���|, ���B��  G�2#�D�\3�T0 k� �$�(T2e   2$    ��"    �  �B�.B�c�rH.�d���|, ���B�� G�2#�D�`3�T0 k� �,�0T2e   2$    ��"    �  �B�/B�k�bL-�h���|, ���B�� K�2'�D�d3�T0 k� �0�4T2e   2$    ��"    �  �B�/B�s�bP,�l���|, ���B�� O�2'�D�l3�T0 k� �4�8T2e   2$    ��"    �  �B�0B�w�bX+�t���|, ���B�� O�2'�Drp3�T0 k� �8�<T2e   2$    ��"    �  �B�$0B��b\+�x���|, ���B�� S�2+�Drt3�T0 k� �<�@T2e   2$    ��"    �  �B�,1B���b\+̀���|, ���B�� W�2+�Dr|3�T0 k� �@�DT2e   2$    �"    �  �E�<1B���Rd-͌���|, �ϜB� [�2/�Dr�3�T0 k� �D�HT2e   2$    �"    �  �E�D2B���Rd.͐���|,  ל@ _� �/�Or�!3�T0 k� �H�LT2e   2$    �"    �  �E�L2B���Rh/͘���|,  ߜ@ c� �3�Or�"3�T0 k� �H�LT2e   2$    ��"    �  �E�T2E���Rl0͠ ���|,  �@  g� �3�Or�$3�T0 k� �L�PT2e   2$    ��"    �  �E�\2E���Rl1ͤ ��|,  �@( `g� �7�Or�%3�T0 k� �P�TT2e   2$    ��"    �  �Ed3E���bp2ͬ ��|,  ��@0 `k� �7�Or�&3�T0 k� �P�TT2e   2$    ��"    �  �El3E���bt3ʹ!��|,  ��@8 `o��7�Or�(3�T0 k� �T �X T2e   2$    ��"    �  �Et3E�ǧbt5ݼ!��|,  �@@ `s��;�Or�)3�T0 k� �T!�X!T2e   2$    ��"    �  �E|4E�ϧbx6��"�'�|,  �@H `s��;�Or�+3�T0 k� �X"�\"T2e   2$    ��"    �  �E�4E�Өbx7��"�/�|,  �@P `w��;�Or�,3�T0 k� �\#�`#T2e   2$    ��"   �  �K��4E�ۨr|8��"�7�|,  �@X `{��?�Or�-3�T0 k� �\$�`$T2e   2$    ��"    �  �K��4E��r|8��#�?�|,  '�@` `{��?�Or�.3�T0 k� �`%�d%T2e   2$    ��"    �  �K��5Eq�r�9��#�G�|,  /�@h `��?�Or�03�T0 k� �`&�d&T2e   2$    ��"    �  �K��5Eq�r�:��#�O�|,  7�@p `���?�Or�13�T0 k� �d'�h'T2e   2$    ��"    �  �K��5Eq��r�;��#�W�|,  ?�@x `���?�Or�23�T0 k� �d(�h(T2e   2$    ��"    �  �K��6Eq����<��$�_�|,  G�@| `���?�Or�33�T0 k� �x%�|%T2e   2$   �"    �  �K��6Er���=� $�g�|,  O�@� `���?�Or�53�T0 k� ��"��"T2e   2$   ��/    �  �K��6Er���>�$�o�|,  W�@� `���?�Or�63�T0 k� ����T2e   2$   ��/    �  �K��6Er���?�%�w�|,  _�@� `���?�Or�73�T0 k� ����T2e   2$   ��/    �  �K��7Er���@�%��|,  g�@� `���?�Os83�T0 k� ����T2e   2$   ��/    �  �K��7Er#���A�%���|,  o�@� `���?�Os93�T0 k� ����T2e   2$   ��/    �  �K��7D�'���A�$&���|,  w�@� `���?�Os:3�T0 k� ����T2e   2$   ��/   �  �K��7D�/���B�,&���|,  �@� `���;�Os;3�T0 k� ����T2e   2$  	 ��/    �  �K��8D�3���C�4&���|,  ��@� `���;�Os<3�T0 k� � �T2e   2$  
 ��/    �  �K��8D�;���D�<&���|,  ��@� `���;�A�=3�T0 k� �	�	T2e   2$   ��/    �  �K��8D�?���E�D'���|,  ��@� `���7�A� >3�T0 k� �$�(T2e   2$   ��/    �  �K��8D�G���E�L'���|,  ��@� `���7�A�$?3�T0 k� �4�8T2e   2$   ��/    �  �K� 8D�K���F�T'���|,  ��@� `���7�A�,@3�T0 k� �H �L T2e   2$   ��/    �  �K�9D�S���G�\'���|,  ��@� `���3�A�0A3�T0 k� �[��_�T2e   2$   ��/    �  �K�9D�W���H�d(���|,  ��@� `� �3�A�4B3�T0 k� �k��o�T2e   2$   ��/    �  �K�9D�_���H�l(���|,  ��@� `��/�A�8C3�T0 k� �����T2e   2$   ��/    �  �K�9D�c���I�t(���|,  Ò@� `��+�A�<D3�T0 k� ������T2e   2$   ��/    �  �K�9D�g���J�x(���|,  ˒@� `�B+�A�@E3�T0 k� ������T2e   2$   ��/    �  �K�$:D�o���J��)���|,  Ӓ@� `�B'�A�DF3�T0 k� ������T2e   2$   ��/    �  �K�(:D�s���K��)���|,  ۑ@� `�B'�A�HG3�T0 k� ������T2e   2$   ��/    �  �K�,:D�w���L��)��|,  �@� `�B#�A�LH3�T0 k� ������T2e   2$   ��/    �  �K�4:D�{���L��)��|,  �@� `�B�A�TI3�T0 k� ������T2e   2$   ��/    �  �K�8:D�����M��*��|,  �@  `�B�A�XJ3�T0 k� ������T2e   2$   ��/    �  �K�<;D�����N��*��!�,  ��@ `�	B�A�\J3�T0 k� ����T2e   2$   ��/    �  �K�@;D�����N��*�'�!�,  �@ `�	B�A�`K3�T0 k� ����T2e   2$   ��/    �  �K�H;D�����O��*�/�!�,  �@ `�
B�A�`L3�T0 k� �+��/�T2e   2$   ��/    �  �K�L;D�����P��*�7�!�,  �@ `�B�A�dM3�T0 k� �;��?�T2e   2$   ��/    �  �K�P;D�����P��+�?�!�,  �@ `�2�A�hN3�T0 k� �K��O�T2e   2$   ��/    �  �K�T;D�����Q��+�G�!�,  �@  `�2 A�lN3�T0 k� �_��c�T2e   2$   ��/    �  �K�X<D�����Q��+�S�!�,  '�@$ `�2 A�pO3�T0 k� �o��s�T2e   2$   ��/    �  �K�`<D�����Q��+�[�!�,  /�@( `�2 A�tP3�T0 k� �����T2e   2$   ��/    �  �K�d<D�����R��+�c�!�,  7�@, `�1�A�xQ3�T0 k� ������T2e   2$   ��/   �  �K�h<D�����R��,�k�!�,  ?�@0 `���A�|Q3�T0 k� ������T2e   2$   (�/    �  �K�l<D�����R��,�s�!�,  G�@4 `���	A�R3�T0 k� ğ����T2e   2$   ��/    �  �K�p<D�����R��,�{�|,  O�@8 `���A�S3�T0 k� ě����T2e   2$   ��/    �  �K�t=D���r�R�,���|,  W�@< `���A�S3�T0 k� ė����T2e   2$   ��/    �  �K�x=D���r�R�,���|,  [�@@ `���A�T3�T0 k� ē����T2e   2$   ��/    �  �K�|=D���r�R�,���|,  c�@D `���A�U3�T0 k� ď����T2e   2$   ��/    �  �K��=D���r�R�-���|,  k�@H `���A�V3�T0 k� ć����T2e   2$   ��/    �  �K��=D���r�R�$-���|,  s�@L `���A�V3�T0 k� ԃ����T2e   2$   ��/    �  �K��=D���2�Q�,-���|,  {�@P `���A�W3�T0 k� �����T2e   2$   ��/    �  �K��=D���2�Q�4-���|,  ��@T `���A�W3�T0 k� �{���T2e   2$   ��/    �  �K��>D���2�Q�<-���|,  ��@X `��A�X3�T0 k� �w��{�T2e   2$   ��/    �  �K��>D���2�Q�D-��|,  ��@\ `��A�Y3�T0 k� �s��w�T2e   2$   ��/    �  �K��>D���2�Q�L.��|,  ��@` `��A�Y3�T0 k� �o��s�T2e   2$   ��/    �  �K��>D���2�Q�P.��!�,  ��@d `��A�Z3�T0 k� �k��o�T2e   2$   ��/    �  �K��>D���2�Q�X.��!�,  ��@d `��!A�Z3�T0 k� �g��k�T2e   2$   ��/    �  �K��>D���2�P�`.��!�,  ��@h `��#A�[3�T0 k� �_��c�T2e   2$   ��/    �  �K��>D���2�P�h.��!�,  ��@l `��$A�\"��T0 k� �W��[�T2e   2$   ��/    �  �K��>D���B�P�p.��!�,  ��@p `��&A�\"��T0 k� �O��S�T2e   2$   ��/    �  �K��?D���B�P�x/��!�,  È@t `��'A�]"��T0 k� �G��K�T2e   2$   ��/    �  �K��?D���B�P��/ �!�,  ˈ@x `��)A�]"��T0 k� �?��C�T2e   2$   ��/    �  �K��?D���B�P��/ �!�,  ӈ@x `��*A�^"��T0 k� �3��7�T2e   2$   ��/    �  �K��?D���B�P��/ �!�,  ۇ@| `��,A�^"��T0 k� �+��/�T2e   2$   ��/    �  �K��?D���B�O��/�!�,  ߇@� `��-A�_"��T0 k� #��'�T2e   2$   ��/    �  �B��?D���B�O��/�!�,  �@� `��/A��_"��T0 k� ���T2e   2$  
 ��/   �  �B��?D��B�O��/'�|,  �@� `��0A��`"��T0 k� ���T2e   2$  	 ��/    �  �B��?D��B�O��0/�|,  ��@� `��2A��`"��T0 k� ���T2e   2$   ��/    �  �B��?D��2�O��07�|,  ��@� `� �3A��a"��T0 k� �����T2e   2$   ��/    �  �B��>D�2�O��0?�|,  �@� `� �4A��a3�T0 k� ����T2e   2$   ��/    �  �E�>D�2�O��0G�|,  �@� `�!�6A��b3�T0 k� ����T2e   2$   ��/    �  �E�>D�2�O��0O�|,  �@� `�!�7A��b3�T0 k� ����T2e   2$   ��/    �  �E�>D�2�O��0W�|,  �@� `�"�8A��c3�T0 k� ��~��~T2e   2$   ��/    �  �E�>D�2�O��0[�|,  #�@� `�"�:A��c3�T0 k� ��}��}T2e   2$   ��/    �  �E�>D�
2�O��0c�|,  '�@� `�#�;A��d3�T0 k� �}��}T2e   2$    ��/    �  �E��>D�2�O��1 k�|,  /�@� `�#�<A��d3�T0 k� �}��}T2e   2$    ,�/    �  �E��>D�2�O��1 s�|,  7�@� `�#�=A��d3�T0 k� �|��|T2e   2$    ��/    �  �E��>D���O��1 {�|,  ?�@� `�$�?A��e3�T0 k� �|��|T2e   2$    ��/    �  �E��>D� ��P��1 ��|,  C�@� `�$�@A��e3�T0 k� �|��|T2e   2$    ��/   �  �E��>D�$��P�1 � |,  K�@� `�%�AA��f3�T0 k� ��|��|T2e   2$    ��/    �  �E��?D�$��P�1 �|,  S�@� `�%�BA��f"s�T0 k� ��|��|T2e   2$    ��/    �  �E��?D�(��P�1 �|,  [�@� `�&�CA��g"s�T0 k� �{|�|T2e   2$    ��/    �  �E� ?D�(��P�1 �|,  _�@� `�&�DA��g"s�T0 k� �o|�s|T2e   2$    ��/    �  �E�?D�,��P�1 �|,  g�@� `�&�EA��g"s�T0 k� �g|�k|T2e   2$    ��/    �  �E�@D�0��P�$1 �|,  o�@� `�'�FA��h"s�T0 k� �_|�c|T2e   2$    ��/    �  �E�@D�0��P�(2 �|,  w�@� `�'�HA��h"s�T0 k� �S|�W|T2e   2$    ��/    �  �E�@D�4 ��P�02�|,  {�@� `�(�IA��h"s�T0 k� �K|�O|T2e   2$    ��/    �  �E�AD�4"��P�42�|,  ��@� `�(�JA��i"s�T0 k� �C|�G|T2e   2$    ��/    �  �E� AD�8$��P�<2�|,  ��@� `�(�KA��i"s�T0 k� �;|�?|T2e   2$    ��/    �  �Es$BD�8&��P�@2�|,  ��@� `�)�LA��j"s�T0 k� �/|�3|T2e   2$    ��/    �  �Es(BD�<'��P�D2��|,  ��@� `�)|MA��j"s�T0 k� �'|�+|T2e   2$    ��/    �  �Es,CD�<)��P�L2��|,  ��@� `�)|NA��j3�T0 k� �|�#|T2e   2$    ��/    �  �Es0CD�@+��P�P2��|,  ��@� `�*xOA��k3�T0 k� �|�|T2e   2$    ��/    �  �Es8DD�@-��P�T2��|,  ��@� `�*xOA��k3�T0 k� �|�|T2e   2$    ��/    �  �Es<ED�D/��P�\2��	|,  ��@� `�*xPA��k3�T0 k� �|�|T2e   2$    ��/    �  �Es@ED�D1��P�`3��
|,  ��@� `�+tQA��l3�T0 k� ��|��|T2e   2$    ��/    �  �EsDFD�H3��P�d3��|,  ��@� `�+tRA��l3�T0 k� ��|��|T2e   2$    ��/    �  �EsHGD�H5��P�l3��|,  ǂ@� `�+pSA��l3�T0 k� ��|��|T2e   2$    ��/    �  �EsLHD�H6��P�p3 �|,  ς@� `�,pTA��l3�T0 k� ��|��|T2e   2$    ��/    �  �EsPID�L8��P�t3|,  Ӄ@� `�,pUA� m3�T0 k� ��|��|T2e   2$    ��/    �  �EsTJD�L:��P�x3|,  ۃ@� `�,lVA� m3�T0 k� ��|��|T2e   2$    ��/    �  �Es\KD�L:��P�|3|,  �@� `�-lVA� m3�T0 k� ��|��|T2e   2$    ��/    �  �Ec`LD�L<��P��3|,  �@� `�-lWA�n3�T0 k� ��|��|T2e   2$    ��/    �  �EcdMLSP=��Q��3� |,  �@� `�-hXA�n3�T0 k� ��|��|T2e   2$    ��/    �  �EchOLSP>��Q��3�(|,  ��@� `�-hYA�n3�T0 k� ��|��|T2e   2$    ��/    �  �EclPLSP@��Q��3�0|,  ��@� `�.hZA�n3�T0 k� ��|��|T2e   2$    ��/    �  �EclQLSTA��Q��3�4|,  �@� `�.dZA�o3�T0 k� ��|��|T2e   2$    ��/    �  �L3pRLSTC��Q��3�<|,  �@� a .d[A�o3�T0 k� ��|��|T2e   2$    ��/   �  �L3tTLSTD��Q��4�D|,  �@� a /d\A�o3�T0 k� ��|��|T2e   2$    ��/    �  �L3xULSXE��Q��4�L|,  �@� a /`]A�p3�T0 k� �|��|T2e   2$    ��/    �  �L3|VLSXF��Q��4�P|,  �@� a /`]A�p3�T0 k� �s|�w|T2e   2$    ��/    �  �L3�WLSXH��Q��4�X|,  '�@� a 0`^A�p3�T0 k� �k|�o|T2e   2$    ��/    �  �L3�YLS\I��Q��4�\|,  +�@�  a 0\_A�p3�T0 k� �c|�g|T2e   2$    ��/    �  �L3�ZLS\J��Q��4�d|,  3�@�  a0\_A�q3�T0 k� �[|�_|T2e   2$    ��/    �  �L3�[LS\K��Q��4�h|,  7�@�  a1\`A�q3�T0 k� �S|�W|T2e   2$    ��/    �  �L3�\LS`M��Q��4�p|,  ?�@�  a1XaA�q3�T0 k� �K|�O|T2e   2$    ��/    �  �L3�]LS`N��Q��4�t|,  G�@�! a1XaA�q3�T0 k� �?|�C|T2e   2$    ��/    �  �L3�^Lc`O��Q��4�||,  K�@�! a2XbA�q3�T0 k� �7|�;|T2e   2$    ��/    �  �L3�_LcdP��Q��4��|,  S�@�! a2XcA�r3�T0 k� �/|�3|T2e   2$    ��/    �  �LC�aLcdQ��Q��4��|,  [�@�! a2TcA�r3�T0 k� �'|�+|T2e   2$    ��/    �  �LC�bLcdR��Q��4��|,  _�@�" a3TdA�r3�T0 k� �|�#|T2e   2$    ��/   �  �LC�cLchS��Q��4��|,  g�@�" a3TeA�r3�T0 k� �|�|T2e   2$    ��/    �  �LC�dLchT��Q��4��|,  k�@�" a3PeA�s3�T0 k� �|�|T2e   2$    ��/    �  �LC�eLchU��Q��5�� |,  s�@�" a3PfA�s3�T0 k� �|�|T2e   2$    ��/    �  �LC�fLchW��Q��5��!|,  {�@�" a4PfA�s3�T0 k� ��|��|T2e   2$    ��/    �  �LC�gLclX��Q��5��!|,  �@�# a4PgA�s3�T0 k� ��|��|T2e   2$    ��/    �  �LC�hLclY��Q��5��"|,  ��@�# a4LgA�s3�T0 k� ��|��|T2e   2$    ��/    �  �LC�iLclZ��Q��5��#|,  ��@�# a4LhA� t3�T0 k� ��|��|T2e   2$    ��/    �  �LC�iLcl[��Q��5��#|,  ��@�# a5LiA� s3�T0 k� ��|��|T2e   2$    ��/    �  �LC�jLcp[��Q��5��$|,  ��@�$ a5LiA� s3�T0 k� ��|��|T2e   2$    ��/    �  �LC�kLcp\��Q��5��$|,  ��@ $ a5LjA� s3�T0 k� ��|��|T2e   2$    ��/    �  �LC�lLcp]��Q��5��%|,  ��@ $ a5HjA� r3�T0 k� ��|��|T2e   2$    ��/    �  �LC�mLct^��Q��6��&|,  ��@ $ a6HkA� r3�T0 k� ��|��|T2e   2$    ��/    �  �LC�nLct_��Q��6��&|,  ��@ $ a6HkA� r3�T0 k� ��|��|T2e   2$    ��/    �  �LC�oLct`��Q��6��'|,  ��@ % a 6HlA� r3�T0 k� ��|��|T2e   2$    ��/    �  �LC�pLcta��Q��6��'|,  ��@% a 6DlA� q3�T0 k� ��|��|T2e   2$    ��/    �  �LC�pLctb��Q��6��(|,  ǌ@% a$6DmA� q3�T0 k� ��|��|T2e   2$    ��/    �  �LC�qLcxc��Q��6��(|,  ˌ@% a$7DmA� q3�T0 k� ��|��|T2e   2$    ��/    �  �LC�rLcxc��R��6��)|,  ӌ@% a(7DnA� q3�T0 k� ��|��|T2e   2$    ��/    �  �LC�sLcxd��R��6��)|,  ۍ@% a(7DnA� p3�T0 k� �|��|T2e   2$    ��/    �  �LC�tLcxe��R��6��*|,  ߍ@& a(7@nA� p3�T0 k� �w|�{|T2e   2$    ��/    �  �LC�uLc|g��R��6��+|,  �@& a08@oA� p3�T0 k� �g|�k|T2e   2$    ��/    �  �LC�vLc|g��R��6��+|,  �@& a08@pA� p3�T0 k� �_|�c|T2e   2$    ��/    �  �LC�wLc|h��R��6��,|,  ��@& a48@pA� o3�T0 k� �W|�[|T2e   2$    ��/    �  �LC�wLc|i��R��6� ,|,  ��@& a88@qA� o3�T0 k� �O|�S|T2e   2$    ��/    �  �LC�xLc�j��R��6�-|,  �@' a88<qA� o3�T0 k� �G�KT2e   2$    ��&    �  �LC�yLc�j��R��6�-|,  �@' a<9<qA� o3�T0 k� �O��S�T2e   2$    ��&    �  �LC�yLc�k��R��6�.|,  �@' a<9<rA� n3�T0 k� �W��[�T2e   2$    ��&    �  �LC�zLc�l��R��6�.|,  �@' a@9<rA� n3�T0 k� �[��_�T2e   2$    ��&    �  �LC�{Lc�m��R��7�/|,  �@' aD9<sA� n3�T0 k� �_��c�T2e   2$    ��&    �  �LC�{Lc�m��R��7�/|,  #�@' aD98sA� n3�T0 k� �g��k�T2e   2$    ��&    �  �LC�|Lc�n��R� 7�0|,  '�@' aH:8sA� n3�T0 k� �k��o�T2e   2$    ��&    �  �LC�}Lc�o��R�7�0|,  +�@' aH:8tA� m3�T0 k� �s��w�T2e   2$    ��&    �  �LC�|Lc�o��R�7� 0|,  3�@' aL:8tA� m3�T0 k� �w��{�T2e   2$    ��&    �  �LC�|Lc�p��R�8�$1|,  7�@' aL:8uA� m3�T0 k� �{���T2e   2$    ��&    �  �LC�|Lc�q��R�8�(1|,  ;�@' aP:8uA� m3�T0 k� ������T2e   2$    ��&    �  �LC�|Lc�q��R�8�(2|,  C�@' aT:8uA� m3�T0 k� ������T2e   2$    ��&    �  �LC�{LS�r��R�8�,2|,  G�@' aX;4vA� m3�T0 k� ������T2e   2$    ��&    �  �LC�{LS�r��R�8�02|,  K�@' aX;4vA� l3�T0 k� ������T2e   2$    ��&    �  �L3�{LS�s��R�8�43|,  S�@' a\;4vA� l3�T0 k� ������T2e   2$    ��&    �  �L3�zLS�t��R�9�43|,  W�@' a`;4wA� l3�T0 k� ������T2e   2$    ��&    �  �L3�zLS�t��R� 9�84|,  [�@' ad;4wA� l3�T0 k� ������T2e   2$    ��&    �  �L3�zLS�u��R�$9�<4|,  _�@' ah<4wA� l3�T0 k� ������T2e   2$    ��&    �  �L3�zEs�u��R�(9�@4|,  c�@' ah<4xA� l3�T0 k� ������T2e   2$    ��&    �  �L3�yEs�v��R�(9�@5|,  g�@' al<0xA� k3�T0 k� ������T2e   2$    ��&   �  �A��yEs�v��R�(9�D5|,  k�@' ap<0xA� k3�T0 k� ������T2e   2$    ��&    �  �A��yEs�v2�R�,9�H6|,  s�@' at<0xA� k3�T0 k� ������T2e   2$    ��&    �  �A��yEs�u2�R�09�L6|,  w�@ ' ax=0yA� k3�T0 k� ������T2e   2$    ��&    �  �A��yA��u2�R�4:�P7|,  {�@ ' a|=0yA� k3�T0 k� ����ÌT2e   2$    ��&    �  �A��yA��u2�R�8:�T7|,  �@ ' a|=0xA� k3�T0 k� �Ì�ǌT2e   2$    ��&    �  �C��xA��u2�R�8:�X8|,  ��@ ' a�=0xA� j3�T0 k� �Ǎ�ˍT2e   2$    ��&    �  �C��xA��t2�R�<:�\9|,  ��@ ' a�>0xA� j3�T0 k� �ˍ�ύT2e   2$    ��&    �  �C��xA��t2�R�@:�`9|,  ��@ ' a�>,xA� j3�T0 k� �ύ�ӍT2e   2$    ��&    �  �C��xAS�t2�R�D:�d:|,  ��@$' a�>,wA� j3�T0 k� �Ӎ�׍T2e   2$    ��&    �  �C��xAS�t2�R�H:�h;|,  ��@$' a�>,wA� j3�T0 k� �׍�ۍT2e   2$    ��&    �  �C��xAS�t2�R�L:l<|,  ��@$' a�>,wA� j3�T0 k� �ۍ�ߍT2e   2$    ��&    �  �ES�xAS�tB�R�P:p<|,  ��@$' a�?,wA� j3�T0 k� �ߎ��T2e   2$    ��&    �  �ES�xAS�tB�R�T:t=|,  ��@$' a�?,vA� j3�T0 k� ����T2e   2$    ��&    �  �ES�xES�tB�R�X:x>|,  ��@$' a�?,vA� i3�T0 k� ����T2e   2$    ��&    �  �ES�xES�sB�R�\:|?|,  ��@(' a�?,vA� i3�T0 k� ����T2e   2$    ��&    �  �ES�wES�sB�R�`:�@|,  ��@(' a�?,vA� i3�T0 k� ����T2e   2$    ��&    �  �EC�wES�sB�R�d:�A|,  ��@(' a�@,vA� i3�T0 k� �����T2e   2$    ��&    �  �EC�wES�sB�R�h;�B|,  ��@(' a�@(uA� i3�T0 k� ������T2e   2$    ��&    �  �EC�wEC�sB�R�l;�C|,  ��@(' a�@(uA� i3�T0 k� ������T2e   2$    ��&    �  �EC�wEC|rB�R�l;�D|,  ��@(' a�@(uA� i3�T0 k� ������T2e   2$    ��&    �  �EC�wEC|r2�R�p;�E|,  ��@(' a�@(uA� i3�T0 k� �����T2e   2$    ��&   �  �C��vECxq2�R�t;�F|,  ��@(' a�@(uA� h3�T0 k� ����T2e   2$    ��&    �  �C��vECxq2�R�x;�G|,  ��@,' a�A(tA� h3�T0 k� ����T2e   2$    ��&    �  �C��vECtq2�R�|;�H|,  Ö@,' a�A(tA� h3�T0 k� ����T2e   2$    ��&    �  �C��uECpp2�R�|;�I|,  ǖ@,( a�A(tA� h3�T0 k� ����T2e   2$    ��&    �  �C��uECpp2�R��;�J|,  ǖ@,( a�A(tA� h3�T0 k� ����T2e   2$    ��&    �  �C��tEClo2�R��;�K|,  ˖@,( a�A(tA� h3�T0 k� ����T2e   2$    ��&    �  �C��tE3hn2�R��;�L|,  ϖ@,( a�B(tA� h3�T0 k� ����T2e   2$    ��&    �  �C��sE3dn2�R��;�L|,  ӗ@,( a�B$sA� h3�T0 k� ����T2e   2$    ��&    �  �C��sE3dm� S��;�L|,  ӗ@,( a�B$sA� h3�T0 k� ����T2e   2$    ��&    �  �C��rE3`l�S��;�L|,  ח@0( a�B$sA� h3�T0 k� ���#�T2e   2$    ��&    �  �C��rE3\l�S��;�M|,  ۗ@0( a�B$sA� g3�T0 k� �#��'�T2e   2$    ��&    �  �C��qE3\k�S��;��M|,  ۗ@0( a�B$sA� g3�T0 k� �#��'�T2e   2$    ��&    �  �C��qCCXj�T��;��N|,  ߗ@0( a�C$sA� g3�T0 k� �'��+�T2e   2$    ��&   �  �C��pCCTi�T��;��N|,  �@0( a�C$rA� g3�T0 k� �+��/�T2e   2$    ��&    �  �C��oCCTh�T��;��N|,  �@0( a�C$rA� g3�T0 k� �+��/�T2e   2$    ��&    �  �C��oCCPh�U��;��N|,  �@0( a�C$rA� g3�T0 k� �/��3�T2e   2$    ��&   �  �C��nCCPg�U��;��N|,  �@0( a�C$rA� g3�T0 k� �3��7�T2e   2$    ��&    �  �K�nCCLf�U��;��O|,  �@0( a�C$rA� g3�T0 k� �3��7�T2e   2$    ��&    �  �K�mCCLf�U��;��O|,  �@4( a�D$rA� g3�T0 k� �7��;�T2e   2$    ��&    �  �K�mCCLe� V��;��P|,  �@4( a�D$rA� g3�T0 k� �7��;�T2e   2$    ��&    �  �K�lCCHe�$V��;��P|,  �@4( a�D$qA� g3�T0 k� �;��?�T2e   2$    ��&    �  �K�lCCHe�$V��;��P|,  ��@4( a�D qA� g3�T0 k� �?��C�T2e   2$    ��&    �  �K�kCCHd�(V��;��P|,  ��@4( a�D qA� f3�T0 k� �?��C�T2e   2$    ��&    �  �K�kCCHd�(V��;��P|,  ��@4( a�D qA� f3�T0 k� �C��G�T2e   2$    ��&    �  �K�kCSHd�(V��;��P|,  ��@4( a�D qA� f3�T0 k� �C��G�T2e   2$    ��&    �  �K�kCSHd3(U��<��P|,  ��@4( a�E qA� f3�T0 k� �G��K�T2e   2$    ��&    �  �K�kCSHd3,U��<��P|,  ��@4( a�E qA� f3�T0 k� �G��K�T2e   2$    ��&   �  �K�kCSHd30U��<��P|,  �@4( a�E pA� f3�T0 k� �K��O�T2e   2$    ��&    �  �                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��� ]�++ � � j}  � �	    � ᝮ     j�� ��    �q           		 Z �          %��    ���  8           d\*         � �δ     d\* �δ           	        	 Z �              ���   0
% 	           O{�     
     �?I     O�� ��    ���   
          D  Z �         �p     ���   0
           <|�   � �
       �d+     <�\ ��    ���              f  Z �           � �  #  ���   8          U�i   � �	    . ���     U�� ŦT    ��             S	 Z �           0�     ���   P
		           H  ��
      B�7�      H�7�                            ���q                ���    P          ��)�        V �I7    �� �x     ��                 �� �         �`     ��H   8            (S        j Q     (S Q*       �                   m �          �     ��@   0
!           J}2         ~ ��     Ja, ��4    �U                 	 �         o�     ��@   H          m
8         � F��     m� F�    �5��                    �         	 i�  �  ��B   (          dpY       �&�     dw�&�    ��                   A �         
 @     ��B   X	
           �J ��     � ��     �J ��                             ���u                ��@                   ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��s�  ��        � �y�    ��h �7�     ��                   x                j  �       �                         ��    ��        � �      ��   �           "                                                �                          � � � � �� � Q � F ��� � �  
   	            
   �   � �� ���L       �� �[� �� \� �� 0\� �D  ]@ �� ]� �D b����J ����X � ˤ _� �� `  � 0_` � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0���� � �� �R� � }`���� � 
�< V� 
�\ W  
�\ W� 
�< W� 
�\ W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���� �  ���3  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"     �j
��   �
� �  �  
� ��    ��     � �       O��  ��     � �      ��    ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �&        �� �T ���        � �+ ��        �        ��        �        ��        �   G�    ����|��        ��                         �$ ( �� ��                                     �                 ����            �� ����%��    � 2                7 Tomas Sandstrom y   4:45                                                                        1  1     �

� �_c�Fwc�VSkj  CC  C$$c~$!	c�4
cV v � s � r �	C.2 �C4* �C73 � C:D �J�8 � J�0 �C+ � C# �J�D � J�< �J�, �J�4 � J�I �c� � �c� � �c� � � c� � �k�> � k�N �	 � � �	!� � �"� � �#� �6$"� q6 %"� �&&� m&'
� | �("�  � )"�2 �*"�  �+*�/6,"� q6 -"� �&.� m& 
� | �  *Oq � *&y u2*y � 3*Oq � *(y � *(y � 6"K � �7"( s � 8"O { p " � � !� p �;!� s* "< s+ "< t, "< u@ "< x                                                                                                                                                                                                                         �� R         �    @ 
             ] P E _  ���� #              	 
�������������������������������������� ���������	�
��������                                                                                          ��    �YE�� ��������������������������������������������������������   �4, ,� @L�@�����V����                                                                                                                                                                                                                                                                                                                                            O� O�                                                                                                                                                                                                                                                \    5    ��  D�J    	  M�  	                           ������������������������������������������������������                                                                                                                                         w     �      �        �        �  �          	  
 	 
 	 	  ��� ��������� � ������ ���� � ������������������� � � ��������������������������� ���������������������� ����������� ��� ���� ��� ������������������ ������������������� �� ��������������� ��������������� ��������������������  ����� � ����            x                      7    ��  R�J   
 T                             �������������������������������������������������������                                                                                                                                        P  5        ��      �       �   �          	 	 
  	 	 	 � ���   � ����������� ������������������������� �  ����������������������������������� ��� �������������������� ����������������������������  ������ ���� ������������������������������� ���������������������� � ������������ �����                                                                                                                                                                                                                                                                                                                               �             


           �   }�                        !                                           '�     'w               ����������������������������  '�   /������������    ������������  '{�������������������������������������ww�ww333wwwwwwww�ww�ww�ww�ww333wwww = E 7               	 
                 � ��� �\         �T�S&+@�IQ+
                                                                                                                                                                                                                                                           
)nY  
                    m      m      d            `      m                                                                                                                                                                                                                                                                                                                                                                                                         @ v  � ��  � ��  � (��  � @��  EZmz  �N :���������������������������������������         :  ���> :�� M        
 	 
�   & AG� �   �              �r�                                                                                                                                                                                                                                                                                                                                     p B J   �     `                 !��                                                                                                                                                                                                                            Y��   �� �� ��      �� B 	      ��� ��������� � ������ ���� � ������������������� � � ��������������������������� ���������������������� ����������� ��� ���� ��� ������������������ ������������������� �� ��������������� ��������������� ��������������������  ����� � ����� ���   � ����������� ������������������������� �  ����������������������������������� ��� �������������������� ����������������������������  ������ ���� ������������������������������� ���������������������� � ������������ �����    ��       ���������������������������������������������������f��ff�fff�ff���������l�ff�ffffl��ff˼fllf������l��̼�ʗ���˹�ffjz�fkyl�l��fƨ�����������������������̼��̉������������������������������f���f�fff�ff�ffl�ff�flfl�l��xl�wwl���l̻�����˺��fl����l�xx��w��̻���l�f�f�ƻ�fl�����ffl�ffffffff���f���̚���ffflffflfffffffffflfffff������������������������l���l������f����������������������������l��lf��f�fff�f��l˪���ww��w�����flflffffffff�̼̙��fww��w��fx�̻�llffff�ffff���fl���f�l�l�˶����fffl��fflfll����ff��ff��lfl�lf��l���l�����������l�������l�������ʼ�j˚��̩��ʨ��ɘ���xxxȈ��ɉ�x���̇�̺������www��ww��xw���x��xk�����������wx��������������x����l�ƈ��Ƈ���w��Ɨ��̩z�̩yf̪�f�������������������������������̙i���ɖ�yɌ��ˌȉ̚ə̩���ə��Ɉ����x�̹x�̹�����������ƺ�������������������ˈ������˙������̫��̺�������˪�������������̸��̗�����̇��̇�����������������������̈���xx����x���w���ɉ��̨���k���̛̻�������������l��Ʀl�Ɗl�l���̻�lk��̺�f̩�l��f�ɫ�ˉ�lɊ�˙���ʚ���˙�˫̼���ɬ�̚��̼�����̼���̬������̼�����˻������������f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff���m�    I      D   "  ��                       B     �   �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �r@  �    � �N ^$   �̞   8  ��  ��   �   �   ��Ҝ     �f ��       p����         �k  �    ��D      �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@     _ 
k ��  _ 
k �$   2\d � ��� �� � ��� �$  v  ��6  �      �       ���� e�����   g���      0 f ^�         �� K             ��`���2�������J����  ��      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                                                �����   �   �   �   ����                                     
�  

  
 � 
 
 
   
   
   
   
  ��                  ��   
   
   
   
   
   
 
 
 � 

  
�                 �   
    �   
    �   
    �   
   
   �  
   �  
   �  
   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    "!  "" "  """ "!    " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "! ""! " ""  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """ "!    " ""  !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         w 
�� ɚ� ���
�˻Ɋ�����������-� �"+ ". "$ "$ �U  Z�  Z�  J�  J�  �D  ��  ��  ɘ ˰ "  �"/�"" "  �  �            g���z��ȩ�����ة�� ���  ̰  ̰  ˰  ��  �  N�� T4�CD  CD0 C40 C30 3;� ܰ �� �� �  �  "  �""�"" �"/���  � �  �      �     �   �   ��  �"" �""  ""   "                 �   ��   �                            � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ��Л�  ��� ��� ������̻��˸��������                    �   P   S                                                                                                                  �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                {`  g`  w                      �  �  ��"� ��� "                               �                        ���� ��� ����                              "  .���"    �     �                                                                                                                                                                                    �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    4U� 4U� 4U� 3UXP�EX��U����  ��                    �  ��� ݼ� �    �    �   �                     �  �  �   �   �   �                   �   �               �  ��� ݼ� w{� �װ vw�      � �������������  �                                �   �                                                                                                  ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                      ��  ��  ���     �     �                                                                                                                                                                                   �ɚ�����˼��˽��̽��˻I���D���DDJ�CEU�4EZ3DJ��D��D�� �� ���  ��  �� "���"��̲
��� ��         @   �   �   ��  ��  ˰  �       �  "�  "   �   "                �                        �  �                      ˢ �+���"����"��"  �   �    �   �" �"� "������     �     �� �� ��
��׊��w٪�|��������            "   "   "       �         �        �   �     �       �   �   �   �   �      �                    ��� ���� �����                                                                                                                                                                                                        �  ��� ��� ��� �ݪ�                       �   �    �z� 
�� ������������ ˍ� ��� ���������ˉ����� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��                    ˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                                         �  ��  �� ��  ��       �  � � �� ��     �      �   �                    ���  ��   �                   � � ����� ��                                                                                                                                                                                    �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   ̻����ߪ����� �                         �  � ��� ��  �   �ˀ ��� ����������+� ""��"�""��"/� ����                                     ��  ��  �                  �  ������� ��             �   �                        �   ��  �   ��   �       �                                                                                                                                  �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �             �  �  �" �.�� "            �   �   �  �  �  �       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��  ��  ���  �   ��  ��  ��  �  �   ��  ��                                                                                                                                                                                       	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                      �   �                           �                        ���� ��� ����                                    � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                                 �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �      �   � � �  ��� ��  �                       �   �                      �������  ���    �                    ��  ��  ���                   ���                                                                                                                                                                          �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                         �   ��   ��                            ����    
�  ��  ��  ��  �����  �   �          ��                           � ��                    ���� �                                                                                                                                                                                                                �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwww""""wwwwwwwGwqGwGwDGwG""""wwwwwwqAqwAwG""""wwwwwwwwDDwwwwwwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwqDDDG""""wwwwwqqADAqq""""wwwwwwqwwwqwqwq""""wwwwqDDDwGq"""$www4ww4Gw4DGw4www4ww4wwwwwwwwwwtwww333DDDGwGGwqwDDwtwwww3333DDDDwGtqGwADqDGwDwwww3333DDDDwwqwwwwDwwDGwwwwww3333DDDDADAGqGqtGwDwwww3333DDDDGqGqGqGqtGwDwwww3333DDDDGqqqwwtDDwwww3333DDDDDDqwqqqwAwtDGwwww3333DDDDwqwqwGqDDGwwwww3333DDDDDGwAwwwwDDtDwwww3333DDDDww4Gw4Gw4Gw4Dww4www43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L����������������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7����������������  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq 

� �_c�Fwc�VSkj !CC C$$c~$"	c�4
cV v � s � r �	C.2 �C4* �C73 � C:D �J�8 � J�0 �C+ � C# �J�D � J�< �J�, �J�4 � J�I �c� � �c� � �c� � � c� � �k�> � k�N �	 � � �	!� � �"� � �#� �6$"� q6 %"� �&&� m&'
� | �("�  � )"�2 �*"�  �+*�/6,"� q6 -"� �&.� m& 
� | �  *Oq � *&y u2*y � 3*Oq � *(y � *(y � 6"K � �7"( s � 8"O { p " � � !� p �;!� s* "< s+ "< t, "< u@ "< x3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������!��9�G�Z��?�K�X�H�K�K�Q� � � � � � � � � �2�0�.�����������������������������������������#��1�K�U�L�L��<�G�T�J�K�X�Y�U�T� � � � � �2�0�.�����������������������������������������"��=�U�S�G�Y��<�G�T�J�Y�Z�X�U�S� � � � � �6�+� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������6�+� � ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                