GST@�                                                            \     �                                               >���      �      b         ���2�������J�������������������        �g     #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    "�j��,  " ��
   �                                                                              ����������������������������������      ��    =b 0Qb 4 114  4c  c  c      	 
      	   
       ��G �� � ( �(                 nn 
)1         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                D   7           @  &   q   �                                                                                 'w w  
)n1n  �    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E 7 �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    R�rBDk�@7� a0 �|3�� L@HDK�<[��MT��8/T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�rBDk�@7� a0 �|3�� M@HDK�<\��MT��8/T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�rBDk�@7� a4 �|3�� M@HDK�@\��Md{��8/T0 k� �E��EU2d  %Q8D"!  ��'    �  R�rBDk�@7� a4 �|3�� N@HDK�@\��Nd{��8/T0 k� �E��EU2d  %Q8D"!  ��'    �  R�rBDk�@7� a4 �|3��N@DDK�D]��Nd{��8/T0 k� �E��EU2d  %Q8D"!  ��'    �  R�rBDk�@7� a8 �|3��N@DDK�H]��Nd{��80T0 k� �E��EU2d  %Q8D"!  ��'   �  R�rBDk�@7� a8 �|3��O@DDK�H^��Nd{��80T0 k� �E��EU2d  %Q8D"!  ��'    �  R�rBDk�@7� a8 �|3��O@DDK�L^��Nd{��80T0 k� �E��EU2d  %Q8D"!  ��'    �  R�rBDk�@7� a< �|3��O@DDK�L_��Nd{��80T0 k� �E��EU2d  %Q8D"!  ��'    �  R�rBDk�@7� a< �|3��P@@DK�P_��Nd{��<0T0 k� �E��EU2d  %Q8D"!  ��'    �  R�rBDk�@7� a< �|3��P@@DK�P_��Odw�4<1T0 k� �E��EU2d  %Q8D"!  ��'    �  R�rBDo�@7� a@ �|3��P@@DK�T`��Odw�4<1T0 k� �E��EU2d  %Q8D"!  ��'    �  R�rBDo�@7� a@ �|3��Q@@DK�T`��Odw�481T0 k� �E��EU2d  %Q8D"!  ��'    �  R�rBDo�@7� a@ �|3��Q@@DK�X`��Otw�481T0 k� �E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aD �|3��Q@@DK�Xa��Otw�482T0 k� �E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aD �|3��R@<DK�\a��Ottd82T0 k� �E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aD �|3��R@<DK�\a��Ottd82T0 k� �E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aD �|3��R@<DK�`b��Pttd82T0 k� �E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aH �|3��R@<DK�`b��Pttd82T0 k� �E��EU2d  %Q8D"!  ��'   �  R�qBDo�@7� aH �|3��S@<DK�db��Ptpd82T0 k� �E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aH �|3��S@<DK�dc��Ptp
d83T0 k� �E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aL �|3��S@8DK�hc��Ptpd83T0 k� �E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aL �|3��T@8DK�hc��Ptpd43T0 k� �E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aL �|3��T@8DK�ld��Ptpd43T0 k� �E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aL �|3��T@8DK�hd��QDpd43T0 k� �|E��EU2d  %Q8D"!  ��'   �  R�qBDo�@7� aP �|3��T@8DK�hd��QDpd43T0 k� �|E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aP �|3��U@8DK�hc��QDpd43T0 k� �|E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aP  |3��U@4DK�hc��QDpd43T0 k� �|E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aT  |3��U@4DK�dc��Q�pd43T0 k� �|E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aT  |3��V@4DK�dc c�Q�ld43T0 k� �|E��EU2d  %Q8D"!  ��'   �  R�qBDo�@7� aT |3��V@4DK�dc c�Q�ld43T0 k� �|E��EU2d  %Q8D"!  ��'    �  R�qBDo�@7� aT |3��V@4DK�dc c�R�l!d43T0 k� �xE�|EU2d  %Q8D"!  ��'    �  R�qBDs�@7� aT |3��V@4DK�dc c�R�l#d43T0 k� �xE�|EU2d  %Q8D"!  ��'    �  R�pBDs�@7� aX |3��W@4DK�`b c�R�l%d03T0 k� �xE�|EU2d  %Q8D"!  ��'    �  R�pBDs�@7� aX |3��W@4DK�`b��R�l&d03T0 k� �xE�|EU2d  %Q8D"!  ��'    �  R�pBDs�@7� aX |3��W@0DK�`b��R�l(d03T0 k� �xE�|EU2d  %Q8D"!  ��'    �  R�pBDs�@7� aX |3��WK�0DK�`b��S�l*d03T0 k� �dD�hDU2d  %Q8D"!  ��'    �  R�pBDs�@7� a\ |3��XK�0D@d`b��S�l,d03T0 k� �TD�XDU2d  %Q8D"!  ��'    �  R�pBDs�@7� a\ |3��XK�0D@d\b��S�l,d03T0 k� �HD�LDU2d  %Q8D"!  ��'    �  R�pBDs�@7� a\ |3��XK�0D@d\b��S�l.d03T0 k� �<D�@DU2d  %Q8D"!  ��'    �  R�pBDs�@7� a\ |3��XK�0D@d\a��S�l/d,3T0 k� �8D�<DU2d  %Q8D"!  ��'    �  R�pBDs�@7� a\ |3��XK�0E@d\a��S�l1d,3T0 k� �4D�8DU2d  %Q8D"!  ��'    �  R�pBDs�@7� a` |3��YK�0E@d\a��S�l3d(3T0 k� �0D�4DU2d  %Q8D"!  ��'    �  R�pBDs�@7� a` |3��YK�0E@�\a��T�p4d(3T0 k� �0D�4DU2d  %Q8D"!  ��'    �  R�pBDs�@7� a` |3��YK�,E@�\`��T�p6d(3T0 k� �,D�0DU2d  %Q8D"!  ��'    �  R�pBDs�@7� a` |3��YK�,E@�\`üT�p7d(3T0 k� �,D�0DU2d  %Q8D"!  ��'    �  R�pBDs�@7� a` |3��YK�,E@�\_üT�p9d$3T0 k� �,D�0DU2d  %Q8D"!  ��'    �  R�pBDs�@7� a` |3��ZK�,E@�\_üT�p:d$3T0 k� �,D�0DU2d  %Q8D"!  ��'    �  R�pBDs�@7� ad |3��ZK�,EE�\^üT�p<d$3T0 k� �(D�,DU2d  %Q8D"!  ��'    �  R�pBDs�@7� ad |3��ZK�,EE�\^üU�p=d 4T0 k� �(D�,DU2d  %Q8D"!  ��'    �  R�pBDs�@7� ad |3��ZK�,EE�\]üU�t?d 4T0 k� �(D�,DU2d  %Q8D"!  ��'    �  R�pBDs�@7� ad |3��ZK�,EE�\]��U�t@d 4T0 k� �(E�,EU2d  %Q8D"!  ��'    �  R�pBDs�@7� ad |3��ZK�,FE�\\��U�tAd4T0 k� �(E�,EU2d  %Q8D"!  ��'    �  R�pBDs�@7� ah |3��[K�,FE�\\��U�tCd4T0 k� �(E�,EU2d  %Q8D"!  ��'    �  R�pBDs�@7� ah |3��[K�(FE�\\��U�tDd4T0 k� �(E�,EU2d  %Q8D"!  ��'    �  R�pBDs�@7� ah |3��[K�(FE�\\��U�tEd4T0 k� �(E�,EU2d  %Q8D"!  ��'    �  R�pBDs�@7� ah |3��[K�(FE�\\��U�tGd4T0 k� �(E�,EU2d  %Q8D"!  ��'    �  R�pBDs�@7� ah |3��[K�(FE�\\��V�tHd4T0 k� �(E�,EU2d  %Q8D"!  ��'    �  R�pBDs�@7� ah |3��[K�(FE�\\��V�xId4T0 k� �(E�,EU2d  %Q8D"!  ��'    �  R�pBDs�@7� ah |3��[K�(FE�\\��V�xJd4T0 k� �$E�(EU2d  %Q8D"!  ��'    �  R�pBDs�@7� al |3��[K�(FE�\[��V�xLd4T0 k� �$E�(EU2d  %Q8D"!  ��'    �  R�pBDw�@7� al |3��[K�(FE�\[��V�xLd5T0 k� �$E�(EU2d  %Q8D"!  ��'    �  R�pBDw�@7� al |3��[K�(FE�\[��V�xL�5T0 k� �$E�(EU2d  %Q8D"!  ��'    �  R�pBDw�@7� al |3��[K�(FE�\[��V�|M�5T0 k� �$E�(EU2d  %Q8D"!  ��'   �  R�pBDw�@7� al |3��[K�(FC�\[��V�|M�4T0 k� �$F�(FU2d  %Q8D"!  ��'    �  R�oBDw�@7� al |3��[K�(GC�\[��W�|M�4T0 k� �$F�(FU2d  %Q8D"!  ��'    �  R�oBDw�@7� al |3��[K�(GC�\[��W�M�4T0 k� �$F�(FU2d  %Q8D"!  ��'    �  R�oBDw�@7� ap |3��[K�$GC�X[��W�Nd4T0 k� �$F�(FU2d  %Q8D"!  ��'    �  R�oBDw�@7� ap  |3��[K�$GC�X[��W�Nd4T0 k� �$F�(FU2d  %Q8D"!  ��'    �  R�oBDw�@7� ap  |3��[K�$GC�X[��W�Od4T0 k� �$F�(FU2d  %Q8D"!  ��'    �  R�oBDw�@7� ap  |3��[K�$GC�X[��W�Od4T0 k� �$F�(FU2d  %Q8D"!  ��'    �  R�oBDw�@7� ap  |3��[K�$GC�X[��W�Pd4T0 k� �$F�(FU2d  %Q8D"!  ��'    �  R�oBDw�@7� ap  |3��[K�$GC�T[��W�Pd4T0 k� �$F�(FU2d  %Q8D"!  ��'    �  R�oBDw�@7� ap  |3��[K�$GC�T\��W�Qd3T0 k� � F�$FU2d  %Q8D"!  ��'    �  R�oBDw�@7� ap  |3��[K�$GC�P\��W�Qd 3T0 k� � F�$FU2d  %Q8D"!  ��'    �  R|oBDw�@7� at  |3��[K�$GC�P\��X�Qd 3T0 k� � F�$FU2d  %Q8D"!  ��'    �  R|oBDw�@7� at $|3��[K�$GC�L\��X�Rd 3T0 k� � F�$FU2d  %Q8D"!  ��'    �  R|oBDw�@7� at $|3��[K�$GC�L\��X�Rc�3T0 k� � F�$FU2d  %Q8D"!  ��'    �  R|oBDw�@7� at $|3��[K�$GC�L\��X�Sc�3T0 k� � F�$FU2d  %Q8D"!  ��'    �  R|oBDw�@7� at $|3� �[K�$GC�L\��X�Sc�3T0 k� � G�$GU2d  %Q8D"!  ��'    �  R|oBDw�@7� at $|3� �[K�$HC�L\��X�Sc�3T0 k� � G�$GU2d  %Q8D"!  ��'    �  R|oBDw�@7� at $|3� �[K�$HC�L\��X�Tc�3T0 k� � G�$GU2d  %Q8D"!  ��'    �  R|oBDw�@7� at $|3� �[K�$HC�H\��X�Tc�3T0 k� � G�$GU2d  %Q8D"!  ��'    �  R|oBDw�@7� at $|3� �[K� HC�H\��X�Tc�3T0 k� � G�$GU2d  %Q8D"!  ��'    �  RxoBDw�@7� ax $|3� �[K� HC�H\��X�Tc�2T0 k� � G�$GU2d  %Q8D"!  ��'    �  RxoBDw�@7� ax (|3� �[K� HC�H\��X�Uc�2T0 k� � G�$GU2d  %Q8D"!  ��'    �  RxoBDw�@7� ax (|3� �[K� HC�H\��X�Uc�2T0 k� � G�$GU2d  %Q8D"!  ��'    �  RxoBDw�@7� ax (|3� �[K� HDH\��Y�Uc�2T0 k� � G�$GU2d  %Q8D"!  ��'    �  RxoBDw�@7� ax (|3� �[K� HDH\��Y�Uc�2T0 k� � G�$GU2d  %Q8D"!  ��'    �  RxoBDw�@7� ax (|3� �[K� HDH\��Y�Uc�2T0 k� � G�$GU2d  %Q8D"!  ��'    �  RxoBDw�@7� ax (|3� �[K� HDH\��YԄUc�2T0 k� � G�$GU2d  %Q8D"!  ��'    �  RxoBDw�@7� ax (|3� �[K� HDH\��YԄUc�2T0 k� �G� GU2d  %Q8D"!  ��'    �  RxoBDw�@7� ax (|3� �[K� HLH\��YԄUc�2T0 k� �G� GU2d  %Q8D"!  ��'    �  RxoBDw�@7� ax (|3� �[K� HLH\��YԄUc�2T0 k� �G� GU2d  %Q8D"!  ��'    �  RxoBDw�@7� a| (|3� �[K� HLH]��YԄUc�2T0 k� �G� GU2d  %Q8D"!  ��'    �  RtoBDw�@7� a| ,|3� �[K� HLH]��YԄUc�2T0 k� �G� GU2d  %Q8D"!  ��'    �  RtoBDw�@7� a| ,|3� �[K� HLH]��Y�Uc�2T0 k� �G� GU2d  %Q8D"!  ��'    �  RtoBDw�@7� a| ,|3�[@ HLH]��Y�Uc�2T0 k� �0H�4HU2d  %Q8D"!  ��'    �  RtoBDw�@7� a| ,|3�[@ HLH]��Y�Uc�2T0 k� �@I�DIU2d  %Q8D"!  ��'    �  RtoBDw�@7� a| ,|3�[@ HLH]��Y�Uc�1T0 k� �LI�PIU2d  %Q8D"!  ��'    �  RtoBDw�@7� a| ,|3�[@ ILH]��Y�Uc�1T0 k� �TJ�XJU2d  %Q8D"!  ��'    �  RtoBDw�@7� a| ,|3�[@ ILH]��Y�Uc�1T0 k� �XJ�\JU2d  %Q8D"!  ��'    �  RtoBD{�@7� a| ,|3�[@ ILH]��YT�Uc�1T0 k� �\J�`JU2d  %Q8D"!  ��'    �  RtoBD{�@7� a| ,|3�[@ IL$H]��YT�Uc�1T0 k� �`J�dJU2d  %Q8D"!  ��'    �  RtoBD{�@7� a| ,|3�[@ IL$H^��YT�Uc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'   �  RtoBD{�@7� a| ,|3�[@ IL$H^��YT�Uc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RtoBD{�@7� a� ,|3�[@ IL$H^��YT�Uc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RtoBD{�@7� a� 0|3�[@IL$H^��YT�Uc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$H_��YT�Uc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$H_��YT|Uc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$H_��YT|Uc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$H_ �Y�|Uc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$H_ �Y�|Uc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$H` �Y�|Uc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$H` �Y�xUc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$H` �Y�xUc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$Ha �Y�xUc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$Da��Y�tUc�1T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$Da��Y�tUc�0T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$Db��Y�pUc�0T0 k� �dJ�hJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 0|3�[@IL$Db��Y�lUc�0T0 k� �`J�dJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 4|3�T[@IL$Db��Y�lUc�0T0 k� �`J�dJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 4|3�T[@IL$Db��Y�lUc�0T0 k� �`J�dJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 4|3�T[@IL$Dc��Y�hUc�0T0 k� �`J�dJU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 4|3�T[@IL$Dc��Y�dUc�0T0 k� �`K�dKU2d  %Q8D"!  ��'    �  RpoBD{�@7� a� 4|3�T[@IL$Dc��Y�`Uc�0T0 k� �`K�dKU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4|3�T[@IL$Dd��Y�\Uc�0T0 k� �`K�dKU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4|3�T[@JL$@d��Y�XUc�0T0 k� �`K�dKU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4|3�T[@JL$@d��Y�TUc�0T0 k� �`K�dKU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4!�3�T[@JL$@e��Y�PUc�0T0 k� �`K�dKU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4!�3�T[@JL$@e��Y�LUc�0T0 k� �`K�dKU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4!�3�T[@JL$@e��Y�LUc�0T0 k� �`K�dKU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4!�3�T[@IL$<f��Y�HUc�0T0 k� �`J�dJU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4!�3��[@IL$<f��Y�HUc�0T0 k� �`J�dJU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4!�3��[@IL$<f��YHUc�0T0 k� �\J�`JU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4!�3��\@IL$<g �YDUc�0T0 k� �\J�`JU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4!�3��\@HL$<g �YDUc�0T0 k� �\I�`IU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4!�3��\@HL$<g �XDUc�0T0 k� �XI�\IU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 4!�3��\@HL$8g �XDUc�0T0 k� �XI�\IU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8!�3��\@HL$8h �XDUc�0T0 k� �XI�\IU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\@GL$8h �XDUc�0T0 k� �XH�\HU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\@GL$8h��XDUc�0T0 k� �TH�XHU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\@GL$8h��XDUc�0T0 k� �TH�XHU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\@GL$8i��XDUc�0T0 k� �TH�XHU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\@GL4i��XTDUc�0T0 k� �PH�THU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\@FL4i��XTDUc�0T0 k� �PG�TGU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\@FL4i��XTDUc�0T0 k� �PG�TGU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\@FL4j��XTDUc�0T0 k� �PG�TGU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\K�FL4j��XTDUc�/T0 k� �8F�<FU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\K�EL4j��X�DUc�/T0 k� �,E�0EU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8|3��\K�EL4j��X�DUc�/T0 k� � D�$DU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8!�3��\K�EL4k��X�DUc�/T0 k� �D�DU2d  %Q8D"!  ��'    �  RloBD{�@7� a� 8!�3��\K�EL4k��X�DTc�/T0 k� �D�DU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� 8!�3��\K�EL4k��X�DTc�/T0 k� �D�DU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� 8!�3��\K�EL4k��X�@Tc�/T0 k� �D�DU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� 8!�3��\K�DL4k��X�@Tc�/T0 k� �C�CU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� 8!�3��\K� DAT4k��X�@Tc�/T0 k� � C�CU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� 8!�3��\K� DAT4k��X�@Tc�/T0 k� ��C� CU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� 8!�3��\K� DAT4k��X�@Tc�/T0 k� ��C� CU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� 8!�3��\K� DAT4k��X�@Tc�/T0 k� ��C� CU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� 8!�3��\K��CAT0k��X�@Tc�/T0 k� ��B� BU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <!�3��\K��CC�0k��X�@Tc�/T0 k� ��B� BU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3��\K��CC�0j��W�@Tc�/T0 k� ��B��BU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3��\K��CC�0j��W�@Tc�/T0 k� ��B��BU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3��\K��CC�0j��W�@Tc�/T0 k� ��B��BU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3��\K��CC�0j��WT@Tc�/T0 k� ��B��BU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3��\K��CC�0j��WT@Tc�/T0 k� ��B��BU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3��\K��BC�0j��WT@Tc�/T0 k� ��A��AU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3��\K��BC�0j��WT@Tc�/T0 k� ��A��AU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3��\K��BC�0j��WT@Tc�/T0 k� ��A��AU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3�T\K��BC�,j��W�@Tc�/T0 k� ��A��AU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3�T\K��BC�,j��W�@Tc�/T0 k� ��A��AU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3�T\K��BC�,j��W�@Tc�/T0 k� ��A��AU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3�T\K��BC�,j��W�@Tc�/T0 k� ��A��AU2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3�T\K��AC�(j��W�@Tc�/T0 k� ��@��@U2d  %Q8D"!  ��'    �  RhoBD{�@7� a� <|3�T\K��AC�(j��W�@Tc�/T0 k� ��@��@U2d  %Q8D"!  ��'    �  ��hB��@.��lӬ]��|+����D��6B����[����3��T0 k� �ϫ�ӫU2d  %Q8D"!  ��" 
   �������gB�#�@.��lӮ]��|+���D��8B����c����3��T0 k� �߫��U2d  %Q8D"!  ��" 
   �������gB�+�@.��lװ]��|+��D��9B����k����3��T0 k� �����U2d  %Q8D"!  ��" 
   �������fB�3�@.��lײ]��|+��E� ;B����s����3��T0 k� �����U2d  %Q8D"!  ��" 
   �������fB�7�@.íl״]��|+��E�<B����w����3��T0 k� ����U2d  %Q8D"!  ��" 
   �������eB�G�E�Ϯl۸헒|+��E�?B���������3��T0 k� ����U2d  %Q8D"!  ��" 
   �������dB�O�E�׮|ۺ헒|+��E�@B���������3��T0 k� ����U2d  %Q8D"!  ��" 
   �������dB�W�E�ۮ|ۼ헒|+�#�E�BB�������Ǆ3��T0 k� ����U2d  %Q8D"!  ��" 
   �������cB�_�E��|߾헒|+�+�E�CB�ð����˄3��T0 k� ����U2d  %Q8D"!  ��" 
   �������cB�g�E��|��헒|+��/�E�$DB�˰����Ӆ3��T0 k� ����U2d  %Q8D"!  ��" 
   �������bB�o�E��|��]��|+��7�B�(FB�ϱ����׆3��T0 k� ����U2d  %Q8D"!  ��" 
   �������bB�w�B^��|��]��|+��;�B�0GB�ױ���߆3��T0 k� ����U2d  %Q8D"!  ��" 
   �������bB��B^��|��]��|+��C�B�4HB�߲����3��T0 k� ����U2d  %Q8D"!  ��" 
   ������ aB΃�B_�|��]��|+��G�B�<JB������3��T0 k� ����U2d  %Q8D"!  ��" 
   ������aB΋�B_�|��]��|+� K�B�@KB������3��T0 k� �#��'�U2d  %Q8D"!  ��"    ������`BΓ�B_�|�����|+� S�B�HLB��з���3��T0 k� �+��/�U2d  %Q8D"!  ��"    ������`BΛ�B_�|�����|+� W�B�LMB���л���3��T0 k� �3��7�U2d  %Q8D"!  ��"    ������ `Bޣ�B_�L�����|/� _�B�TOB���п��3��T0 k� �7��;�U2d  %Q8D"!  ��"    ������(_Bޫ�B_'�L�����|/� c�B�\PB��п��3��T0 k� �?��C�U2d  %Q8D"!  ��"    ������<^B޻�B_3�L�����|/� o�B�hRB���ǳ�3��T0 k� �O��S�U2d  %Q8D"!  ��"    ������D^B�ÆB_;�L�����|/� s�B�pSB���Ǵ�3��T0 k� �S��W�U2d  %Q8D"!  ��"    ������L^B�ˆB_C�	\�����|/� w�B�xTB�'��˶'�3��T0 k� �[��_�U2d  %Q8D"!  ��"    ��� �T]B�φBoK�	\�����|/� �B��UB�/��˷/�3��T0 k� �c��g�U2d  %Q8D"!  ��"    ��� �\]B�ׇBoO�	\�����|3����B��VB�7��ϸ3�3��T0 k� �k��o�U2d  %Q8D"!  ��"    ��� �d]B�߇BoW�	\�����|3����B��XB�?��Ϲ;�3��T0 k� �s��w�U2d  %Q8D"!  ��"    ��� �l\B��Bo_�	\�����|3����B��YB�G��ϺC�3��T0 k� �����U2d  %Q8D"!  �"    ��� �t\B��Bog�	l�����|3����B��ZB�O��ϼG�3��T0 k� ������U2d  %Q8D"! ��/    ��� �|\E��H�k�	l�����|3����B��[B�W��ӽO�3��T0 k� ������U2d  %Q8D"! ��/    ��� Є[E��H�s�	l�����|3����B��\B�_��ӾW�3��T0 k� ������U2d  %Q8D"! ��/    ��� Ќ[E�H�{�	l�����|3����B��]B�g��ӿ_�3��T0 k� ������U2d  %Q8D"! ��/    ��� !И[E�H��	l����|3����B��^B�o����c�3��T0 k� ������U2d  %Q8D"! ��/    ��� &РZE�H��,����|3����B��_B�w����k�3��T0 k� ������U2d  %Q8D"! ��/    ��� +ШZE�H���,���{�|3����B��`B�����.s�3��T0 k� ������U2d  %Q8D"! ��/    ��� 0аZE#�H���,���w�|3����B��`Bއ����.w�3��T0 k� ������U2d  %Q8D"! ��/    ��� 4иYE+�H���,���w�|3����B��aBޏ����.�3��T0 k� ������U2d  %Q8D"! ��/    ��� 8��YE3�H���,���s�|3����B��bBޗ����.��3��T0 k� �����U2d  %Q8D"! ��/    ��� <��YE�;�H���,���o�|3����B��cBޟ����.��3��T0 k� ����U2d  %Q8D"! ��/    ��� @��XE�C�I��,���k�|3����B� dBާ����.��3��T0 k� ����U2d  %Q8D"! ��/    ��� D��XE�K�I��,���g�|3����B�eB������.��3��T0 k� �#��'�U2d  %Q8D"! ��/    ��� H��XE�S�I��,���g�|3����B�fB������.��3��T0 k� �/��3�U2d  %Q8D"! ��/    ��� L��WE�[�I��,���c�|3� ��B�gB���@��.��3��T0 k� �;��?�U2d  %Q8D"! ��/    ��� P��WD�_�I��,���_�|3� ��B�$gB�ǻ@��.��3��T0 k� �K��O�U2d  %Q8D"! ��/    ��� T��WD�g�I�����[�|3� ��B�,hB�ϻ@��.��3��T0 k� �W��[�U2d  %Q8D"! ��/    ��� X� VD�o�I�����W�|3� �B�8iB�׼@�����3��T0 k� �c��g�U2d  %Q8D"! ��/    ��� \�VD�w�I�����S�|3� �B�@jB�߼@���è3��T0 k� �o��s�U2d  %Q8D"! ��/    ��� `�VD��I�����O�|3� �B�HkB��@���ǩ3��T0 k� �{���U2d  %Q8D"! ��/    ��� d�UE���I����O�|3� �B�PkB��@���Ϫ3��T0 k� ������U2d  %Q8D"! ��/    ��� h� UE���I�� �K�|3� �B�\lB���@���ӫ3��T0 k� ������U2d  %Q8D"! ��/    ��� l�(UE���I���G�|3� '�B�dmB���@���۬3��T0 k� ������U2d  %Q8D"! ��/    ��� p�0TE���I���G�|3� /�B�lmB��@����3��T0 k� ������U2d  %Q8D"! ��/    ��� t�8TE���I���C�|3� 3�B�tnB��0����3��T0 k� ������U2d  %Q8D"! ��/    ��� x�@TE���I���C�|3� ;�B݀oB��0����3��T0 k� ������U2d  %Q8D"! ��/    ��� |�HTE���I����?�|3� ?�B݈pB��0����3��T0 k� ������U2d  %Q8D"! ��/    ��� ��PSE���I����;�|3� G�BݐpB�'�0�����3��T0 k� ������U2d  %Q8D"! ��/    ��� ��XSE�ÎI���	�;�|3� K�B��qB�/�0�����3��T0 k� ������U2d  %Q8D"! ��/    ��� ��`SE�ˎI��� �7�|3� S�B��rE�7�0����3��T0 k� ������U2d  %Q8D"! ��/    ��� ��hRB�ӎI���$�7�|3� W�B��rE�?�0���3��T0 k� ��U2d  %Q8D"! ��/    ��� ��pRB�׏I���(�3�|3� _�B��sE�G�0���3��T0 k� ��U2d  %Q8D"! ��/    ��� ��xRB�ߏE���,�3�|3� c�B��tE�O�0���3��T0 k� � �$U2d  %Q8D"! ��/    ��� �рQB��E���0�/�|3� g�E��tE�W�0���3��T0 k� �,�0U2d  %Q8D"! ��/    ��� �шQB��E���4�+�|3� o�E��uE�_� ���3��T0 k� �8�<U2d  %Q8D"! ��/    ��� �ѐQB���E���8�+�|3� s�E��uE�g� ��'�3��T0 k� �D	�H	U2d  %Q8D"! ��/    ��� �јPB���E���<�'�|3� w�E��vD�o� ��+�3��T0 k� �P�TU2d  %Q8D"! ��/    ��� �ѠPB��E��}D�#�|3���E��wD�w� ��3�3��T0 k� �\�`U2d  %Q8D"! ��/    ��� �ѨPB��E�}H��|3����E��wD�� ��;�3��T0 k� �l�pU2d  %Q8D"! ��    ��� ���OB��E#�}L��|3����E� xD߇� ��?�3��T0 k� �x�|U2d  %Q8D"! ��    ��� ���OB��E'�}P��|3����E�xDߏ� ��G�3��T0 k� ����U2d  %Q8D"! ��    ��� ���OB�#�E+�}T��|3����E�yE��� ��O�3� T0 k� ����U2d  %Q8D"! ��    ��� ���NB�+�E3�}X��|3����E�yE��� ��S�3� T0 k� ����U2d  %Q8D"! ��    ��� ���NB�3�E7�}\��|3����E�$zE��� ��[�3� T0 k� ����U2d  %Q8D"! ��    ��� ���MB�;�E�;�}`��|3����E�0zE��� ��c�3� T0 k� ����U2d  %Q8D"! ��    ��� ���MB�C�E�C�}d��|3����E�8{E�����g�3�T0 k� ����U2d  %Q8D"! ��    ��� ���LB�K�E�G�mh��|3����E�@{E������o�3�T0 k� ����U2d  %Q8D"! ��    ��� ���LB�S�E�O�ml��|3����E�L|E������w�3�T0 k� ����U2d  %Q8D"!  ��    ��� ���KB�[�E�S�mp��|3����ET|E������3�T0 k� �� �� U2d  %Q8D"!  -�    ��� ��KB�c�E�W�mt���|3����E\|E�������3�T0 k� ��"��"U2d  %Q8D"!  ��    ��� ��JB�g�E�_�mx���|3����Eh}E�������3�T0 k� �#�#U2d  %Q8D"!  ��    ��� ��IB�o�E�c�mx���|3����Ep}E�������3�T0 k� �%�%U2d  %Q8D"!  ��    ��� ��IB�w�E�k�m|L��|3����E|}E��� ���3�T0 k� �'� 'U2d  %Q8D"! ��    ��� ��$HB��E�s�]�L��|3����E�~F������3�T0 k� �()�,)U2d  %Q8D"! ��    ��� ��,HB���E�w�]�L��|3����E�~F�������3�T0 k� �4*�8*U2d  %Q8D"! ��    ��� ��4GB���E��]�L�|3����B��F�������3�T0 k� �@,�D,U2d  %Q8D"! ��    ��� ��<FB���E���]�L�|3���B��F ������3�T0 k� �P.�T.U2d  %Q8D"! ��    ��� ��DFB���E���]�,�|3���B��F ������3�T0 k� �\0�`0U2d  %Q8D"! ��    ��� ��LEB���B���]�,�|3���B���F ������3�T0 k� �h1�l1U2d  %Q8D"! ��    ��� ��TDB���B���M�,�|3��/�B��F ���
���3�T0 k� �t3�x3U2d  %Q8D"! ��    ��� ��\CB���B���M�,�|3��;�B��D�#������3�T0 k� �|5��5U2d  %Q8D"! ��     ��� �RdCB���B���M�,�|3��G�B��D�+������3�T0 k� ��4��4U2d  %Q8D"! ��     ��� �RlBB�ÕB���M�,�|3��S�B��D�/������3�	T0 k� ��3��3U2d  %Q8D"! ��     ��� �RtAB�˖B���M���|3��_�B��~D�7�������	T0 k� ��2��2U2d  %Q8D"! ��     ��� �R|@B�ӖB��� ����|3��k�B��~D�?�������
T0 k� ��1��1U2d  %Q8D"! ��     ��� �R�@B�ۖB��� ����|3��w�B��~D�G�������
T0 k� ��0��0U2d  %Q8D"! ��     ��� �R�?B��B��� ����|3����B� ~D�O�������
T0 k� ��/��/U2d  %Q8D"! ��     ��� �R�>B��B��� ����|3����B�~D�S������T0 k� ��.��.U2d  %Q8D"! ��     ��� �R�=B��B��� ��,�|3����B�}D�[������T0 k� ��-��-U2d  %Q8D"!  ��     ��� �R�<B���B��� ��,�|3����B�}D�c������T0 k� ��,��,U2d  %Q8D"!  ��     ��� �R�;B���B��� m�,�|3����B�$}D�k������T0 k� ��,��,U2d  %Q8D"!  ��     ��� �R�;B��B��� m�,�|3����B�0}D�s����#��T0 k� ��+��+U2d  %Q8D"!  ��     �   �R�:B��B��� m�,�|3����B�8|D�w����+��T0 k� ��*��*U2d  %Q8D"!  /�     �  �b�9B��B�� m���|3����B�D|D�����3��T0 k� ��)��)U2d  %Q8D"!  ��     �  �b�8B��B�� m���|3����B�L|D�����;��T0 k� ��(��(U2d  %Q8D"!  ��     �  �b�7B�'�B�� m���|3����B�T|D�����C��T0 k� ��'��'U2d  %Q8D"!  ��     �  �b�6B�/�B�� ���|3����B�`|D�����K��T0 k� ��&��&U2d  %Q8D"!  ��     �  �b�5B�7�B�#� ���|3����B�h{D�����S��T0 k� � %�%U2d  %Q8D"!  ��     �  �b�4B�?�B�+� ����|3����B�p{D����[��T0 k� �$�$U2d  %Q8D"!  ��     �  �b�3B�G�B�3� ����|3���B�|{D���� _��T0 k� �#�#U2d  %Q8D"!  ��     �  ���2B�K�B�;� ����|3���Bτ{D����!g��T0 k� �&�&U2d  %Q8D"!  ��     � 	 ��1B�S�B�C�����|3���Bϐ{D����"o��T0 k� � (�$(U2d  %Q8D"!  ��     � 	 ��0B�[�B�K�����|3��#�BϘzD����#�w��T0 k� �()�,)U2d  %Q8D"!  ��     � 	 ��/B�c�B�S�����|3��+�E��zD�����$���T0 k� �0*�4*U2d  %Q8D"!  ��     � 	 ��/B�k�B�_�����|3��7�E��zD�����%����T0 k� �8+�<+U2d  %Q8D"!  ��     � 	 ��$.B�s�B�g�����|3��?�E��yD���� %����T0 k� �@+�D+U2d  %Q8D"!  ��     � 	 ��(-B�{�B�o�����|3��G�E��yD����&����T0 k� �D+�H+U2d  %Q8D"!  ��     � 	 ��0,B���B�w�����|3��O�E��yD����'����T0 k� �L*�P*U2d  %Q8D"!  ��     � 	 ��8+B���B������|3��W�E��xD����(����T0 k� �T)�X)U2d  %Q8D"!  ��     � 	 ��@*B���B�������|3��_�E��xD����)����T0 k� �\(�`(U2d  %Q8D"!  ��     � 	 ��H*B���B������#�|3��g�E��wD���� *����T0 k� �d(�h(U2d  %Q8D"!  ��     � 	 ��P)B���B������'�|3��o�B��wD����(*����T0 k� �l,�p,U2d  %Q8D"!  ��     � 	 ��X(B���Bџ����+�|3��w�B��vD���,+����T0 k� �t.�x.U2d  %Q8D"!  ��     � 	 �d'B���Bѧ����/�|3���B� vD���4,����T0 k� �|/��/U2d  %Q8D"!  ��     � 	 �l'B���Bѯ����7�|3����B�uE��<-����T0 k� ��0��0U2d  %Q8D"!  ��     � 	 �t&B���Bѷ����;�|3���B�uE��D.����T0 k� ��0��0U2d  %Q8D"!  ��     � 	 �|&B�ǚBѿ����?�|3���B�tE��L.����T0 k� ��1��1U2d  %Q8D"!  ��     � 	 ��%B�ϚB������C�|3���B�$sE#��T/����T0 k� ��1��1U2d  %Q8D"!  ��     � 	 ��%B�ךB������K�|3���B�,sE+��X0����T0 k� ��1��1U2d  %Q8D"!  ��     � 	 ��%B�ߚB������O�|3���B�8rF/��`0����T0 k� ��1��1U2d  %Q8D"!  ��     � 	 ��$B��B������[�|3���B�HqF?��p2���T0 k� ��1��1U2d  %Q8D"!  ��     � 	 ��$B��B������c�|3����B�TpFC��x2���T0 k� ��1��1U2d  %Q8D"!  ��     � 	 ��$B���B������g�|3����C \oFK���3���T0 k� ��2��2U2d  %Q8D"!  ��     � 	 ��$B��B�����o�|3����C dnFP �4�#��T0 k� ��4��4U2d  %Q8D"!  ��     � 	 ��$B��B�����s�|3����C lnFT�4�+���T0 k� ��5��5U2d  %Q8D"!  ��     � 	 ��$B��B�����{�|3�2��C xmF\�5�3���T0 k� ��6��6U2d  %Q8D"!  ��     � 	 ��$B��B����̓�|3�2��C �lF`�6�;���T0 k� ��7��7U2d  %Q8D"!  ��     � 	 ��$B�#�B�#���͇�|3�2��E�lFh�6�C���T0 k� ��8��8U2d  %Q8D"!  ��     � 	 ��$B�+�B�+��͏�|3�2��E�kE�p��7�K���T0 k� ��8��8U2d  %Q8D"!  ��     � 	 ��%B�7�B�?��͟�|3�3�E�iE�|��8�[���T0 k� ��8��8U2d  %Q8D"!  ��     � 	  ��%B�?�B�G��ݣ�|3�C�E�iE��	��9�c���T0 k� ��9��9U2d  %Q8D"!  ��     � 	  �%B�G�B�O�� ݫ�|3�C�E�hE��
��9�k���T0 k� ��9��9U2d  %Q8D"!  ��     � 	  �&B�O�B�W��$ݳ�|3�C�E�hI���:�s���T0 k� ��:� :U2d  %Q8D"!  ��     � 	  �&B�W�B�_��,ݻ�|3�C�B��gI���;�{���T0 k� �:�:U2d  %Q8D"!  ��     � 	  �'B�_�B�g��4���|3�C'�B��fI���;����T0 k� �;�;U2d  %Q8D"!  ��     � 	  � (B�g�B�o��<���|3�C+�B��fI���<����T0 k� �;�;U2d  %Q8D"!  ��     � 	  �((B�o�B�w��D���|3�C3�B��eI���=����T0 k� �<�<U2d  %Q8D"!  ��     � 	  �,)B�w�B���L���|3�C7�B��dI!��=����T0 k� � =�$=U2d  %Q8D"!  ��     � 	  �4*B��I���T���|3�C?�B��dI!��>����T0 k� �$>�(>U2d  %Q8D"!  ��     � 	  �@+B���I���d���|3�3K�B�cI!��@����T0 k� �4?�8?U2d  %Q8D"!  ��     � 	  �H,B���I���l���|3�3O�B�bI!��$@����T0 k� �8@�<@U2d  %Q8D"!  ��     � 	  �L-B���I���t��|3�3W�B�bI��,A����T0 k� �@A�DAU2d  %Q8D"!  ��     � 	  �T.B���I���|��|3�3[�B�$aI��4B�����T0 k� �HB�LBU2d  %Q8D"!  ��     � 	  �\/B���I"������|3�3c�B�0`I��<C����T0 k� �LC�PCU2d  %Q8D"!  ��     � 	  �`1B���I"������|3��g�B�8`I��DC����T0 k� �TD�XDU2d  %Q8D"!  ��     � 	  �h2E���I"�����'�|3��o�B�@_I��LD��� T0 k� �XF�\FU2d  %Q8D"!  ��     � 
  �p4E�˝I"�����7�|3��w�B�T^I!��\F��� T0 k� �dH�hHU2d  %Q8D"!  ��     �   �x5E�ϝI�����?�|3���B�\^I!��dG��� T0 k� �lI�pIU2d  %Q8D"!  ��     �   �|7E�םI�����G�|3����B�h]I!��lH���� T0 k� �pK�tKU2d  %Q8D"!  ��     �   Ԅ8E�ߝI�����O�|3����B�p]I!��tH��� T0 k� �tL�xLU2d  %Q8D"!  ��     �   Ԉ9E��I�����W�|3����B�x\I!��|I���T0 k� �|N��NU2d  %Q8D"!  ��     �   �;E��I�����c�|3����B��\E����J���T0 k� ��O��OU2d  %Q8D"!  ��     �   �<E���I"�����k�|3����B��[E����K���T0 k� ��P��PU2d  %Q8D"!  ��     �   �?E��I"�����{�|3����B��ZE����N�'��T0 k� ��T��TU2d  %Q8D"!  ��     �   �AD��I"�������|3����B��ZE����O�/��T0 k� ��U��UU2d  %Q8D"!  ��     �  ��CD��I"�������|3����B��ZE����P�7��T0 k� ��W��WU2d  %Q8D"!  ��     �  ��DD��I�������|3����B��YEq���Q�?��T0 k� ��X��XU2d  %Q8D"!  ��     �  ��FD�#�I�����|3����B��YEq���R�G�"T0 k� ��Z��ZU2d  %Q8D"!  ��     �  ��GD�+�I�����|3����B��XEq���T�K�"T0 k� ��[��[U2d  %Q8D"!  ��  
   �  ��KD�;�I�����|3����B��WEq���V�[�"T0 k� ��^��^U2d  %Q8D"!  ��  
   �  ��LD�C�I#��$ο�|3����B��WD����X�c�"T0 k� �|`��`U2d  %Q8D"!  ��  
   �  ��ND�G�I#��,���|3����B��WD����Y�k�"T0 k� �|a��aU2d  %Q8D"!  ��  
   �  ČOD�O�I#��8���|3����B��VD����Z�s�"T0 k� �xa�|aU2d  %Q8D"!  ��  
   �  ČQD�W�I#��@���|3����B�VD����\�{�"T0 k� �ta�xaU2d  %Q8D"!  ��  
   �  ĈSD�_�I#��H���|3����B�UD����]���"T0 k� �pb�tbU2d  %Q8D"!  ��  
   �  ĈTD�g�I��P���|3����B�UD����_���"T0 k� �pb�tbU2d  %Q8D"!  ��  
   �  ĄWD�s�I��`���|3����B�,TD� ��a���"T0 k� �le�peU2d  %Q8D"!  �  
   �  ĀYD�{�I��h �|3����B�4TF ��c����T0 k� �hf�lfU2d  %Q8D"!  �  
   �  �|[DユI��p �|3���B�@TF��d����T0 k� �dh�hhU2d  %Q8D"!  ��  
   �  �|]E���@#��x �|3���B�HSF��f����T0 k� �dj�hjU2d  %Q8D"!  ��     �  �x^E���@#��� �|3���B�PSF� h����T0 k� �\k�`kU2d  %Q8D"!  ��     �  �pbE���@'��� +�|3���B�dRFsk����T0 k� �Tn�XnU2d  %Q8D"!  ��     �  �ldE���@'� o� 3�|3���B�lRFsl����T0 k� �Lk�PkU2d  %Q8D"!  ��     �  �heE���@+� o� ;�|3���B�xQE�sm����T0 k� �Hj�LjU2d  %Q8D"!  ��     �  �dgE���@+� o� C�|3���B��QE�so����T0 k� �Di�HiU2d  %Q8D"!  ��     �  �\hBC��@/� o� G�|3���B��QE� sp����T0 k� �<i�@iU2d  %Q8D"!  ��     �  �XjBC��@/� o� O�|3���B��PE� �r����T0 k� �8e�<eU2d  %Q8D"!  �     �  �TkBCë@/� o� W�|3�4�B��PE�!�q���"$T0 k� �4a�8aU2d  %Q8D"!  ��    �  �LlBC˫@3� o� _�|3�4�K��PB� !� q���"$T0 k� �0]�4]U2d  %Q8D"!  ��    �  �HnBCϬ@3� o� g�|3�4�K��PB�$"�$q��"$T0 k� �,Z�0ZU2d  %Q8D"! ��    �  �DoBC׬@3� o� k�|3�4�K��OB�("�(p��"$T0 k� �(V�,VU2d  %Q8D"! ��    �  �<pBCۭ@7� o� s�|3�4�K��OB�,#�(p��"$T0 k� �$R�(RU2d  %Q8D"! ��    �  �8rBC�@7� o� {�|3�$�K��OB�0#�,p��"$T0 k� � N�$NU2d  %Q8D"! ��    �  �0rBC�@7� o� �|3�$�K��NB�4$�0o�#�"$T0 k� �J� JU2d  %Q8D"! ��    �  �,sBC�@;� o� ��|3�#��K��NB�8$s4o�+�"$T0 k� �G�GU2d  %Q8D"! ��    �  �$tBC�@;� o� ��|3�#��K��NB�<$s4o�3�"$T0 k� �C�CU2d  %Q8D"! ��    �  � uBC��@;� o� ��|3�#��K��NB�@%s8n�;�"$T0 k� �?�?U2d  %Q8D"! ��    �  �vBC��@?� o� ��|3����K��MB�D%s<n�C�"$T0 k� �;�;U2d  %Q8D"! ��    �  �wBD�@?� o� ��|3����K��MB�L&s@n�K��T0 k� �7�7U2d  %Q8D"! ��    �  �xBD�@?� ` ��|3����K��MB�P&�@n�S��T0 k� �4�4U2d  %Q8D"! ��    �  �yBD�FCC� ` ��|3����K�LB�X'�Dm�c��T0 k� ��,� ,U2d  %Q8D"! ��/    �  � zBD�FCC� ` ��|3����K�LB�`'�Hm�k��T0 k� ��(��(U2d  %Q8D"! ��/    �  ��{BD�FCC� ` ��|3����K�LE�d(�Hm�s��T0 k� ��$��$U2d  %Q8D"! �/    �  ��|BD�FCG� `  ��|3����K� KE�h)�Lm�w��T0 k� ��%��%U2d  %Q8D"! ��/    �  ��|BD#�FCG� `$ ��|3����K�(KE�p)�Lm���T0 k� ��&��&U2d  %Q8D"! ��/    �  ��|BD'�E�K� `( ��|3����K�0KE�t*�LmC���T0 k� ��'��'U2d  %Q8D"! ��/    �  ��}BD3�E�O� `4 ��|3����K�<KE��+�PmC���T0 k� ��)��)U2d  %Q8D"! ��/    �  ��}BD7�E�W� `8 ��|3���K�DJD҄,SPmC���T0 k� ��*��*U2d  %Q8D"! ��/    �  ��}BD;�E�_� `< ��!�3���K�HJDҌ,SPmC���T0 k� ��+��+U2d  %Q8D"!  ��/    �  ��}BD?�B�g� `D ��!�3���K�PJDҐ-SPlC���T0 k� ��,��,U2d  %Q8D"!  ��/    �  ��~BDC�B�o� `H ��!�3���K�TJDҘ.SPlӯ��T0 k� ��-��-U2d  %Q8D"!  ��/    �  ��~BDG�B�w� `L ��!�3���K�\IDҜ/SPlӷ��T0 k� ��.��.U2d  %Q8D"!  ��/    �  �~BDK�B�� `P ��!�3����K�`IDҤ0�Plӻ��T0 k� ��/��/U2d  %Q8D"!  ��/   �  �BDO�B��� `T ��!�3����K�hIDҨ0�Pl����T0 k� ��0��0U2d  %Q8D"!  /�/    �  �~BDW�B��� `\ �!�3����K�tIDҴ2�Tl����T0 k� ��2��2U2d  %Q8D"!  ��/    �  �~BD[�B��� `d �!�3����K�xHDҼ3�Tl����T0 k� ��2��2U2d  %Q8D"!  ��/    �  S�~BD_�B��� `h �!�3����K��HD��4�Tl����T0 k� ��3��3U2d  %Q8D"!  ��/    �  S�}BDc�B��� `l �!�3��� K��HD��5�Tk����T0 k� ��4��4U2d  %Q8D"!  ��/    �  S�}BDg�B��� `p �|3�C�K��HD��6�Tk����T0 k� ��5��5U2d  %Q8D"!  ��/    �  S�}BDk�B��� `t �|3�C�K��HD��7�Tk����T0 k� ��6��6U2d  %Q8D"!  ��/    �  S�}BDo�B��� `x �|3�C�K��GD��8�Tj����T0 k� ��7��7U2d  %Q8D"!  ��/    �  S�|BDs�B��� `| #�|3�C�K��GD��9�Tj����T0 k� ��8��8U2d  %Q8D"!  ��/    �  S�|BDw�B��� `� '�|3�C�K��GD��:�Ti����T0 k� ��9��9U2d  %Q8D"!  ��/    �  S�|BD{�B��� `� /�|3�C�K��GE��<�Th���T0 k� ��;��;U2d  %Q8D"!  ��/    �  S|{BD�B��� `� 3�|3�C�K��GE� =cTh���T0 k� ��<��<U2d  %Q8D"!  ��/    �  Sx{BD��O��� `� 7�|3�C�K��FE�>cTg���T0 k� ��?��?U2d  %Q8D"!  ��'    �  Sp{BD��O��� `� ;�|3�C�K��FE�?cTf���T0 k� ��@��@U2d  %Q8D"!  ��'    �  Sl{BD��O��� `� ?�|3�C�K��FE�@cTe���T0 k� ��A��AU2d  %Q8D"!  ��'    �  Sh{BD��O��� `� C�!�3�C�	K��FE�AcTe�#��T0 k� ��B��BU2d  %Q8D"!  ��'    �  S`zBD��O��� `� K�!�3�S�K��FB�,B�Tc�/��T0 k� ��C��CU2d  %Q8D"!  ��'    �  S\zBD��O�� `� O�!�3�S�K��EB�0C�Tb�3��T0 k� ��C��CU2d  %Q8D"!  ��'    �  S\zBD�O�� `� S�!�3�S�K��EB�8D�Ta�7��T0 k� ��B��BU2d  %Q8D"!  ��'    �  SXzBD�O�� `� W�!�3�S�K��EB�@E�T`�?��T0 k� ��B��BU2d  %Q8D"!  ��'    �  STyBD�O�� `� W�!�3�S�K��EB�HF�T_�C��T0 k� ��B��BU2d  %Q8D"!  ��'    �  SLyBD{�O�� `� _�!�3�S�K��EB�XGT]�O��T0 k� ��B��BU2d  %Q8D"!  ��'    �  SHyBD{�O�� `� c�!�3�S�K��EB�\HT\�S��T0 k� ��B��BU2d  %Q8D"!  ��'    �  SDyBD{�O�� `� g�!�3�S�K��DB�dIT[�W��T0 k� ��A��AU2d  %Q8D"!  ��'    �  S@yBD{�O�� `� k�|3�S�K��DB�lJTZ�[��T0 k� ��A��AU2d  %Q8D"!  ��'    �  S<xBD{�O�� `� k�|3�c�K��DB�tJTX�_��T0 k� ��A��AU2d  %Q8D"!  ��'    �  S8xBDw�O�� `� s�|3�c�K��DB��LTX�k��T0 k� ��A� AU2d  %Q8D"!  ��'    �  S4xBDw�O�� `� w�|3�c�K� DI�MTW�o�� T0 k� � A�AU2d  %Q8D"!  ��'    �  S0xBDw�O�� `� {�|3�c�K�DI�M�XV�s�� T0 k� � A�AU2d  %Q8D"!  ��'    �  S,xBDw�O�� `� {�|3�c�K�DI�N�XU�w��!T0 k� �A�AU2d  %Q8D"!  ��'    �  S(wBDs�O�� `� �|3�c�K�DI�N�\T�{��!T0 k� �A�AU2d  %Q8D"!  ��'    �  S(wBDs�O�� `� ��|3�c�K�DI�O�\T���!T0 k� �A�AU2d  %Q8D"!  ��'    �  S$wBDs�O�� `� ��|3�c�@DI�O�`S���"T0 k� � B�$BU2d  %Q8D"!  ��'    �  S wBDs�O�#� `� ��|3�c�!@DI#�O�dR���"T0 k� �4C�8CU2d  %Q8D"!  ��'    �  SwBDo�O�#� `� ��|3�c�$@DI#�P�hP���#T0 k� �DD�HDU2d  %Q8D"!  ��'    �  SvBDo�@'� `� ��|3�s�&@DI#�P�lO���#T0 k� �PE�TEU2d  %Q8D"!  ��'    �  SvBDo�@'� `� ��|3�s�'@DI#�Q�pO��� $T0 k� �XE�\EU2d  %Q8D"!  ��'    �  SvBDo�@'� `� ��|3�s�)@ DI�Q�tN��� $T0 k� �\E�`EU2d  %Q8D"!  ��'    �  SvBDo�@'� `� ��|3�s�+@ DI�Q�xM��� %T0 k� �dE�hEU2d  %Q8D"!  ��'    �  SvBDo�@+� `� ��|3�s�-@$DI�Q�|L��� %T0 k� �hE�lEU2d  %Q8D"!  ��'    �  SvBDk�@+� `� ��|3�#�.@(DI�Q��K��� %T0 k� �lE�pEU2d  %Q8D"!  ��'    �  SvBDk�@+� `� � |3�#�0@(DI�Q��K���$&T0 k� �pE�tEU2d  %Q8D"!  ��'    �  SvBDk�@/� `� � |3�#�2@,DI#�Q��J���$&T0 k� �pE�tEU2d  %Q8D"!  ��'    �  S uBDk�@/� `� � |3�#�4@,DI#�Q��I���$&T0 k� �tE�xEU2d  %Q8D"!  ��'    �  S uBDk�@/� `� � |3�#�5@0DI#�Q��I���$'T0 k� �xE�|EU2d  %Q8D"!  ��'    �  R�uBDk�@/� `� � |3�#�7@4DI#�Q��H���$'T0 k� �xE�|EU2d  %Q8D"!  ��'    �  R�uBDg�@3� a  � |3�#�9@4DI#�Q��Gԏ��('T0 k� �|E��EU2d  %Q8D"!  ��'    �  R�uBDg�@3� a  � |3�#�;@8DI�Q��Gԏ��((T0 k� �|E��EU2d  %Q8D"!  ��'    �  R�uBDg�@3� a � |3���<@8DI�Q��Hԏ��((T0 k� �E��EU2d  %Q8D"!  ��'    �  R�uBDg�@3� a � |3���=@<DI�Q��Hԏ��((T0 k� �E��EU2d  %Q8D"!  ��'    �  R�uBDg�@7� a � |3���>@<DI�Q��Hԋ��()T0 k� �E��EU2d  %Q8D"!  ��'    �  R�tBDg�@7� a �|3���?@@DI�Q��Hԋ��()T0 k� �E��EU2d  %Q8D"!  ��'    �  R�tBDg�@7� a �|3���@@@DK� Q��ID���,)T0 k� �E��EU2d  %Q8D"!  ��'    �  R�tBDc�@7� a �|3���B@DDK� Q��ID���,*T0 k� �E��EU2d  %Q8D"!  ��'    �  R�tBDg�@7� a �|3���B@DDK�R��ID���,*T0 k� �E��EU2d  %Q8D"!  ��'    �  R�tBDg�@7� a �|3���B@HDK�R��ID���,*T0 k� �E��EU2d  %Q8D"!  ��'    �  R�tBDg�@7� a �|3���C@HDK�S��JD���,*T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�tBDg�@7� a �|3���D@LDK�S��JD���,+T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�tBDg�@7� a �|3���E@LDK�T��JD���0+T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�tBDg�@7� a �|3���E@PDK�T��JD���0+T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�tBDg�@7� a �|3�C�F@PDK�U��KD���0+T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDg�@7� a �|3�C�G@PDK�U��KD���0,T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDg�@7� a  �|3�C�G@TDK�V��KD���0,T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDg�@7� a  �|3�C�H@TDK� V��KD���0,T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDg�@7� a  �|3�C�H@PDK�$W��KT���0-T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDg�@7� a$ �|3�C�I@PDK�$W��LT���4-T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDg�@7� a$ �|3�C�I@PDK�(X��LT���4-T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDg�@7� a( �|3�C�J@PDK�,X��LT���4-T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDk�@7� a( �|3�C�J@LDK�,Y��LT��4-T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDk�@7� a( �|3�C�K@LDK�0Y��LT��4.T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDk�@7� a, �|3���K@LDK�4Z��LT��4.T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDk�@7� a, �|3���L@LDK�4Z��MT��4.T0 k� ��E��EU2d  %Q8D"!  ��'    �  R�sBDk�@7� a0 �|3�� L@HDK�8[��MT��4.T0 k� ��E��EU2d  %Q8D"!  ��'    �                                                                                                                                                                              � � �  �  �  c A�  �J����   �      � \��B� ]�%!%   �� o<�     
	  � �v�     o<� �{      ��                  %          N�     ���   0	          ��s-  $ $       ��@    ��s-�@           
             > �         p     ���   0	%          ����         �R    �����R           
         �� �          `     ���   8	           %    5	      cn'     % cf       y   
            	 A�m          �     ���   8	          '�    9     . O}C     '� Ou      {   
            
   �t           �0     ���   P			         ��p�  ��
      B�)9    ��p��)9           
                ���>              �  ���    P           \L�  � �	   V�9     \rj�=    ���<                $	 Z           �     ��`   H%          A�� � �
     j �Y)     A�h ��#    ���               q  Z           ��    ��h   8�           j#3 : : 	  ~
Y�     jd
��    ���C               ? Z �        /`�    ��@   	@
           W
z  � �
     � �5�     W"� �F�    ���                 Z          	  ���    ��`   H	$
          TT�  > >    ��     TY�R�    ���                Z         
 ��     ��@   H
!
          /�? ��
	      � �B     /�� ��    ���                  ����              F  ��@      0                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          @��  ��        � ��     @�� ���    ���                  x                j  �       �                          @    ��        � �       @   �           "                                                �                          � c O� �
 � ��� � �       
          	
   �   J �� ���F       $ `o� � p�   p� �$ @k� ˤ l` �� l� #� `t� $d u���� ���� ����  ����. ����< ����J ����X � �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0� ���� ����� � 
�| V ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����    ���   ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    "�j�� , " �
� �  �  
�  A    ��     � �      ��    ��     �       A    ��     � �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �'��      ��t1  ���        �:T ���        �        ��        �        ��        �     ��     A����O        ��                         ���   � ����                                     �                 ����             A ����%��     2���2            23/36 (63%) chuk th    4:41                                                                        5  5     �AB�Ia B�Q �
c� � c� � c� �c�0 �c�( �c�@ � 	� �
kj �kp �kt � � �cV: �cZ: �c\" �c_ � cc2 � cd! �k~@ � k�H � k�8 �	� � �	� � �� � �� � �K � �c�. � c�> �J� � � J� � � "� � !"�) �"� �#
�" �$"� � � %"� � �&"� � �'*� � �("� � )"�) �*� �+
�" � ," � �-!� � �." � �/" � �0" � �1!� � �2" � �3* � 4*Hr � 5*Kb � 6)�r �7*z � 8*Or � *(z � :*Qj � ;)�r �<*z � =*Rr � *&z �  )�B                                                                                                                                                                                                                         �� R              @ 
       �     R P E ^  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��    �8)�� ��������������������������������������������������������   �4, 3� * /�� R�� ݃	��@~�	@��9                                                                                                                                                                                                                                                                                                                                ~�M�                                                                                                                                                                                                                                              e  
  2    ��  D�J    	  7�  	                           ������������������������������������������������������                                                                                                                                        �      �      &        �        �  �          	  
 	 
 	 	 ��� ��� ������������������������� �� �������� ������������� ��� ���������������������� �� �������������� � � �� �������� �� ������������ � ������� ���� ������� �����  � � ��� ������������������� ������������������������������� �� ����������            x                      $      �   H�J      *]                             ������������������������������������������������������                                                                                                                                         x       �      �        �    �   �          
 	  
	 
 	 	 ���������������������� ��� ����������������� �� ������������� ������������� �� �  ����������� ������������ �� �������� � ���� ���� �������������������������� ������������  ����������� � ��������������������������� ������������� ������ ����� ���             _                                                                                                                                                                                                                                                                                         
                    �             


           �   }�    �    wwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwww % K ?               	                  � gM(x �\                                                                                                                                                                                                                                                                                      
)n1n  �              e            `                  l                                                                                                                                                                                                                                                                                                                                                                                                              � @� �  � ��  � ��  � 2��  � 2��  � ��  �����F����������������I����������F������������        <  ���B :� u	
        	 �   & AG� �   �   
           � �                                                                                                                                                                                                                                                                                                                                      p B C   �      ��  #             !��                                                                                                                                                                                                                            Y 
 	 �� �� Ѱ�      �� @ 	     ��� ��� ������������������������� �� �������� ������������� ��� ���������������������� �� �������������� � � �� �������� �� ������������ � ������� ���� ������� �����  � � ��� ������������������� ������������������������������� �� �������������������������������� ��� ����������������� �� ������������� ������������� �� �  ����������� ������������ �� �������� � ���� ���� �������������������������� ������������  ����������� � ��������������������������� ������������� ������ ����� ���   �� �     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    A   $   1   �  @                       B     �   �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p����  c@ F �    �      �f ��     �f �$ ^$ �@      ����� ��   �����    ����@ ��   ����@ �$ ^$  /   �        ^ 
j� �� ^ 
j� �$ ^$ � ��� �� � ��� �$ " �  ��"  �      �       b�������2����   g���        f ^�         ��        b      ��C`���2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                                    �����   �   �   �   ����                                     	�  		  	 � 	 	 	   	   	   	   	  ��                  ��   	   	   	   	   	   	 	 	 � 		  	�                 �   	    �   	    �   	    �   	   	   �  	   �  	   �  	   �                                      
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "! ""! " "" """ "!   " ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  ""   "! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "! ""! " "" """ "!   " ""            """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                    ""  ."  �"    �   ��  �   �                  �  �  �  �                                       �  �   ��                     �    � �  ��                  ���                              �   ���                            �   �                                                                                                        �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   �   �"  ""  !� �� ��  �               �   ������  ��                      �   �                      �������  ���    �                             	�                                                                                                                                                                                                  �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �           ��    ��                                 ��            �   �   �   ��                               �� " ��   "                       �    ���  ��                    ��  ��  ��� ���                                                                                                                                                                                                          �   �  �  �  ��  ��  C�  U=  UJ  DZ  D  E  �4 
�: ���+��"��""� """ ""   �   �                        ɪ��ɪw̚�p�������������˻��۽��ݸ�̲-ۻ"""�""�2"�@  �C  �D  �T  D@  �   �   �   "�  "     �� �  �                                        ܰ ˻ �ݚ��w{`  g`  w                      �  �  ��"� ��� "                        "  �"     �                       �������  ���    �                    ��  ��  ���   ���� �                                                                                                                                                                                                                 ��	����ɪ�ܙ����ݼ "-� "� J.��#��C>Z�C U�D �Z�#�U"�C"�� ���                �  �˰ ̻� �wp ׶� �vp �w� ɪ� ��� ��� �ۙ ��� �
� �" 0�" 0.�@ "�            ����˰ + �"  "" "  � �     �  �  ��  �   �           �   �   �   �   ��  ��  ��  ��  ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                            ��  ��  ���   ���� �                                                                                                                                                                                                   �  ��� ��� ��� �ݪ�                       �   �    �z� 
�� ������������ ˍ� ��� ���������ˉ����� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��                    ˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                                         �  ��  �� ��  ���"!�����                            �  �� Ș ��  ��  �      �     �                                      � ����ݼ� ����                                                                                                                                                                    �  ��� ݻ� g�� bm� ggz�'w���������������˛������ˊۼ�����˻������H�DH�@U�DPT�E X�T H�P H�@ Ȥ� ̻� ˘ "�� � ���/�"" �""/���               �   �                                                     �  �                      � �                       ���           �                      �  �  �          ����  �   �             ����                         � "            � "�",�"+� ",                       "  .���"    �     �                              �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                      ��  ��  ���                                      � ���� ��   � � �  �  �   �   �   �                                                                                                                          � �� �������ۛ˽���� �ͼ ��+ �""�B.�R#Z�C U�D �T Z� �; � �� ��� ��  ��� ˽� �wp ��� �vp �w� ��� ˙� ̻� �۰ �ِ ��� Ш� �� >�" 3��.30" ��  �   �                �"/ "" ""  ��  ��                       �  �  ��  �   �   �   �   �   �   ��  ��  ��  ��    ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                     ��  ��  ��� �   ��  ���   �                 ���������������������  ��  ��  ��  �   �    �          �         �                                                                                            ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                      ��� ���� �����                                                                                                                                                                                              � 
��	�˽���w��{k��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            �  �  �  ��  �           �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                      �   �   �      �                                                                            �               �  �  ��  �   �   �       ���                                                                                                                                                                                                    �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��                  �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��           	 
          
        ((((((( 
	(((( ����������������             ! " # $ % & '   ( $ % ) ! " # * ('(&(%($(#("(! (((���������������� + , -   . / 0 1  	 2         3       4 (((((((2	10/(.(-(,(+���������������� 5 6   7   8 9 1 :   $ % ) ! " #   ; ) ! " # $ % ) (#("(!()(%($ :198(((7(6(5����������������    <     = 8 0 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>108(=((( (<���������������� L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L����������������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7����������������  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(�����������������333333333333333333333333333333333333333333333333333333333333����  
�fD
��L���"��������������������D" � j  "  B   J jF� ����
��� �����
���� ����
��� �����
��� 0 q����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqAB�Ia B�Q �
c� � c� � c� �c�0 �c�( �c�@ � 	� �
kj �kp �kt � � �cV: �cZ: �c\" �c_ � cc2 � cd! �k~@ � k�H � k�8 �	� � �	� � �� � �� � �K � �c�. � c�> �J� � � J� � � "� � !"�) �"� �#
�" �$"� � � %"� � �&"� � �'*� � �("� � )"�) �*� �+
�" � ," � �-!� � �." � �/" � �0" � �1!� � �2" � �3* � 4*Hr � 5*Kb � 6)�r �7*z � 8*Or � *(z � :*Qj � ;)�r �<*z � =*Rr � *&z �  )�B3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������#� ��9�K�Z�X��5�R�O�S�G� � � � � � � � � � �/�.�7�������������������������������������������.�G�\�K��7�G�T�Y�U�T� � � � � � � � � �/�.�7�������������������������������������������3�M�U�X��5�X�G�\�I�N�[�Q� � � � � � � �/�.�7�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������/�.�7� �� �������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                