GST@�                                                           �`�                                                      ��     �  H            ���2���$�	 J�����������H�������        �g     	#    ����                                d8<n    �  ?     b`����  �
fD�
�L���"����D"� j   " B   J  jF�"      �j* , . ���
��
�"   "D�j��
� " ��
  �                                                                               ����������������������������������      ��    ??= 000 554 881                  

    

             ��� 44� � ���                 YY� 	         ::�����������������������������������������������������������������������������������������������������������������������������=o  0  4g  1                      �                         �  �  �  �                  E�            8 �����������������������������������������������������������������������������                                ��  -   �  �   @  #   �   �                                                                                '    YY	�  E�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�9O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E * �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    K�|-DXIl�]	\�PE�L���]�A\H&BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�|-DX@��]	\�PD�H#��]�A\H&BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�|-@Y@��]	\�PD�D#��]�A\H&BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K� {-<Y@��]	\�PD�@#��]�A\H&BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�${-<Y@��] ��PD�< #��]�A\H'BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�({-8Z@��] ��PD�< #��]�A\H'BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�,{-8ZA�] ��PD�8!#��]�A\H'BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�0{-4[A�] ��PD�4"#��]�A\H'BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�4{-4[A�] ��PD�0"#��]�A\H'BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�8{-0[A�] ��PD�0##��]�A\H'BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�@{-0\A�] ��PD�,$#��]�A\H'BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�D{-,\A�] ��PD�($#��]�A\H'BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�H{-,]A�] ��PD�(%���]�A\H'BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�Lz-(]A�] ��PD�$&���]�A\H(BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�Pz-(]A�]�PD� '���]�A\H(BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_   � �8E�Tz-$^A�]�PD� (���]�A\H(BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�Xy-$^A�]�PD�)���]�A\H(BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�\y- ^A�]�PD�*���]�A\H(BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�`x _A�]�PD�+���]�A\H(BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�dx_A�]�PD�,���]�A\H(BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�hw_A�]��PD�-���]�A\H(BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�lw`A�]��PD�/���]�A\H(BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�lv`A�]��PD�0���]�A\D(BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�pv`A�]��PD�1#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�tu�aA�]��PD�2#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�xt�aA�]��PD�4#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�xt�aA�]��PD�5#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�|s�aA�]��PD�7#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8E�|s�aA�]��PD� 8#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8C�r�aA�\��PD� 9#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8C�r�aA�\��PD��;#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8C�q�aA�\��PD��<#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8C�p�aK��\��PD��>#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8C�p�aK��\��PD��>#��]�A\D)BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8DS��Ct1C����C��|,	�LA��F ���04E3p^�dT0 k� ����� 2d q&�1D"3Q  ��'    �  ;DS��Sp0C����C��|,	�LA��F ���04E3l^�hT0 k� ����� 2d q&�1D"3Q  ��'    �  9DS��Sp/C����C��|,	�LA��F ���03E3h^�lT0 k� ����� 2d q&�1D"3Q  ��'    �  6DS��Sl-C���ۻC��|,	�HA��F ���03E3d^�tT0 k� ����� 2d q&�1D"3Q  ��'    �  3DS��Sl,C���׺C��|,	�DA��F ���,2E3`^�xT0 k� ����� 2d q&�1D"3Q  ��'    �  0Dc�Sl+C�{��ӹC���|,	�DA��F ���,1E3\^�|T0 k� ����� 2d q&�1D"3Q  ��'    �  -Dcw�Sh*C�w��˸C���|,2@A��E����,0E3\^��T0 k� ����� 2d q&�1D"3Q  ��'    �  *Dcs�Sh)C�o��ǸC��|,2@A!��E����,/E3X^��T0 k� ����� 2d q&�1D"3Q  ��'    �  'Dck�Sh(C�k��D w�|,2<A!��E����(.E3X^��T0 k� �{��� 2d q&�1D"3Q  ��G    �  $Dcc�Sd'C�c��D o�|,2<A!��E����(-E3T^��T0 k� �s��w� 2d q&�1D"3Q  ��G    �  !DcW�S`%C�W��D _�|,24A!��B����(-E#P^��T0 k� �_��c� 2d q&�1D"3Q  ��G    �  DcO�c`$C�S��D W�|,24Eы�B����$,E#L^��T0 k� �[��_� 2d q&�1D"3Q  ��G    �  DcG�c\#C�K���APO�|,20Eу�B���$,E#L^��T0 k� �W��[� 2d q&�1D"3Q  ��G    �  Dc?�c\!C�C���APG�|,2,E�{�B��� +E#L
^��T0 k� �S��W� 2d q&�1D"3Q  ��G    �  Dc;�cX C�?���AP?�|,2(E�s�B��� *E#H^��T0 k� �K��O� 2d q&�1D"3Q  ��G    �  D33�cXC�7���AP;�|,B( E�k�E��� )E#H^��T0 k� �C��G� 2d q&�1D"3Q  ��G    �  D3+�cTC�/���AP3�|,B$ E�c�E���'E#H^��T0 k� �;��?� 2d q&�1D"3Q  ��G    �  D3�cPC�#�w�AP#�|,B�E�O�E���%E#D^��T0 k� �'��+� 2d q&�1D"3Q  ��G    �  	D3�cPC��o�AP�|,B�E�G�E�{��#E#D ^��T0 k� ���#� 2d q&�1D"3Q  ��G    �  D3�cLC��g�AP�|,B�E�?�@�{��"E#G�^��T0 k� ���� 2d q&�1D"3Q  ��G    �  D3�cHC��_�AP�|,B�E�7�@�{��"EG�^��T0 k� ���� 2d q&�1D"3Q  ��G    �   D3�cHC��W�AP�|,B�E�/�@�{��!EG�^��T0 k� ���� 2d q&�1D"3Q  ��G    � ��D2��SDC���O�A_��|,B�E�'�@�{�� EG�^��T0 k� ���� 2d q&�1D"3Q  ��G    � ��D2��SDC���G�A_��|,B�E��@�{�� EK�^��T0 k� ������ 2d q&�1D"3Q  ��G    � ��D2��S@C���?�A_� |,B�E��A {��EK�^��T0 k� ������ 2d q&�1D"3Q  ��G    � ��D2��S<C���3�A_� |,Q��E��A {��EK�^��T0 k� ������ 2d q&�1D"3Q  �G    � ��DB��S<C���+�A_�|,Q��EQ�A {�� EK�^��T0 k� ������ 2d q&�1D"3Q  ��G    � ��DB��8
C����A_�|,Q��EP��A {�� EO�^r�T0 k� ������ 2d q&�1D"3Q  ��G    � ��DB��8	C����A_�|,Q��EP��A {��$ES�^r�T0 k� ������ 2d q&�1D"3Q  ��G    � ��DB��8C���A_�|,Q��EP��AP{��$ES�^r�	T0 k� ����� 2d q&�1D"3Q  ��G    � ��DB��8C����A_�|,Q��EP��AP{��$EW�^r�T0 k� ����� 2d q&�1D"3Q  ��G    � ��DB��4D����A_�|,Q��EP��APw��$E�W�^r�T0 k� ����� 2d q&�1D"3Q  ��G    � ��DB��4D����A_�|,Q��EP��APw��(E�[�^r�T0 k� ����� 2d q&�1D"3Q  ��G    � ��DB��#4D����A_�|,Q��EP��APw��(E�_�^r�T0 k� ����� 2d q&�1D"3Q  ��G    � ��DB��#4 D���ۢA_�|,Q��EP��C�w��(E�c�^r�T0 k� ����� 2d q&�1D"3Q  ��G    � ��DB��#7�D���ӡK�|,a��A`��C�o��(E�c�^r�T0 k� ����� 2d q&�1D"3Q  ��G    � ��DR��#7�D��ˠK�|,a��A`��C�k��(E�g�^r�T0 k� �s��w� 2d q&�1D"3Q  ��G    � ��DR��#;�Dw�ῠK�|,a��A`��C�g��,E�k�^��T0 k� �g��k� 2d q&�1D"3Q  ��G    � ��DR��#;�Do�ᷟK�|,a��A`��C�c��,E�k�^��T0 k� �_��c� 2d q&�1D"3Q  ��G    � ��DR��#;�Dc�ᯟK�|,a��A`��C�_��,E�o�^�� T0 k� �S��W� 2d q&�1D"3Q  ��G    � ��DR{�3;�DS�ᛞE�!�,a��A`��C�S��0
E�s�^���T0 k� �G��K� 2d q&�1D"3Q  ��W    � ��DRs�3?�DK�ᓝE�!�,a��A`��C�O��0E�w�^��T0 k� �/��3� 2d q&�1D"3Q  �W    � ��DRk�3?�DC�ዝE�!�,a��G���C�G��0E�{�^��T0 k� ���� 2d q&�1D"3Q  ��_    � ��DRc�3?�D;��E|!�(a��G���C�C��4E��^��T0 k� ���� 2d q&�1D"3Q ��_    � ��DR_�3C�D3��w�Ex!�(a��G��C�;��4E���^��T0 k� ������ 2d q&�1D"3Q ��_    � ��DRW�3C�D'��o�Et!�(a��G�w�C�7��8Es��`C�T0 k� ������ 2d q&�1D"3Q ��_    � ��DbO�3C�D��g�Ep!�(Q{�G�s�E�/��8Es��`C�T0 k� ������ 2d q&�1D"3Q ��_    � ��DbG�3G�D��_�El!�(Qw�G�o�E�+��<Es��`C�T0 k� ������ 2d q&�1D"3Q ��_    � ��Db7�3G�D��K�Eo`!�(Qg�G�c�E���C�Es��`C�T0 k� ������ 2d q&�1D"3Q ��_    � ��Db3�3K�D���C�Eo\|(Qc�G�_�E���G�Es��`S�T0 k� �w��{� 2d q&�1D"3Q ��_    � ��Db+�3K�D���;�EoX|$Q[�G�[�E���K�Es��`S�T0 k� �c��g� 2d q&�1D"3Q ��_    � ��Db#�3O�C����/�EoT|$QS�G�S�C���K�Es��`S�T0 k� �O��S� 2d q&�1D"3Q ��_    � ��Db�3O�C����'�EoL|$QK�G�O�C����O�Ec��`S�T0 k� �;��?� 2d q&�1D"3Q ��_    � ��Db�3O�C����EoH	|$QG�G�K�C����S�Ec��`S�T0 k� �'��+� 2d q&�1D"3Q ��_    � �|Db�3S�C����EoD	|$�?�G�G�C����W�Ec��`S�T0 k� ���� 2d q&�1D"3Q ��_    � �wDb�3S�C����Eo<
|$�7�G�C�C����[�Ec��`S�T0 k� ����� 2d q&�1D"3Q ��_    � �sD1��3S�C����Eo8
|$�/�G�?�P����_�Ec��`S�T0 k� ������ 2d q&�1D"3Q ��_    � �oD1��3W�C�� ��Eo4|$�+�G�;�P����_�D3��`c�T0 k� ������ 2d q&�1D"3Q ��_    � �kD1��3W�C�� �Eo,|$�#�G�3�P����c�D3��`c#�T0 k� ������ 2d q&�1D"3Q ��_    � �gD1��3W�C�� �E_(| ��G�/�P����g�D3��`c'�T0 k� ������ 2d q&�1D"3Q ��_    � �dD1��3[�C�� ߔE_ !� ��G�+�P����k�D3��`c+�T0 k� ������ 2d q&�1D"3Q ��_    � �aD1��3[�C��PӔE_!� ��G�'�P����k�D3��`c+�T0 k� ������ 2d q&�1D"3Q ��_    � �^D1��3[�C��P˓E_!� ��G�#�P����k�D3��`c/�T0 k� �o��s� 2d q&�1D"3Q ��_    � �[D1��3[�C��PÓE_!� ���G��P����o�D3��`c3�T0 k� �[��_� 2d q&�1D"3Q ��_    � �XD1��3[�C��P��E_!� ���G��P����s�D3��`c7�T0 k� �G��K� 2d q&�1D"3Q ��_    � �VD1��3_�C�s�P��E_!� ���G��P����w�D3��`c?�T0 k� �3��7� 2d q&�1D"3Q ��_    � �TD1��3_�C�k�P��E^�!� ���G��P����{�D3��`cC�T0 k� ���� 2d q&�1D"3Q ��_    � �RD1��3_�C�c�P��E^�!� ���G��P����{�D3��`cG�T0 k� ���� 2d q&�1D"3Q ��_    � �PDA��3_�C�[�P��E^�!� ���G��P�����DC��`cK�T0 k� ������ 2d q&�1D"3Q ��_    � �NDA��3_�C�S�P��EN�!� ���G��P���s�DC��`cK�T0 k� ������ 2d q&�1D"3Q ��_    � �LDA��3c�C�K�P��EN�!� �ǿG��P���s�DC��`cK�T0 k� ������ 2d q&�1D"3Q ��_    � �JDA��3c�C�C�@w�EN�| �G��P��s�DC��Z�K�T0 k� ������ 2d q&�1D"3Q ��_    � �HDA��3c�C�7�@o�EN�| �G���P�{�s�DC��Z�K�T0 k� ������ 2d q&�1D"3Q ��_    � �GDA��3c�C�/�@g�EN�| �C���P�s�s�DC��Z�K�T0 k� ������ 2d q&�1D"3Q ��_    � �FDA�3c�D'�@_�E��| �C���P�o�s��DC��Z�K�T0 k� �w��{� 2d q&�1D"3Q ��_    � �EDAw�3g�D�@S�E޼| �C���C�g�s��DC��Z�K�T0 k� �c��g� 2d q&�1D"3Q ��_    � �DDAo�3g�D�@K�E޴| �C���C�c�s��DC��Z�K�T0 k� �O��S� 2d q&�1D"3Q ��_    � �CDAg�3g�D�@C�Eެ|  ��C���C�[�s��DC��Z�K�T0 k� �;��?� 2d q&�1D"3Q  ��_    � �BDAc�3g�D�@7�Eޤ|  ��C���C�W�s��DC��Z�K�T0 k� �'��+� 2d q&�1D"3Q  ��_    � �ADQ[�3g�D ��@/�Eޜ|  ��C���C�O�c��DS��Z�K�T0 k� ���� 2d q&�1D"3Q  .�_    � �@DQS�3g�D ��@'�Eޔ|  {�C���C�G�c��DS��`3K�T0 k� ����� 2d q&�1D"3Q  ��_    � �?DQK�3g�D ����C��  s�C���C�C�c��DS��`3K�T0 k� ������ 2d q&�1D"3Q  ��_    � �>DQC�3g�D ����C��  k�C���C�;�c��DS��`3O�T0 k� ������ 2d q&�1D"3Q  ��_    � �=DQ?�3g�D ����C�|�  c�C���C�3�c��DS��`3O�T0 k� ������ 2d q&�1D"3Q  ��_    � �<DQ7�3g�D �����C�t�  [�C���C�/�	���Ec��`3O�T0 k� ������ 2d q&�1D"3Q  ��_    � �;DQ/�3g�D�����C�l�  S�C���C�'�	���Ec��Z�S�T0 k� ������ 2d q&�1D"3Q ��_    � �:DQ'�3g�D����C�d�  K�C���A_�	���Ec��Z�S�T0 k� ������ 2d q&�1D"3Q ��_    � �9DQ�3g�D����C�\�  C�C���A_�	���Ec��Z�W�T0 k� �o��s� 2d q&�1D"3Q ��_    � �8DQ�3g�D���ےC�T� ;�C���A_�	���Ec��Z�W�T0 k� �[��_� 2d q&�1D"3Q ��_    � �8DQ�3g�D���ӒC�L� 3�C���A_�	Ã�Ec��Z�[�T0 k� �G��K� 2d q&�1D"3Q �_    � �8Da�3g�D���ǓC�D� +�C���A_�	Ã�ES��Z�_�T0 k� ,K��O� 2d q&�1D"3Q ��_    � �8Da�3g�D�����C�8� #�C���A^��	Ã�ES��Z�c�T0 k� ,K��O� 2d q&�1D"3Q ��_    � �8D`��3g�D�����C�0� �C���A^��	Ã�ES��Z�c�T0 k� ,K��O� 2d q&�1D"3Q ��_    � �8D`��3g�D�����C�(� �C���A^��	Ã�ES��Z�g�T0 k� ,K��O� 2d q&�1D"3Q ��_    � �8D`��3g�D{����C� � �C���A^��	���ES��Z�k�T0 k� ,K��O� 2d q&�1D"3Q ��_    � �8D`��3k�Ds����C�� ��C�{�A^��	���C���Z�o�T0 k� ,K��O� 2d q&�1D"3Q ��_    � �8D`��3k�C�k����C�� ��Dw�A^��	���C���Z�w�T0 k� �O��S� 2d q&�1D"3Q ��_    � �8D`��3k�C�c����C�� �Do�A^��	���C��Z�{�T0 k� �O��S� 2d q&�1D"3Q ��_    � �8D`��3k�C�[���C� � �Dg�A^��	���C��Z��T0 k� �O��S� 2d q&�1D"3Q ��_    � �8D`��3k�C�O��w�C��� �ߩD_�A^��	Ã�C��ZÃ�T0 k� �O��S� 2d q&�1D"3Q ��_    � �8D`��3k�C�G��o�C��� �רDW�A^��	Ã�C��ZÇ�T0 k� �O��S� 2d q&�1D"3Q	 ��_    � �8D0��3k�C�?��g�EM�� �ϨDO�A^��	Ã�C��ZË�T0 k� <O��S� 2d q&�1D"3Q	 ��_    � �8D0��3k�C�7��[�EM�� �ǧDG�A^��	Ã�C��ZÏ�T0 k� <O��S� 2d q&�1D"3Q
 ��_    � �8D0��3k�C�/��S�EM�� ￧D;�A^��	Ã�C��ZÓ�T0 k� <S��W� 2d q&�1D"3Q
 ��_    � �8D0��3k�C�'��K�EM�� ﷦D3�A^��	���C��Z×�T0 k� <S��W� 2d q&�1D"3Q ��_    � �8D0��3k�C���C�EM�� ﯦD+�A^��	���C��Z×�T0 k� <S��W� 2d q&�1D"3Q ��_    � �8D0��3k�C���;�EM�� 痢D#�A^��	���C��ZÛ�T0 k� �S��W� 2d q&�1D"3Q ��_    � �8D0��3k�C���/�EM�� D�A^��	���C��Zß�T0 k� �S��W� 2d q&�1D"3Q ��_    � �8D0��3k�C���'�EM�� D�A^��	���C��Zã�T0 k� �S��W� 2d q&�1D"3Q ��_    � �8D0��3k�C�����EM�� D�A^��	Ã�C��Zç�T0 k� �W��[� 2d q&�1D"3Q ��_    � �8D0�3k�C�����EM�� D��A^��	Ã�C��Zë�T0 k� �W��[� 2d q&�1D"3Q ��_    � �8D0w�3k�C�����C��� �{�D��A^��	Ã�E��Zï�T0 k� ,W��[� 2d q&�1D"3Q ��_    � �8D0o�3k�C�����C��� �s�D��A^��	Ã�E��Zï�T0 k� ,W��[� 2d q&�1D"3Q ��_    � �8D@g�3k�C������C�|� �k�D��A^��	Ã�E��Zó�T0 k� ,W��[� 2d q&�1D"3Q ��_    � �8D@_�3k�C�����C�t� �c�D��A^����E��Z÷�T0 k� ,W��[� 2d q&�1D"3Q ��_    � �8D@[�3k�C�����C�l� �[�D��A^{����E��Z÷�T0 k� ,W��[� 2d q&�1D"3Q ��_    � �8D@S�3k�C�����C�d� �S�D��A^w����E��Zû�T0 k� �[��_� 2d q&�1D"3Q ��_    � �8D@K�3k�C����ۥC�\� �K�D��A^s����E��Zû�T0 k� �[��_� 2d q&�1D"3Q ��_    � �8D@C�3k�C����ϦC�T� �?�C��A^o����D3��Zÿ�T0 k� �[��_� 2d q&�1D"3Q ��_    � �8D@?�3k�D���ǧC�L� �7�C��A^k�S��D3��Zÿ�T0 k� �[��_� 2d q&�1D"3Q ��_    � �8D@7�3k�D��ο�C�@� �/�C��A^g�S��D3��Z���T0 k� �[��_� 2d q&�1D"3Q ��_    � �8D@/�3k�D��η�EM8� �'�C��A^_�S��D3�Z���T0 k� L[��_� 2d q&�1D"3Q ��_    � �8D@'�3k�D��ί�EM0� �C��A^[�S��D3w�Z���T0 k� L_��c� 2d q&�1D"3Q ��_    � �8D@#�3k�D��Χ�EM(� �C��A^W�S��ESs�Z���T0 k� L_��c� 2d q&�1D"3Q ��_    � �8DP�3o�D{�Ο�EM � �C��A^W�S��ESo�Z���T0 k� L_��c� 2d q&�1D"3Q �_    � �8DP�3o�E�s�N��EM� �A^�A^S�S��ESk�Z���T0 k� L_��c� 2d q&�1D"3Q �_    � �8DP�3o�E�g�N��E�� ��A^w�A^O�S��ESg�Z���T0 k� �_��c� 2d q&�1D"3Q ��_    � �8DP�3o�E�_�N��E�� ^��A^o�A^K�S��ESc�Z���T0 k� �_��c� 2d q&�1D"3Q ��_    � �8D_��3o�E�W�N{�E� � ^�A^g�C�G�S��ES_�Z���T0 k� �_��c� 2d q&�1D"3Q ��_    � �8D_��3o�E�O�Ns�E��� ^�A^_�C�C�S��ES[�Z���T0 k� �c��g� 2d q&�1D"3Q ��_    � �8D_��3o�E�G�Nk�E��� ^ߚA^W�C�?�S��ASW�Z���T0 k� �c��g� 2d q&�1D"3Q ��_    � �8D_��3o�E�?�Nc�E��� ^ךA^O�C�7�S��ASS�Z���T0 k� ,c��g� 2d q&�1D"3Q ��_    � �8D_��3o�E�7�N[�E��� ^ϚA^G�C�3�S��ASO�Z���T0 k� ,c��g� 2d q&�1D"3Q ��_    � �8D_��3o�E�+�NS�E��� ^ǙA^?�E^/�S��ASK�Z���T0 k� ,c��g� 2d q&�1D"3Q ��_    � �8D_��3o�E�#�>K�E��� ^ÙA^7�E^+�S��ASG�Z���T0 k� ,c��g� 2d q&�1D"3Q ��_    � �8Do��3o�E��>C�E��� ^��A^3�E^'�S��ASC�Z���T0 k� ,g��k� 2d q&�1D"3Q ��_    � �8Do��3o�E��>;�Eܼ� ^��A^+�E^�S��AS?�Z���T0 k� �g��k� 2d q&�1D"3Q ��_    � �8Do��3o�D?�>3�Eܴ� ^��A^#�E^�S��AS;�Z���T0 k� �g��k� 2d q&�1D"3Q ��_    � �8Do��3o�D?�>+�Eܬ� ^��A^�EN�S��AS7�Z���T0 k� �g��k� 2d q&�1D"3Q ��_    � �8Do��Co�D>��N'�E�� ^��A^�EN�S��AS3�Z���T0 k� �g��k� 2d q&�1D"3Q ��_    � �8Do��Co�D>��N�E�� ^��A^�EN�S��AS/�Z���T0 k� �g��k� 2d q&�1D"3Q
 ��_    � �8Do��Co�D>��N�E�� ^��A^�EN�S��AS/�Z���T0 k� <g��k� 2d q&�1D"3Q
 ��_    � �8Do��Co�D>��N�E�� ^��A^�EM��S��AS+�Z���T0 k� <k��o� 2d q&�1D"3Q	 ��_    � �8Do��Co�D>��N�E�� ^��A]��P}��S��AS'�Z���T0 k� <k��o� 2d q&�1D"3Q	 ��_    � �8Do� Co�D>��N�E�x� ^�A]��P}��S��AS#�Z���T0 k� <k��o� 2d q&�1D"3Q ��_    � �8Do� Co�D>��M��E�p� ^{�A]��P}��S��AS�Z���T0 k� <k��o� 2d q&�1D"3Q ��_    � �8D?|Co�D>��M��E�h� ^s�A]��P}��S��AS�Z���T0 k� �k��o� 2d q&�1D"3Q ��_    � �8D?tCo�DN��]��E�`� ^o�A]��P}��S��AS�Z���T0 k� �k��o� 2d q&�1D"3Q ��_    � �8D?pSo�DN��]��E�T� ^g�A]��P���S��AS�Z���T0 k� �o��s� 2d q&�1D"3Q ��_    � �8D?hSo�DN��]��E�L� ^c�A]��P���S��AS�Z���T0 k� �o��s� 2d q&�1D"3Q �_    � �8D?`So�DN��]��E�D� ^_�A]��P���S��AS�Z���T0 k� �o��s� 2d q&�1D"3Q ��_    � �8D?XSo�DN��]��E�D�  ^W�A]��P���S��AS�Z���T0 k� ,o��s� 2d q&�1D"3Q ��_    � �8D?TSo�DN�����E�<�#�^S�A]��P���S��AS�Z���T0 k� ,o��s� 2d q&�1D"3Q ��_    � �8D?LSo�DN�����E�4�#�^O�A]��P���S��AS�Z���T0 k� ,o��s� 2d q&�1D"3Q ��_    � �8D?DSo�DN{����E�,�#�^G�A]��P���S��AS�Z���T0 k� ,s��w� 2d q&�1D"3Q ��_    � �8D?<So�DNs����E�(�#�^C�A]��P���S��AS�Z���T0 k� ,s��w� 2d q&�1D"3Q  ��_    � �8D?8So�DNk����E� �#�^?�A]��P}��S��AR��Z���T0 k� �s��w� 2d q&�1D"3Q  ,�_    � �8D?0�o�DNc����E��#�^7�A]��P}��S��AR��Z���T0 k� �s��w� 2d q&�1D"3Q  ��_    � �8DO(�o�D^[����E��#�^3�A]��P}��S��AR��Z���T0 k� �s��w� 2d q&�1D"3Q  ��_   � �8DO$�o�D^S����E��#�^/�A]��P}��S��AR��Z���T0 k� �s��w� 2d q&�1D"3Q ��_   � �8DO	�o�D^K����E��'�^+�A]��P}��S��AR��Z���T0 k� �s��w� 2d q&�1D"3Q ��_    � �8DO	�o�D^C����F��'�^'�A]� C���S��AR��Z���T0 k� Lw��{� 2d q&�1D"3Q ��_    � �8DO
�k�D^;����F��'�^�A]� C���S��AR��Z���T0 k� Lw��{� 2d q&�1D"3Q ��_    � �8DO
�k�D^3����F��+�^�A]� C���S��AR��Z���T0 k� Lw��{� 2d q&�1D"3Q ��_    � �8DO �g�D^+����F��+�^�A]� C���S��AR��Z���T0 k� Lw��{� 2d q&�1D"3Q ��_    � �8DN��g�D^#����F��/�^�A]� C���S��AR��Z���T0 k� Lw��{� 2d q&�1D"3Q ��_    � �8DN��g�D^ ���D���/�^�A]| C���S��AR��Z���T0 k� �w��{� 2d q&�1D"3Q ��_    � �8DN��c�D^���D���3�^�A]x C���S��AR��Z���T0 k� �{��� 2d q&�1D"3Q ��_    � �8DN��_�D^���D���7�^�A]t C���S��AR��Z���T0 k� �{��� 2d q&�1D"3Q ��_    � �8D^�S_�Dn ���D���7�^�A]p C�{�S��AR��Z���T0 k� �{��� 2d q&�1D"3Q ��_    � �8D^�S[�Dm����D���;�]��A]l C�w�S��AR��Z���T0 k� �{��� 2d q&�1D"3Q ��_    � �8D^�SW�Dm����D���?�]��A]h C�s�S��AR��Z���T0 k� ,{��� 2d q&�1D"3Q ��_    � �8D^�SS�Dm����D���C�]��A]d C�k�S��AR��Z���T0 k� ,{��� 2d q&�1D"3Q ��_    � �8D^�SS�Dm���D���G�]�A]` C�g�S��AR� Z���T0 k� ,{��� 2d q&�1D"3Q ��_    � �8D^�SO�Dm��{�D�� �K�]�A]\ C�c�S��AR� Z���T0 k� ,���� 2d q&�1D"3Q ��_    � �8D^�CK�Dm��w�Dۼ"�O�]�A]X C�[�S��AR� Z���T0 k� ,���� 2d q&�1D"3Q ��_    � �8L>�CG�Dm��s�D۸#�S�]�A]T C�W�S��AR� Z���T0 k� ����� 2d q&�1D"3Q ��_    � �8L>�CC�L=�	�o�D�$�W�]�A]P C�O�S��AR� Z���T0 k� ����� 2d q&�1D"3Q ��_    � �8L>�C?�L=�
�o�D�%!\[�]ߎA]L C�K�S��AR�Z���T0 k� ����� 2d q&�1D"3Q ��_    � �8L>�C;�L=��k�D�&!\_�]ߎA]H C�C�S��AR�Z���T0 k� ����� 2d q&�1D"3Q ��_    � �8L>��7�L=��g�D�'!\c�]ێA]D C�;�S��AR�Z���T0 k� ������ 2d q&�1D"3Q ��_    � �8L>��3�L=��c�D�)!\g�]׎A]@ C�7�S��AR�Z���T0 k� <����� 2d q&�1D"3Q ��_    � �8L>��/�L=��_�D�*!\k�]ӍA]@ C�/�S��AR�Z���T0 k� <����� 2d q&�1D"3Q ��_    � �8L>|�+�L=��_�L{�+!\o�]ύA]< C�+�S��AR�Z���T0 k� <����� 2d q&�1D"3Q ��_    � �8L>t�#�L=��[�L{�,!\o�]ˍA]8 C�#�S��AR�Z���T0 k� <����� 2d q&�1D"3Q ��_    � �8L>p��L=��W�L{�-!ls�]ˍA]4 C��S��AR�Z���T0 k� <����� 2d q&�1D"3Q ��_    � �8L>h��L=��S�L{�/!lw�]ǍA]0 C��S��AR�Z���T0 k� ������ 2d q&�1D"3Q ��_    � �8L>`��L=x�O�L{�0!l{�]ÍA],C��S��AR�Z���T0 k� ������ 2d q&�1D"3Q  $�_    � �8L>X��L=t�K�L{�1!l�]��A],C��S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��_    � �8L>T��L=l�K�L{�2!l��]��A](C���S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��_    � �8LNL��L=h�G�L{�3!l��]��A]$C���S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��_    � �8LND��LM`�C�L{�4!l��]��A] C���S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��_    � �8LN@���LM\�?�L{�5!l��]��A] C���S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��_    � �8LN8���LMT�?�L{�6!l��]��A]EL��S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��_    � �8LN0��LMP�;�L{�7!l��]��A]EL��S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��_    � �8LN,��LMH�7�L{�8!l��]��A]EL��S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��_    � �8LN$��LMD�7�L{�9!l��]��A]EL��S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��_    � �8LN��LM<�3�L��:!l��]��A]EL��S��AR�Z���T0 k� ������ 2d q&�1D"3Q  $�_    � �8LN�ےLM8�/�L��;!l��]��A]C���S��AR�Z���T0 k� <����� 2d q&�1D"3Q  ��X    � �8LN�דLM4�/�L��<!l��]��A]C���S��AR�Z���T0 k� <{��� 2d q&�1D"3Q  ��X    � �8LN �ϔLM,�+�L��=!l��]��A]C���S��AR�Z���T0 k� <k��o� 2d q&�1D"3Q  ��X    � �8LN �˔LM(�'�L��>!l��]��A]C���S��AR�Z���T0 k� <_��c� 2d q&�1D"3Q  ��X    � �8LM�!�ÕLM$�'�L��?!l��]��A]C���S��AR�Z���T0 k� <S��W� 2d q&�1D"3Q  ��X    � �8LM�"���LM �#�L��@!l��]��A] C�{�S��AR�Z���T0 k� �K��O� 2d q&�1D"3Q  ��X    � �8LM�"���LM��L��A!l��]��A] C�s�S��AR�Z���T0 k� �?��C� 2d q&�1D"3Q  ��X    � �8LM�#���LM��L��B!l��]��A\�C�g�S��AR�Z���T0 k� �7��;� 2d q&�1D"3Q  ��X    � �8LM�#���LM��L��C!l��]��A\�C�_�S��AR�Z���T0 k� �+��/� 2d q&�1D"3Q  ��X    � �8LM�$���LM��L��C!l��]��A\�C�S�S��AR�Z���T0 k� ���#� 2d q&�1D"3Q  ��X    � �8LM�$���LM��L��D!l��]��A\�C�K�S��AR�Z���T0 k� ���� 2d q&�1D"3Q  ��X    � �8LM�%���LM ��L��E!l��]��A\�C�?�S��AR�Z���T0 k� ���� 2d q&�1D"3Q  ��X   � �8LM�&���LL� ��L�|F!l��]��A\�C�7�S��AR�Z���T0 k� ���� 2d q&�1D"3Q  ��X    � �8LM�&���LL� ��L�|G!l��]��A\�C�/�S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8LM�'���LL�!��L�|G!l��]��A\�C�#�S��AR�Z���T0 k� ���� 2d q&�1D"3Q  ��X    � �8LM�'��LL�!��L�xH!lð]��A\�C��S��AR�Z���T0 k� ���� 2d q&�1D"3Q  ��X    � �8LM�(�w�LL�"��L�xI!lï]�A\�C��S��AR�Z���T0 k� �ߪ�� 2d q&�1D"3Q  ��X    � �8LM�(�o�LL�"��L�xJ!lǮ]�A\�C��S��AR�Z���T0 k� �ש�۩ 2d q&�1D"3Q  ��X    � �8LM�)�k�LL�#��L�xJ!lǭ]{�A\�C���S��AR�Z���T0 k� �˧�ϧ 2d q&�1D"3Q  ��X    � �8LM�*�c�LL�#��L�tK!lˬ]{�A\�C���S��AR�Z���T0 k� �æ�Ǧ 2d q&�1D"3Q  ��X    � �8LM�*�[�LL�$��L�tL!lϬ]w�A\�C��S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8LM�+�S�LL�$���L�tL!lϫ]w�A\�C��S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8LM�+�O�LL�%���L�pM!lӪ]s�A\�C�߰S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8LM�,�G�LL�%���L�pN!lө]s�A\�C�׮S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8LM|,�?�LL�&���L�pO!lר]o�A\�EKϭS��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8LMt-�7�LL�&���L�pO!lק]o�A\�EKǫS��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8LMp-�3�LL�'���L�lP!lק]o�A\�EK��S��AR�Z���T0 k� ������ 2d q&�1D"3Q  )�X    � �8LMh.�+�LL�'���L�pP!lۦ]k�A\�EK��S��AR�Z���T0 k� ˗���� 2d q&�1D"3Q  ��X    � �8LM`/�#�LL�'���L�pQ!lۥ]k�A\�EK��S��AR�Z���T0 k� ˏ���� 2d q&�1D"3Q  )�X    � �8LM\/��LL�(���L�tQ!lߤ]g�A\�EK��S��AR�Z���T0 k� ˏ���� 2d q&�1D"3Q  )�X    � �8LMT0��LL�(���L�tR!lߤ]g�A\�I{��S��AR�Z���T0 k� ˋ���� 2d q&�1D"3Q  /�X    � �8LMP0��LL�)���L�tR!l�]g�A\�I{��S��AR�Z���T0 k� ˋ���� 2d q&�1D"3Q  ��X    � �8LMH1��LL�)���L�xS!l�]c�A\�I{��S��AR�Z���T0 k� ;����� 2d q&�1D"3Q  ��X    � �8L=D1���LL�)���L�xS!l�]c�A\�I{��S��AR�Z���T0 k� ;����� 2d q&�1D"3Q  ��X    � �8L=<2���L<�*���L�xS!l�]_�A\�I{��S��AR�Z���T0 k� ;����� 2d q&�1D"3Q  ��X    � �8L=82��L<�*���L�|T!l�]_�A\�E۫�S��AR�Z���T0 k� ;����� 2d q&�1D"3Q  ��X    � �8L=03��L<�*���L�|T!\�]_�A\�E۫�S��AR�Z���T0 k� ;����� 2d q&�1D"3Q  ��X    � �8L=(3��L<�+���L��U!\�][�A\�E۫�S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8L=$4�ۺL<�+���L��U!\�][�A\�E۫�S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X   � �8D=5�ӼL<�,���L��U!\�][�A\�Eۯ�S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8D=5�˽D<�,���L{�V!\�]W�A\�A���S��AR�Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8D=6�ǾD<�,���L{�V!\�]W�A\�A���S��AR�	Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8D=6῿D<�-���L{�W!\�]W�A\�A���S��AR�	Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8D=7��D<�-���L{�W!\�]S�A\�A���S��AR�	Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8D<�8��D<�.���L{�W!\��]S�A\�A���S��AR�	Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8D<�8��D<�.���L{�X!\��]S�A\�E���S��AR�	Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8D<�9��D<�/���DۈX���]O�A\�E���S��AR�	Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8D<�:��D<�/���DیY���]O�A\�E���S��AR|	Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E��;��E�|0���DیY���]O�A\�E���S��AR|	Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E��;��E�x1���DېY���]K�A\�E���S��AR|	Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E��<��E�t1���DېZ���]K�A\�F��S��AR|	Z���T0 k� ����û 2d q&�1D"3Q  ��X   � �8E��=�w�E�p2���F�[���]K�A\�F��S��AR|	Z���T0 k� �Ǻ�˺ 2d q&�1D"3Q  ��X    � �8E��=�o�E�l3���F�[���]K�A\�F��S��AR|	Z���T0 k� �ϻ�ӻ 2d q&�1D"3Q  ��X    � �8E��>�g�E�h4���F�\���]G�A\�F��S��ARx	Z���T0 k� �׼�ۼ 2d q&�1D"3Q  ��X    � �8E�?�c�E�d4���F�\���]G�A\�F��S��ARx
Z���T0 k� �۽�߽ 2d q&�1D"3Q  ��X    � �8E�@�[�E�\5���F�]���]G�A\�B[��S��ARx
Z���T0 k� �׾�۾ 2d q&�1D"3Q  ��X    � �8E�@�S�E�X6���E��]���]C�A\�B[��S��ARx
Z���T0 k� �׿�ۿ 2d q&�1D"3Q  ��X    � �8E��A�K�E�T7���E��^���]C�A\�B[��S��ARx
Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E��BC�E�P8���E��^���]C�A\�B[��S��ARx
Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E��C;�E�L9���E��_���]C�A\�B[��S��ARx
Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E��C3�E�H:���E��_���]?�A\�B[��S��ARx
Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E��D/�E�D;���B��`���]?�A\�B[��S��ARt
Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E��E'�E�@<���B��a���]?�A\�B[��S��ARt
Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E�|F�E�<=���B��a���]?�A\�B[øS��ARt
Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E�xG�E�8>���B��a���]?�A\�B[ùS��ARt
Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E�pG!�E�4?���B��b���];�A\�BkǺS��ARt
Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E�pG!�E�0@���B��b���];�A\�Bk˻S��ARt
Z���T0 k� ������ 2d q&�1D"3Q  ��X    � �8E�lH!�E�(A���B��c���];�A\�BkϼS��ARt
c��T0 k� ������ 2d q&�1D"3Q  ��X    � �8FhI ��F$C���B��c���];�A\�BkϾS��ARt
c��T0 k� ������ 2d q&�1D"3Q  ��X    � �8F`K ��F D���B��d���]7�A\�BkӿS��ARp
c��T0 k� ������ 2d q&�1D"3Q  ��X    � �8F\L ��FE̿�B��d���]7�A\�Bk��S��ARp
c��T0 k� ������ 2d q&�1D"3Q  ��X    � �8FXM ��FF̿�B��e���]7�A\�Bk��S��ARpc��T0 k� ������ 2d q&�1D"3Q  ��X    � �8FPO ��FH̿�B��f���]7�A\�Bk��S��ARpc��T0 k� ������ 2d q&�1D"3Q  ��X    � �8FLQ��FI̻�B��f���]3�A\�Bk��S��ARpc��T0 k� ����� 2d q&�1D"3Q  ��X    � �8FHR��FK̻�B��f���]3�A\�Bk��S��ARpc��T0 k� ���� 2d q&�1D"3Q  ��X    � �8FDS��FL̻�B��g���]3�A\�B{��S��ARpc��T0 k� ���� 2d q&�1D"3Q  ��X   � �8F@U��FM<��B� g���]3�A\�B{��S��ARpc��T0 k� ���� 2d q&�1D"3Q  ��X    � �8F<V��F N<��B�h���]3�A\�B{��S��ARpZ���T0 k� ���� 2d q&�1D"3Q  ��X    � �8E�8W��E��P<��B�h���]/�A\�B{��S��ARlZ���T0 k� ���� 2d q&�1D"3Q  ��X    � �8E�4Y��E��Q<��B�h���]/�A\�B{��S��ARlZ���T0 k� ���� 2d q&�1D"3Q  ��X    � �8E�4Y��E��R<��B�j���]/�A\�H��S��ARlZ���T0 k� ���� 2d q&�1D"3Q  ��X    � �8E�4Z��E��S<��B� k���]/�A\�H��S��ARlZ���T0 k� ���� 2d q&�1D"3Q  ��X    � �8E�4Z@��E��S<��B�$l���]/�A\�H��S��ARlZ���T0 k� ���� 2d q&�1D"3Q  ��X    � �8E�4[@��E��T<��B�(m���]/�A\�H��S��ARlZ���T0 k� ���� 2d q&�1D"3Q  ��X    � �8E�4[@��E��U<��B�0n���]+�A\�H��S��ARlZ���T0 k� ���#� 2d q&�1D"3Q  ��X   � �8E�4\@��E��VL��E�4o���]+�A\�H��S��ARlZ���T0 k� �#��'� 2d q&�1D"3Q  ��X    � �8E�4\@��E��WL��E�<q���]+�A\�H��S��ARlZ���T0 k� �'��+� 2d q&�1D"3Q  ��X    � �8B�4]@��B��XL��E�@r���]+�A\�H��S��ARlZ���T0 k� �+��/� 2d q&�1D"3Q  ��X    � �8B�4]@��B��YL��E�Hs���]+�A\�H��S��ARlc��T0 k� �/��3� 2d q&�1D"3Q  ��X    � �8B�4^@��B��ZL��E�Lt���]+�A\�H�#�S��ARhc��T0 k� �/��3� 2d q&�1D"3Q  ��X    � �8B�4^@�B��[L��E�Tu���]'�A\�H�'�S��ARhc��T0 k� �3��7� 2d q&�1D"3Q  ��X    � �8B�8_@w�B��\L��E�Xv���]'�A\�H�'�S��ARhc��T0 k� �7��;� 2d q&�1D"3Q  ��X    � �8B�8_�s�B��]L��E�`w���]'�A\�H�+�S��ARhc��T0 k� �;��?� 2d q&�1D"3Q  ��X    � �8B�8`�k�B��^L��E�hx���]'�A\�H�/�S��ARhc��T0 k� �?��C� 2d q&�1D"3Q  ��X    � �8K�<`�g�B��_L��E�ly���]'�A\�H�3�S��ARhc��T0 k� �C��G� 2d q&�1D"3Q  ��X    � �8K�<a�_�B��`L��E�tz���]'�A\�H�7�S��ARhc��T0 k� �C��G� 2d q&�1D"3Q  ��X    � �8K�<a�[�B��aL��E�|{���]'�A\�H�7�S��ARhc��T0 k� �G��K� 2d q&�1D"3Q  ��X    � �8K�@b�S�B��b\��E��{���]#�A\�H�;�S��ARhc��T0 k� �?��C� 2d q&�1D"3Q  �X    � �8K�@b�O�B��c\��E��|���]#�A\�H�?�S��ARhc��T0 k� �3��7� 2d q&�1D"3Q ��_    � �8K�Dc�G�B� d\��E��}���]#�A\�H�C�S��ARhZ���T0 k� �+��/� 2d q&�1D"3Q ��_    � �8K�Dc�?�B� e\��E��}���]#�A\�H�C�S��ARhZ���T0 k� �#��'� 2d q&�1D"3Q ��_    � �8K�Dd�;�B�f\��E��~���]#�A\�H�G�S��ARhZ���T0 k� ���� 2d q&�1D"3Q ��_   � �8K�Hd�3�B�g\��E��~���]#�A\�H�K�S��ARhZ���T0 k� � �  2d q&�1D"3Q ��_    � �8K�He�+�B�g\��E�����]#�A\�H�K�S��ARdZ���T0 k� �� 2d q&�1D"3Q ��_    � �8K�He�'�B�g\��E�����]#�A\�H�O�S��ARdZ���T0 k� ���  2d q&�1D"3Q ��_    � �8K�Lf��B�h\��E�����]�A\�H�S�S��ARdZ���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�Lf��B�i\��E������]�A\�H�S�S��ARdZ���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�Pg��E�j\��E�Ȁ���]�A\�H�W�S��ARdZ���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�Pg��E�jl��E�����]�A\�H�[�S��ARdZ���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�Th��E�kl��E�����]�A\�H�[�S��ARdZ���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�Xh���E�ll��E��~���]�A\�H�_�S��ARdZ���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�Xi���E�ml��E��~���]�A\�H�c�S��ARdZ���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�\i���E�ml��E��}���]�A\�H�c�S��ARdZ���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�\j���E�nl��CL�}���]�A\�H�c�S��ARdZ���T0 k� ���� 2d q&�1D"3Q	 ��_    � �8K�`j���E� oܧ�CL�|���]�A\�H�c�S��ARdZ���T0 k� ���� 2d q&�1D"3Q	 ��_    � �8K�dj���E�$oܧ�CL�|���]�A\�H�c�S��ARdZ���T0 k� ���� 2d q&�1D"3Q	 ��_    � �8K�dk�� E�$oܧ�CM {���]�A\�H�c�S��ARdZ���T0 k� ���� 2d q&�1D"3Q	 ��_    � �8K�hk��E�(pܫ�CMz���]�A\|H�g�S��ARdZ���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K�ll�E�(pܫ�CMy���]�A\|H�g�S��ARdZ���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K�ll�K�,qܫ�E�y���]�A\|H�g�S��ARdZ���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K�pl�K�0rܯ�E�x���]�A\xH�g�S��ARdZ���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K�tm�K�4rܯ�E�w���]�A\xH�g�S��ARdZ���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K�tm�K�4sܳ�E� v���]�A\xH�g�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K�xn�K�8sܳ�E�$u���]�A\xH�g�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K�|n�K�<tܳ�E�,t���]�A\tBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K�|o�K�<tܷ�E�0s���]�A\tBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K��o�	K�@uܷ�E�4r���]�A\t	BLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K��o�x
K�Duܷ�E�8q���]�A\t
BLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K��p�pK�Dv��E�@o���]�A\t
BLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K��p�hK�Hw� E�Dn���]�A\pBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K��q�`K�Hw� E�Hm���]�A\pBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K��q�XK�Lx�E�Ll���]�A\pBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K��q�PK�Px�E�Pj���]�A\pBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q
 ��_    � �8K��rOHK�Py�E�Ti���]�A\pBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q	 ��_    � �8K��rO@K�Ty��E�Xh���]�A\lBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q	 ��_    � �8K��rO8K�Ty��E�Xf���]�A\lBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q	 ��_    � �8K��sO0K�Xz��E�\e���]�A\lBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q	 ��_    � �8K��sO(K�\z��E�`d���]�A\lBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��tO K�\{��E�db���]�A\lBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��tOK�`{��E�da���]�A\hBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��t�K�`|��E�h`���]�A\hBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��u�K�d|��E�h^���]�A\hBLg�S��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��u� K�d}��	E�l]���]�A\hBLd S��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��v��K�h}��	E�l[���]�A\hBLd S��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��v��K�h}��
E�pZ���]�A\hBLdS��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��v��K�l~��E�pY���]�A\dBLdS��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_   � �8K��w��K�l~��LtW���]�A\dBLdS��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��w��K�p��LtV���]�A\dBLdS��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��x��K�p��LxU���]�A\dBLdS��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��x��K�t��LxT���]�A\dBLdS��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��x��K�t���LxR���]�A\dBLdS��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��y޼ K�t���L|Q���]�A\`BLdS��AR`Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K��y� K�x��L|P���]�A\`BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��z�!K�x��L�O���]�A\`BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��z�"K�|��L�N���]�A\`BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ,�_    � �8B��z�#K�|��L�M���]�A\`BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8B��{�$K̀~��L-�L���]�A\`BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8B��{N�%K̀~��L-�K���]�A\`BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8B��{N�%K̀~��L-�I���]�A\\BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8B��|N|&K̄~��L-�H���]�A\\BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E��|Nt'K̄}��L-�G���]�A\\BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E��}Nl(K̈}��L-�F���]�A\\BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E��}Nd)K̈}��L-�E���]�A\\BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E��}N\*K̈}��L-�D���]�A\\BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E��~�T+Ǩ}��L-�C���]�A\\BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E��~�L,Ǩ|��L-�B���]�A\\BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E��~�D-Ǩ|��L-�B���]�A\XBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E��~�<.K̐|��L-�A���]�A\XBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E� ~�4/K̐|��L-�@���]�A\XBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E�~�00K̐|��L-�?���]�A\XBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E��(1K̔{��L-�>���]�A\XBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_   � �8E�� 2K��{��L-�=���]�A\XBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E��3K��{��L-�<���]�A\XBLd	S��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E�~�4K��{��L-�;���]�A\XBLd	S��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8E�~�5K��{��L-�;���]�A\XBLd	S��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_   � �8E�$~� 6K��zL�L-�:���]�A\XBLd	S��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�(~��7K��zL�L-�9���]�A\TBLd
S��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�,~��8B��zL�L-�8���]�A\TBLd
S��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�0~��9B��zL�L-�7���]�A\TBLd
S��AR\Z���T0 k� ���� 2d q&�1D"3Q ��_    � �8K�8~��:B��zL�L-�7���]�A\TBLd
S��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�<~��:B��yL�L-�6���]�A\TBLd
S��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�@~��;B��yL�L-�5���]�A\TBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�D~��<E��yL�L-�4���]�A\TBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  /�_    � �8K�H~��=E��xL�L-�3���]�A\TBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�P~��=E��xL� L-�2���]�A\TBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�T~��>E��wL�!L-�1���]�A\TBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�X~��?E��wL�"L-�0���]�A\TBLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_   � �8K�\~��@E��v\�#L-�0���]�A\P BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�`~��AE��v\�$L-�/���]�A\P BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�h~��BE��u\�%L-�.���]�A\P BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�l}�BE��t\�&L-�-���]�A\P BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�p}�CE��s\�(L-�,���]�A\P BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�t}�DCL�s\�)L-�,���]�A\P!BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�x}�ECL�r\�*L-�+���]�A\P!BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}�ECL�q\�,L-�*���]�A\P!BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}�FCL�p\�-L-�)���]�A\P!BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}�GCL�o\�/L-�)���]�A\P!BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}�HCL�n\�0L�(���]�A\P"BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}�HCL�ml�2L�'���]�A\P"BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}�ICL�ll�4L�'���]�A\P"BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}�JCL�kl�5L�&���]�A\P"BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}�JCL�jl�7L�%���]�A\L"BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}�KC\�hl�9L�%���]�A\L#BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}-�KC\�gl�;C�$���]�A\L#BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}-�LC\�f	\�=C�#���]�A\L#BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}-�MC\�e	\�>C�#���]�A\L#BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_   � �8K�}-�MC\�d	\�@C�"���]�A\L#BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�}-|NI\�c	\�AC�"���]�A\L#BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-xOI\�b	\�CE݀!���]�A\L$BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-tOI\�a	\�DE݀!���]�A\L$BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-pPI\�`	l�FE�| ���]�A\L$BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-lPI\�_	l�GE�x ���]�A\L$BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-lQIl�_	l�HE�x���]�A\L$BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-hQIl�^	l�IE�t���]�A\L$BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-dRIl�]	l�KE�p���]�A\L$BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-`RIl�]	\�LE�p���]�A\L%BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-`SIl�\	\�ME�l���]�A\L%BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-\SI\�\	\�NE�h���]�A\L%BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-XTI\�\	\�NE�d���]�A\L%BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-XTI\�\	\�OE�d���]�A\H%BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-TUI\�\	l�OE�`���]�A\H%BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K��|-PUI\�\	l�OE�\���]�A\H%BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_   � �8K� |-PVIl�]	l�OE�X���]�A\H&BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�|-LVIl�]	l�PE�T���]�A\H&BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�|-HWIl�]	l�PE�P���]�A\H&BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_    � �8K�|-HWIl�]	\�PE�L���]�A\H&BLdS��AR\Z���T0 k� ���� 2d q&�1D"3Q  ��_   � �8                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��� ]�(�(� � � pd�  > >    ����
     p�)��`u    �q�            Z�8          �p�     ���   H


 

           a=R   > > 
	   ��D�     a=R�D�           	         "	 Z�8         `  �  ���    	!
           \�  � �	    �4��     \��4��           
         F	 Z�8�        �@�     ���  H
           PΒ   � �	    �>��     PΒ�>��    �                	 Z�8          �P�  (  ���   0	 

          >%�  J J
     .�>1(     >���>�E    ���             # Z�8          ��  
  ���   @	
          ���4  11      B�=SX    ���4�=SX                              �@             �  ���    8

 '            ��[          V�A�H    ��[�A�      ��              	  I �         �     ��@   0
&


          )۸         j���     )����    ,��                 �         �     ��@   (
 
           n� $ $       ~��v     ^6��v     �                � A         ـ     ��H   0	
          ��I�   H	      � ���    ��I� ���                    	�� �         	 �     ��@   H	$
          �M  S	     � �%�     �M �%�                        
    �         
 `     ��@   03 
          ������	      � ��v    ���� ��v                           	  ���b             O  ��@    P		 5                   ��      �                                                                           �                               ��        ���          ��                                                                 �                          �t  ��        ���p�     �{��a�    i�� "                  x                j  �   �   �                              ��        ���         ��           "                                                �                         ���D�4�>�>�=�A�� � � �������  
     	          
  <   �R� ��C       �� �`� �� a� �� 0a� �D  b@ �� b� 1d g  GD `[� H 0\� Hd \� H� ]  �D d����< ����J ����X � 
�| V ���� � �  u� 
�< V� 
�� V� 
�\ W  
�< W� 
�| W� 
�\ W� � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }`���� � �� ^� � `^� �� _` �� _� � _� 	�� `t� 	�d u� 	�� u� 	��  u� �� w@ � �w` �$ x� �$ �e� �$ f� �D f� �d g  Є g  Ф g@ �� �`� �� a� � a� �$  b  �d b@ �� b` �� �c@ ¤ 0d@ � d� �$ d� �  }` �D  }����� � 
�\ W  
�| W� 
�| W� 
�| W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����8�� �� �  ������  
�fD
��L���"����D" � j  "  B   J jF�"      �j * , .��
��
��"   "D�j�
�� " �
� �  �  
� ��    ��     ��  �   ��   ��     ��=           ��     ��      ��  � ��   � � 	�         LL     �    ��        MM     �    ��        a�         �    ��  �_ '      �� �T ���        � � �  ���        �        ��        �        ��        �    ��    ���� 
��        ��                         T�) , 	�� ��                                     �                 ����             ��� ���%��   �8��           �    16 Brett Hull ne                                                                                    4  4      �� �� �% � �$ � �kj" kr �k~  k� �	KH � 
K@ �K0 �K8 � KM �CB � �CF � � CJ { �C: � C"J �C#J �C&J � C(= �K.) �K69 � K8! �cV p � c^ x �B�L � B�\ tJ�[ } J�S �"� � �  "� � �!"� } �"*� �#"� � $"�
%� �
&
�X '"K s8 (*D{X  *KkX  *HkH +*PkX  *Hk
-
�@  *Gs
/
�@  *Gs@  *Hs8 2*L{X  *KkH 4*PkX  *Hk �6� � �7
� � x8" � �  *Hg {:" � �  *Hg �  *R{ �=*(s � >*Qs �  )�{                                                                                                                                                                                                                         �� P        �    @ 
        �     _ P E d  ��                    �������������������������������������� ���������	�
��������                                                                                          ��    �L�� ��������������������������������������������������������   �4, C  < �� ��� � � �� ��)��@�A��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       D    ,     ��  0$�J      �  	                           ������������������������������������������������������                                                                                                                                        �    ��                     r��                  
   ���� � �������������  � ���������� �������������� �������������� � ���� ���������������������������� � �������������� ���������������������� � ����������� ������ � ��������� �������������������������������� ���� ������ ���������������                                  (    7         D��J      VT                              ������������������������������������������������������                                                                                                                                      	      �    ���                        �  �            
 	    ��������������������������������� �������������������������������� ��� ����� ���������  �   ��������� ������ �� � � ��������������� ��������������� ��������������� ���� ����� ���������������� �������������� ���������������                                                                                                                                                                                                                                                                                              
         	                    �             


             �   }�         ���.                Y�                                Z  0�  Z                     ������������  V      L*��������������������������������������������������������  6���������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 8 F <                                  � J��  �`�                                                                                                                                                                                                                                                                                        YY	�  E�                m                  b            m                                                                                                                                                                                                                                                                                                                                                                                                                       Z �  Z�  0�  
N  (�  Bm	 �� � �V ����  �˶�w��H���� ������������                ���D : � |          �   &  AG� �   �                    �                                                                                                                                                                                                                                                                                                                                        7 H           ,             !��                                                                                                                                                                                                                            Y��   �� �� ��      �� @      ���� � �������������  � ���������� �������������� �������������� � ���� ���������������������������� � �������������� ���������������������� � ����������� ������ � ��������� �������������������������������� ���� ������ ������������������������������������������������ �������������������������������� ��� ����� ���������  �   ��������� ������ �� � � ��������������� ��������������� ��������������� ���� ����� ���������������� �������������� ���������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     C   !   C    �                         @     �   ���������J      ��     ��         �      �      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �� ��  � ��     � ��   	 ��   p �� �� ��  � ��     �� �� �z     `d �$ ^$ �@    ��    ��   ~ � ��     ��   � ��     � �����6�������� J ��   	 ��  �  ��  �� �� `� �� �� �z `� �� �$   ��       �  ��   �������2���� g���        f ^�         ���             �����2�������J��1 ���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                                                         �� �����虙������(��������������񙙘�!                �  �������                           �       �  "(� """ �"" ""  "   �      �   �"��"""�"""�"""�"""�����������������������������������""�".�"/��"���!���.���/���-���""����������.���-������/�������   ��  �  .� /�� "�� "� "-�                                ""�  �(��""! ("" �"  �"   ����������������陙����.��� 陙/���.���"���"!��"��".���!♒""����������������̎���""�""",""/ �-� /� "�� "�� . /� �                    �                                           ""陂".��""� � �          �"(��(""������� ��        ""!�"!������������           ��     �                       wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  "!  " ! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """"! "   "      ""                                                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  "!  " ! " ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         � 
��	�˽���w��{k��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            �  �  �  ��  �           K�  ��� ڬ� ۻ� +�" """ """ �"" ��"/����� ��   ��  ��  ��                        �          �   � � �  ��� ��  �                                                     �               �  �  ��  �   �   �                             �   �  �      � �������������               �  �     �   �  �  �                     �   �� �       �  �  ��  �   �   �   �                                     � 
��	�˽���w��{k��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            �  �  �  ��  �           / �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw     �� ���  ��                    ���� �                                                                                                                                                                                         w 
�� ɚ� ���
�˻Ɋ�����������-� �"+ ". "$ "$ �U  Z�  Z�  J�  J�  �D  ��  ��  ɘ ˰ "  �"/�"" "  �  �            g���z��ȩ�����ة�� ���  ̰  ̰  ˰  ��  �  N�� T4�CD  CD0 C40 C30 3;� ܰ �� �� �  �  "  �""�"" �"/���  � �  �      �     �   �   ��  �"" �""  ""   "                 �   ��   �                            � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���    �   ��  �   ��   �       �                                                                                                                                  w 
�� ɚ� ���
�˻Ɋ�����������-� �"+ ". "$ "$ �U  Z�  Z�  J�  J�  �D  ��  ��  ɘ ˰ "  �"/�"" "  �  �            g���z��ȩ�����ة�� ���  ̰  ̰  ˰  ��  �  N�� T4�CD  CD0 C40 C30 3;� ܰ �� �� �  �  "  �""�"" �"/���  � �  �      �     �   �   ��  �"" �""  ""   "                 �   ��   �                            � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                                                                                                                                                                �  �˰ ��� w�� k}� gg��j�� ���
���	������ ��� ���˸�,̽�+�ӊ��8� �D 8�U�E �@ �� 	��  ��  � "" """/���  �                                 �   ��  ��  ��  ��� ̽� ̉  ɘ  �40 DD@ EU@ S3C  4M  ��  ��  *�  "�  "  ����� � �  �                          �   �                           �   �  "������"    /   �  �   ��                                �   �                      �������  ���    �    �����                                            "  "  "    �   ��  ���  � �    �                                                                                                                                              ̰ �̽ ͻ���ݪ�	������������ ˍ� ��� ��̌�����˘����� D� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��              �  �˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                     �  ��  �� ��  ��/�� �                                         �  ��  �� ��  ���ڀ �Ͱ ��� �� �̰��˰ ��� ���                     �                               �   �   ��  ���   ˰  ̹  ��@ ��UP�EEXDTD��         �  �� �  �� ��                                                                                                                                       	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w"   "   "  �� ��                   ����������                                ��  ��  ���                                                                                                                                                                                                  	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                       �  ��  �       �       �                "   "   "  �� ��                   ����������                                ��  ��  ��� ���                                                                                                                                                                                                  �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �                         �� �  �        �  �  ��  �   �                              �   �                      �������  ���    �              �  �� ��  �    � ���                                                �   ���                            �   �                                                                                                   ̰ �� ̻ {�����vz� w��  ��  ��  ̘  	�  
� "��,̻�"�� "#3  34  D  
�  �  " "" """ ! ��  ��                               ˹� �ɩ ��� �͋ ��� ��� ��̀��Ȑ���лܹнȝ0ݙ�@43�PCD�@@E�@ E�@ U�� H�  K�  �   ��    �� "�" ���                          �  �   ��  �  ��                �   �   �   "   "   "  !�    ��                              �                        ���� ��� ����                            ��  ��  ���                   ���                                      ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                     	�  �� �� ���ܙܽɪ�͚�����͙ͼ̨��̄DC"�D32�C33�333�33P330X̽ 
�� ˪  "   ""/"""�����vv ��p ��  ��  ̽  ˸  ɚ  ��  ؛  -�� .ܰ .��  �"  �   .   "�                   � �  ��            Z   Z   Z   Z  Z  �� �� �� "� "" "" ""/ ����   �   � ���� �� ����                    �� ��������p��}`     �  ��  ��  ww  ��  vv  w"   "   "  �� ��                   ����������                    � ��                    ���� �                           �   ��  ���  � �    �                                                                                                                                         �   � �� ˚�̹����	��̚���ȭ�̻������ �� H�� �ED�EU�UDDT3�EDӻ�Cݻ�ؽ����ݽ	�ݍ����ݲ �ݰ�ۏ��/��"  ���      ���  w�  ��  ��� ��� ��� ͻ���ة��ڌ�̽���������虄�DD �DC"33��33� 3;� ��� ً� ݸ  ��� ٲ �ݲ  �"� "/  �� �   �      �           �   �   �   ɀ  ��  ��                          �� �� �� +�"�"/� ��      �             ��     �   �  ��  ��  �   �            �   �   �   �    �                             �          �                        �         �  �� �  �� ��                                                                                                                                                   �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""��������D�M����""""�������D�M�M""""�����AMAD������""""��������D��""""������MM�����""""���������D�""""������������������""""������������������������"""$���4���4���4���4���4���4ffffffffffffffffff333DDDffffffffffffffffffffffff3333DDDDafaafffaffDDffff3333DDDDfFfFDfFFfFffdFffff3333DDDDfaffaffaffafffDfffff3333DDDDADAFaFadFfDffff3333DDDDafffDfdFdffff3333DDDDDDFFDfFFfdFffff3333DDDDAffAffaffafffDffffff3333DDDDffffffffffffffffffffffff3333DDDDfff4fff4fff4fff4fff4fff43334DDDD"""������������������""""������������������������""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""���������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��������������D�����3333DDDDI����D��DI����3333DDDDADAIA����D������3333DDDD��������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=LL����������D����3333DDDD    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����������A������ x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx""""�������I�I������ w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww""""�������I��D���I�������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(�D�M�D���M������3333DDDD �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""�����AMAD������ M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M""""������������������ � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�fFfFDfFFfFffdFffff3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DDFFDfFFfdFffff3333DDDD 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5""""wwwwwwwGGD x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x""""wwwwwwqwAqwAwA w w x y�������H���������������������������������H������yxww""""wwwwqwqAwAqAqAq  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(A�A�A�A��LD�����3333DDDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,�A�LDL�L�D�L�����3333DDDD +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+""""wwwwwwDGAD 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5""""wwwwqqDAAq =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=""""wwwwwwwGGwGGwGwGw     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( UQUUQUUQUUQUUUDUUUUU3333DDDD � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � �DEQQUUDUTEUUUU3333DDDD � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � �""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq� �� �% � �$ � �kj" kr �k~  k� �	KH � 
K@ �K0 �K8 � KM �CB � �CF � � CJ { �C: � C"J �C#J �C&J � C(= �K.) �K69 � K8! �cV p � c^ x �B�L � B�\ tJ�[ } J�S �"� � �  "� � �!"� } �"*� �#"� � $"�
%� �
&
�X '"K s8 (*D{X  *KkX  *HkH +*PkX  *Hk
-
�@  *Gs
/
�@  *Gs@  *Hs8 2*L{X  *KkH 4*PkX  *Hk �6� � �7
� � x8" � �  *Hg {:" � �  *Hg �  *R{ �=*(s � >*Qs �  )�{3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������.�G�R�K��2�G�]�K�X�I�N�[�Q� � � � � � ��=�@�������������������������������������������=�K�K�S�[��<�K�R�G�T�T�K� � � � � � � �=��;�����������������������������������������!��,�X�K�Z�Z��2�[�R�R� � � � � � � � � � ��=�@�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������=��;� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ������������������=�@� ��!������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������,�-��.�/�0�1�2������������������������� �!�"�3�4�#�#�#�#�#�#�#�#�$������������������%�&�'�(�)�)�)�)�)�)�)�)�)�)�*�+������������������5�6���7�8�9�:�;�<�=�>�?�������������������� �!�"�#�#�#�#�#�#�#�@�4�#�$������������������%�A�B�C�D�E�F�G�H�I�J�K�L�M�N�O�����������������P�Q�R�S�T�U�V�W�X�Y�W�Z�[�\�]�^��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            