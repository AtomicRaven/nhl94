GST@�                                                            \     �                                               �����     �  ��  �        ���2�������ʳ������������������        6i     #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF��    
 �j@ b ����
��
��     �j�� (*&��
  �                                                                               ����������������������������������      ��    a bQb  111  c c  	     
                g  	                  �$ !2"         =:=�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             FF  )          == �����������������������������������������������������������������������������                                 d  �   d  d�   @  #   �   �                          �                                                     '    !�2"$  )FF    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�=O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE | �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ރ�Iob��-��	�P=Z3��1���C�`%�<z�t|C�T0 k� �\�`	e2D Q%1D"Q  ��     � �J�{�Iob��-���L=Z3��1���C�X%�8z�p|C�T0 k� �W��[�	e2D Q%1D"Q  ��     � �H�s�Iob��-���H=Z3��1���C�L%�4{�l|C�T0 k� �O��S�	e2D Q%1D"Q  ��     � �G�k�Iob��-���D=Z3��1���C�D%�4{�h|C�T0 k� �G��K�	e2D Q%1D"Q  ��     � �F�c�Iob��-���@=Z3��1���C�8%�0|�h|C�T0 k� �;��?�	e2D Q%1D"Q  ��     � �E�[�I_b�-���<=Z3��1��C�0%�0|�d|C�T0 k� �3��7�	e2D Q%1D"Q  ��     � �D�S�I_b�-���8=Z3��|1��C�$%�,{�`|C�T0 k� �+��/�	e2D Q%1D"Q  ��     � �C�K�I_b�-���4=Z3��t1��C�%�,{�\|C�T0 k� �#��'�	e2D Q%1D"Q  ��     � �B�C�I_b�-���0=Z3��l2��C�%�({�X|C�T0 k� ����	e2D Q%1D"Q  ��     � �A�;�I_b�-���,=Z3��d2��C�%�({�P|C�T0 k� ����	e2D Q%1D"Q  ��     � �@�3�C�b�-���$=Z3��\2��C� %�$z�L|C�T0 k� ����	e2D Q%1D"Q  ��     � �?�+�C�a�|-��� =Z3��P2��C��%�$z�H|C�T0 k� ����	e2D Q%1D"Q  ��     � �>�#�C�a�t-���=Z3��H2��D�%
N z�D|C�T0 k� �����	e2D Q%1D"Q  ��     � �=��C�a�l-���=Z3��@2�s�D�%
N y�@|C�T0 k� ������	e2D Q%1D"Q  ��     � �<��C�a�`-���=Z3��82�k�D�%
Ny�8|C�T0 k� ������	e2D Q%1D"Q  ��     � �;��C�a�X-���=Z3�02�c�D�%
Ny�4|C�T0 k� ������	e2D Q%1D"Q  ��     � �:���C�`�P-���=Z3�(2�[�D�%
Nx�0|C�T0 k� ������	e2D Q%1D"Q  ��     � �9�� C�`�H-��� =Z3� 3�O�EO�%
Nx�(|C�T0 k� ������	e2D Q%1D"Q  ��     � �8�� C�_�@-���=Z3�3�G�EO�%
Nw�$|C�T0 k� ������	e2D Q%1D"Q  ��     � �8�� C�_�4,����=Z3�3�?�EO�%
Nw|C�T0 k� ������	e2D Q%1D"Q  ��     � �8�� E�^�$,���=Z3� 3�+�EO�%
Nv|C�T0 k� ������	e2D Q%1D"Q  ��     � �8��E� ]?,���=Z3� �3�#�EO�$
Nu|C�T0 k� ������	e2D Q%1D"Q  ��     � �8��E� ]?+���=Z3� �3��EO�$
N u|C�T0 k� ������	e2D Q%1D"Q  ��     � �8��E��\?+���=Z3� �3��EOx$
]�t |C�T0 k� ������	e2D Q%1D"Q  ��     � �8��E��\? +��=Z3� �3��EOp$
]�s�|C�T0 k� ������	e2D Q%1D"Q  ��     � �8��E��[>�*{��=Z3��3��C�d#
]�r�|C�T0 k� �{���	e2D Q%1D"Q  ��     � �8��E��Z>�*w��=Z3��4��C�\#
]�r�|C�T0 k� �s��w�	e2D Q%1D"Q  ��     � �8��E��Z>�*s��=Z3��4��C�P#
]�q�|C�T0 k� �k��o�	e2D Q%1D"Q  ��     � �8]� E��Y>�)o��=Z3��4��C�H" ��p�|C�T0 k� �g��k�	e2D Q%1D"Q  ��     � �8]� E��X>�)k��=Z3��4��C�@" ��o�|C�T0 k� �c��g�	e2D Q%1D"Q  ��     � �8]t C��W>�(c��=Z3��4��C�,! ��n�|C�T0 k� �S��W�	e2D Q%1D"Q  ��     � �8]l C��V>�'[��=Z3��4��C�   ��n�|C�T0 k� �H �L 	e2D Q%1D"Q  ��     � �8]d C��VN�'W��=Z3��4��C� ��m�|C�T0 k� �@�D	e2D Q%1D"Q  ��     � �8]\ C��UN�&S�|=Z3��4��C���m�|C�T0 k� �8�<	e2D Q%1D"Q  ��     � �8]T C��TN�%O�t=Z3��4��C���l�|C�T0 k� �0�4	e2D Q%1D"Q  ��     � �8]L C��TN�%G�l=Z3��|4��C����l�|C�T0 k� �(�,	e2D Q%1D"Q  ��     � �8]H C��SN�$C�d=Z3��p5��C����l�|C�T0 k� �$�(	e2D Q%1D"Q  ��     � �8]C�C�SN�$;�\=Z3��h5��C����l�|C�T0 k� ��	e2D Q%1D"Q  ��     � �8];�C�RN�#7�T=Z3��`5�C��M�l�|C�T0 k� ��	e2D Q%1D"Q  ��     � �8]+�C�QNp"�+�D=Z3��P5k�C��M�l�x|C�T0 k� ����	e2D Q%1D"Q  ��     � �8]#�C�PNh!�'��<=Z3��H5c�C��M�l�l|C�T0 k� ����	e2D Q%1D"Q  ��     � �8]�C��PN\ ���4=Z3��@5W�C��M�l�d|C�T0 k� ����	e2D Q%1D"Q  ��     � �8]�C��O^T ���,=Z3��85O�C��M�l�\
|C�T0 k� ����	e2D Q%1D"Q  ��     � �8]�C��O^L���$=Z3��05C�C��M�l�T
|C�T0 k� ����	e2D Q%1D"Q  ��     � �8]�C��N^D���=Z3��(5;�C��M�m�L
|C�T0 k� ����	e2D Q%1D"Q  ��     � �8\��C��N^<���<Z3�� 5�3�C��=�m�@	|C�T0 k� ����	e2D Q%1D"Q  ��     � �8\��C�|M^4����<Z3��5�'�C��=�n�8	|C�T0 k� ����	e2D Q%1D"Q  ��     � �8\��C�pL^$����<Z3��5��C�x=�n�(	|C�T0 k� ����	e2D Q%1D"Q  ��     � �8\��C�hL^����<Z3�� 6��C�p=�o� |C�T0 k� ����	e2D Q%1D"Q  ��     � �8\��C�`K^����;Z3���6��C�h��p�|G�T0 k� ����	e2D Q%1D"Q  ��     � �8L��C�XK^�۰��;Z3���6���I~`��p�|G�T0 k� ����	e2D Q%1D"Q  ��     � �8L��DPJ^�Ӱ��;bs���6���I~X��q�|G�T0 k� ��	��		e2D Q%1D"Q  ��     � �8L��DHJm��˰��;bs���6���I~P��q�|K�T0 k� ��
��
	e2D Q%1D"Q  ��     � �8L��D8Im����:bs���6���I~@͌p��|L T0 k� ����	e2D Q%1D"Q  ��     � �8|��D0Im����9bs���6���I�<͈p���L T0 k� �x�|	e2D Q%1D"Q  �     � �8|��D(Hm����9bs��6���I�4͈p���PT0 k� �p�t	e2D Q%1D"Q $�    � �8|��DH]����8bs��6���I�,̈́p���PT0 k� �t�x	e2D Q%1D"Q ��    � �8|��DG]����7bs��6���I� �|o���LT0 k� �x�|	e2D Q%1D"Q ��    � �8���DG]����6bs��6���EN�xo���LT0 k� �x�|	e2D Q%1D"Q  ��    � �8���D�F]�����6bs��6���EN�to]��HT0 k� �|��	e2D Q%1D"Q  ��    � �8���D�F]�{���5Z3��6݇�EN�po]��HT0 k� �|��	e2D Q%1D"Q  ��    � �8���D�E]�s���4Z3��6��EN�lo]��HT0 k� ܀��	e2D Q%1D"Q  ��    � �8���D�E]�c��x2Z3�p7�k�EM��do]��DT0 k� ܄��	e2D Q%1D"Q  ��    � �8���D�D	��[��p1Z3�h7�_�EM��`o]� �@T0 k� ܈��	e2D Q%1D"Q  ��    � �8���E]�D	��S��h0Z3�`7�W�EM�
�\o]� �@T0 k� ����	e2D Q%1D"Q  ��    � �8��E]�C	��K��d/Z3�X7�O�EM�	�To]� �@T0 k� ����	e2D Q%1D"Q  ��    � �8�{�E]�C	�|C��\.Z3�P7�C�EM��Po]��<T0 k� ����	e2D Q%1D"Q  ��    � �8�{�E]�C	�t;��X-Z3�H7�;�EM��Lo]w��<T0 k� ����	e2D Q%1D"Q  ��    � �8�w�E]�B	�p3��P,Z3�@7�/�E=��Do]o��8T0 k� ����	e2D Q%1D"Q  ��    � �8�s�EM�A	�`#��D)Z3�07��E=��<o]_��8T0 k� ����	e2D Q%1D"Q  ��    � �8�s�EM|@	�\��@(b��(7��E=��4o	�S��4T0 k� ����	e2D Q%1D"Q  ��    � �8�o�EMt@	�T��8&b�� 7��E=��0o	�K��4T0 k� ����	e2D Q%1D"Q  ��    � �8�o�EMh?	�P��4%b��7���E=��(o	�G��4T0 k� ����	e2D Q%1D"Q  ��    � �8�k�C�X>	�D��("b��7���E=� �n	�7��0T0 k� ����	e2D Q%1D"Q  ��    � �8Lk�C�L>	�<�$!b����7���E=���n	�/��0T0 k� ����	e2D Q%1D"Q  ��    � �8Lg�C�D=	�8�b����7���E=���n	�'��,	T0 k� ����	e2D Q%1D"Q  ��    � �8Lc�C�<<	�4�b����7���E=���m	�#��,	T0 k� ����	e2D Q%1D"Q  ��    � �8Lc�C�0<	�0ۨb����7���E=���m	���,	T0 k� ����	e2D Q%1D"Q  ��    � �8<[�C� :	�$�˨b����7��E=w���l	���(
T0 k� ����	e2D Q%1D"Q  ��    � �8<[�EM:	� �èZ3���8��E-s���l	���(
T0 k� ����	e2D Q%1D"Q  ��    � �8<[�EM9	�໨Z3���8���E-k���k	���$
T0 k� �� �� 	e2D Q%1D"Q  ��    � �8<X EM8	�೨ Z3��8���E-g���j	���� T0 k� ��!��!	e2D Q%1D"Q  ��    � �8�XEL�7	�ࣧ�Z3�ި8���E-_���i	����T0 k� ��"��"	e2D Q%1D"Q  ��    � �8�TEL�6	������Z3�ޠ8��E-W���h	����T0 k� ��#��#	e2D Q%1D"Q  ��    � �8�TE��5	������Z3�ޘ8�w�E-S���g	����T0 k� ��#��#	e2D Q%1D"Q  ��    � �8�TE��4	������Z3�ސ8�o�E-O���f	����T0 k� ��#��#	e2D Q%1D"Q  ��    � �8�TE��3	��{���	Z3�ހ8�_�E-G���d	����T0 k� ��"��"	e2D Q%1D"Q  ��   � �8�P	E̼2	� �s���Z3��x8�W�E-G���c	����T0 k� ��!��!	e2D Q%1D"Q  ��    � �8�P
I|�1	���k���Z3��p8�O�E-C���b	����T0 k� ��!��!	e2D Q%1D"Q  ��    � �8�PI|�1	���c���Z3��h8�G�E?���a	����T0 k� ��!��!	e2D Q%1D"Q  ��    � �8�PI|�/	���S���Z3��X8�7�E;���_	���|T0 k� �x!�|!	e2D Q%1D"Q  ��    � �8�PI|�.	���K��� Z3��P8/�E7���^���|T0 k� �p�t	e2D Q%1D"Q  �    � �8�LG|�.	���C����Z3��H8'�E7���]���|T0 k� �h�l	e2D Q%1D"Q ��    � �8�LG|�-	���;����Z3��<8�E3���[ܻ�|T0 k� �d�h	e2D Q%1D"Q ��   � �8�LG|t,	���+����Z3��,8�E3���Yܳ�|T0 k� �T�X	e2D Q%1D"Q ��    � �8�LG|l+	���#����Z3��$8�E3���Wܯ��T0 k� �L�P	e2D Q%1D"Q ��    � �8�LG�d*	�������Z3��8�E3��|Vܧ��T0 k� �D�H	e2D Q%1D"Q ��   � �8�HG�\*	�� ����Z3��8�E3��xT���T0 k� �<�@	e2D Q%1D"Q ��    � �8�HG�L)�� ����Z3��7��E3��lQ���T0 k� �0	�4		e2D Q%1D"Q ��    � �8�HG�H(�������Z3�=�7��E3��hP���T0 k� �(�,	e2D Q%1D"Q ��    � �8�HG�@'������Z3�=�7��E�3��dN���T0 k� � �$	e2D Q%1D"Q ��    � �8�HG�@'������Z3�=�7��E�3�`L���T0 k� ��	e2D Q%1D"Q ��    � �8�HG�8'��ۣ���Z3�=�6��E�7�XI�{��T0 k� ����	e2D Q%1D"Q ��    � �8�HG�4(��ӣ��Z3���6���E�7�TG�s��T0 k� ����	e2D Q%1D"Q ��    � �8�HG�0(��ˣ��Z3���5���E�;�PF�o�� T0 k� �����	e2D Q%1D"Q ��    � �8�HG�((��ã��Z3���5���E�;�LD�g���T0 k� ������	e2D Q%1D"Q ��    � �8�HG� (����Z3��4���E�?�H@�[���T0 k� ���#;P 	e2D Q%1D"Q  �    � �8�HG�)�
���Z3��4���D�C�D?�S���T0 k� ���#;P 	e2D Q%1D"Q �    � �8 �HG�),�	���Z3��4���D�C�D=�K���T0 k� ���#;P 	e2D Q%1D"Q��    � �8 �HG�),����Z3���3���D�G�@;�G���T0 k� ���#;P 	e2D Q%1D"Q��    � �8 �HG�),����Z3���3���D�G�<9�?���T0 k� ���#;P 	e2D Q%1D"Q��    � �8 �HEL),�_����Z3���2K��BMO�86�3���T0 k� ���#KP 	e2D Q%1D"Q��    � �8<HEL),�_{��#�Z3��|2K��BMO�44�/���T0 k� ���#KP 	e2D Q%1D"Q��    � �8<HEL *,�_s��'�Z3��x2K��BMS�44�'���T0 k� ���#KP 	e2D Q%1D"Q��    � �8<HEK�+,|_k��+�Z3��p1K��BMS�02�#���T0 k� ���#KP 	e2D Q%1D"Q��    � �8<HEK�+,t _c��/�Z3��h1K��BMW�01����T0 k� ���#KP 	e2D Q%1D"Q��    � �8<HN��,,s�O[��/�Z3��`1K��BMW�L,/����T0 k� ���#[P 	e2D Q%1D"Q��    � �8,LN��,,k�OS��3�Z3��\0K��BM[�L,.����T0 k� ���#[P 	e2D Q%1D"Q��    � �8,LN��.,_�OC��;�Z3��L0K��BM_�L,.����T0 k� ���#[P 	e2D Q%1D"Q��    � �8,PN��/,W�O;��?�Z3��H/K��BM_�L(-�����T0 k� ���#[P 	e2D Q%1D"Q��    � �8,TN��/,S��3��C�Z3��@/K��BMc�L(-�����T0 k� ���#kP 	e2D Q%1D"Q��    � �8�TN��0,K��+��G�Z3��8/K��BMc�L$,����T0 k� ���#kP 	e2D Q%1D"Q��    � �8�XN��1,C��#��G�Z3��4.K��BMc�L +����T0 k� ���#kP 	e2D Q%1D"Q��    � �8�\ N˼1,?����K�Z3��,.K��BMg�L *����T0 k� ���#kP 	e2D Q%1D"Q��    � �8�` N˸2,;����O�Z3��(.K��BMg�L*����T0 k� ���#kP 	e2D Q%1D"Q��    � �8�d N˴3,3����O�Z3�� .K��BMk�L)����T0 k� ���#�P 	e2D Q%1D"Q��    � �8�d!Nˬ4,/����S�Z3��-K��BMk�L(����T0 k� ���#�P 	e2D Q%1D"Q��    � �8�h!N˨4,'�����S�Z3��-K��BMo�L(����T0 k� ���#�P 	e2D Q%1D"Q��    � �8�l"Nˤ5	�#����W�Z3��-K��BMo�L(����T0 k� ���#�P 	e2D Q%1D"Q��    � �8�p#Nˠ5	�����W�Z3��,K��BMo�L(����T0 k� ���#�P 	e2D Q%1D"Q��    � �8�x$N˔7	���ۥ�[�Z3�� ,K��BMs�L'����T0 k� ���#�P 	e2D Q%1D"Q��    � �8�|%Nː7	���ӥ�[�Z3���,K��BMw�L'K����T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��%Nˌ8	���˦�[�Z3���+K��BMw�L'K����T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��&N˄9	���æ�[�Z3���+K��BMw�L'K����T0 k� ���#�P 	e2D Q%1D"Q ��   � �8��'Nˀ9	������[�Z3���+K��BM{�L'K����T0 k� ���#�P 	e2D Q%1D"Q .�    � �8��(N�|:	�������[�Z3���+K��BM{�L'K����T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��)N�x:	�������_�Z3���*K��BM�L'K����T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��*N�t;	�������_�Z3���*K��BM�L'K����T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��+Ap;	�������[�Z3���*K��BM�L'K����T0 k� ���#�P 	e2D Q%1D"Q  �    � �8��+Ap<	�������[�Z3���*K��BM��L'K����T0 k� ���#�P 	e2D Q%1D"Q ��    � �8L�,Ap=	�������[�Z3���)K��BM��L'K����T0 k� ���#�P 	e2D Q%1D"Q ��    � �8L�-At=	�������[�Z3���)K��BM��L&K����T0 k� ���#�P 	e2D Q%1D"Q ��    � �8L�.At>	������[�Z3���)K��BM��L&K����T0 k� ���#�P 	e2D Q%1D"Q ��    � �8L�/At>���Nw��[�Z3���(K��BM��L&K����T0 k� ���#�P 	e2D Q%1D"Q ��    � �8L�1At?���No��W�Z3���(K��BM��L&K���� T0 k� ���#�P 	e2D Q%1D"Q ��    � �8,�2Ax?���Ng��T Z3���(K��BM��L&K���� T0 k� ���#�P 	e2D Q%1D"Q ��    � �8,�4Ax@���NW��PZ3���'K��BM��L&K���� T0 k� ���#�P 	e2D Q%1D"Q ��    � �8,�6AxA���NO��PZ3���'K��BM��L&K����!T0 k� ���#�P 	e2D Q%1D"Q ��    � �8,�7A|A���NK��PZ3���'K��BM��L&K����!T0 k� ���#�P 	e2D Q%1D"Q ��    � �8,�8A|B���NC��LZ3���&K��BM��L%K����!T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��9A|B���>;��LZ3���&K��BM��L%K����!T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��;A|B���>3��HZ3���&K��BM��L%K��{�!T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��<A�C��>+��D	Z3���&K��BM��L%K�{�"T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��>A�C��>#��DZ3���%K��BM��L%K�{�"T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��?A�D��>��@Z3���%K��BM��L%K{�{�"T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��AA�D��>��<Z3���%K��BM��L%Kw�{�"T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��BA�E��>��<Z3���%K��BM��L%Kw� ;�"T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��CA�E��>��8Z3���$K��BM��L%Ks� ;�#T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��EA�E��>��4Z3���$K��BM��L%Ko� ;�#T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��FA�F��=���0Z3���$K��BM��L%Ko� ;�#T0 k� ���#;P 	e2D Q%1D"Q ��    � �8��HA�F��M���0Z3���$K��BM��L%Kk� ;�#T0 k� ���#;P 	e2D Q%1D"Q ��    � �8��JA�G��M��,Z3���#K��BM��L%Ko� ;�#T0 k� ���#;P 	e2D Q%1D"Q ��    � �8�KA�G���M��(Z3���#K��BM��L%Ko� ;�#T0 k� ���#;P 	e2D Q%1D"Q ��    � �8�MA�G���M��$Z3���#K��BM��L%Ko���#T0 k� ���#;P 	e2D Q%1D"Q ��    � �8�NA�H���Mۿ� Z3���#K��BM��L%Ko���$T0 k� ���#KP 	e2D Q%1D"Q ��    � �8�PA�H���M���Z3���#K��BM��L%Ks���$T0 k� ���#KP 	e2D Q%1D"Q ��    � �8�QA�H���M���Z3���"K��BM��L%Ks���$T0 k� ���#KP 	e2D Q%1D"Q ��    � �8	<�RL��I�������Z3���"K��BM��L%Ks���$T0 k� ���#KP 	e2D Q%1D"Q ��    � �8	<�TL��I�������!Z3���"K��BM��L%Ks���$T0 k� ���#KP 	e2D Q%1D"Q ��    � �8	<�UL��J���ݿ��"Z3���"K��BM��L%Ks���$T0 k� ���#[P 	e2D Q%1D"Q ��    � �8	<�VL��J���ݻ��$Z3���"K��BM��L$Kw���$T0 k� ���#[P 	e2D Q%1D"Q ��    � �8	<�WL��J���ݷ��%Z3���!K��BM��L$Kw���$T0 k� ���#[P 	e2D Q%1D"Q ��    � �8	L�XL��K���ݯ�� 'Z3���!K��BM��L$Kw���%T0 k� ���#[P 	e2D Q%1D"Q ��    � �8	L�YL��K���ݫ���)Z3���!K��BM��L$Kw���%T0 k� ���#[P 	e2D Q%1D"Q ��    � �8	L�ZL��K���ݧ���*Z3���!K��BM��L$K{���%T0 k� ���#kP 	e2D Q%1D"Q ��    � �8	L�[L��L���ݟ���,Z3���!KÖBM��L$K{���%T0 k� ���#kP 	e2D Q%1D"Q ��    � �8	L�\L��L���ݛ���.Z3��� KÖBM��L$K{���&T0 k� ���#kP 	e2D Q%1D"Q ��    � �8,�]M�L���ݗ���/Z3��� KÖBM��L$K{���&T0 k� ���#kP 	e2D Q%1D"Q ��    � �8,�^M�L���ݓ���1Z3��� KǕBM��L$K{���&T0 k� ���#kP 	e2D Q%1D"Q ��    � �8,�_M�M���ݏ���2Z3��� KǕBM��L$K���&T0 k� ���#�P 	e2D Q%1D"Q ��    � �8,�`M�M���݇���4Z3��� KǕBM��L$K���'T0 k� ���#�P 	e2D Q%1D"Q ��    � �8,�aM�M�������6Z3��� K˕BM��L$K���'T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�bM�N�������7Z3���K˔BM��L$K���'T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�cM�N����{���9Z3���K˔BM��L$K���'T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�dM�N����w���;Z3���KϔBM��L$K���'T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�fM�O����o�ݼ>Z3���KϔBM��L$K����(T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�gL��O���k�ݸ?Z3���KӓBM��L$K����(T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�hL��O���g�ݴAZ3���KӓBM��L$K����(T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�iL��O����c�ݬBZ3���KӓBM��L$K����)T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�iL��P���_�ݨDZ3���KӓBM��L$K����)T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�jL��P���[��EZ3���KגBM��L$K����)T0 k� ���#�P 	e2D Q%1D"Q ��   � �8��kL��P��W��GZ3���KגBM��L$K����)T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��lL��P��S��HZ3���KגBM��L$K����)T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��mL��Q��O��JZ3���KےBM��L$K����*T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��mL��Q��K��KZ3���KےBM��L$K����*T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��nA�Q��G��LZ3���KۑBM��L$K����*T0 k� ���#�P 	e2D Q%1D"Q ��    � �8|�oA�Q��C��NZ3���KۑBM��L$K����*T0 k� ���#�P 	e2D Q%1D"Q ��    � �8|�oA�R��?��|OZ3���KߑBM��L$K����*T0 k� ���#�P 	e2D Q%1D"Q ��    � �8|�pA�R#��;��tPZ3���KߑBM��L$K����+T0 k� ���#�P 	e2D Q%1D"Q ��    � �8|�qA�R'��7��lRZ3���KߑBM��L$K����+T0 k� ���#�P 	e2D Q%1D"Q ��    � �8} qA�R+��7��hSZ3���KߐBM��L$K����+T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}rA�R/��3��`TZ3���K�BM��L$K����+T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}rA�S7��/��\UZ3���K�BM��L$K����+T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}sA�S;��+��TVZ3���K�BM��L$K����+T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}sA�S?��'��LXZ3���K�BM��L $K����,T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}tA�S�C��#��HYZ3���K�BM��L $K����,T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}tA�S�K��#��@ZZ3���K�BM��L $K����,T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}uA�T�O����<[Z3���K�BM��L $K����,T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}vA�T�S����4\Z3���K�BM��L $K����,T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}vA�T�W����,]Z3���K�BM��L $K����,T0 k� ���#�P 	e2D Q%1D"Q ��    � �8� wA�T�[����$^Z3���K�BM��L $K����,T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�$wA�T�_���� _Z3���K�BM��L $K����-T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�$xA�U�c����`Z3���K�BMÓL $K����-T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�(xA�U�g����aZ3���K�BMÓL$$K����-T0 k� ���$P 	e2D Q%1D"Q ��    � �8�,xA�U�k����bZ3���K�BMÓL$$K����-T0 k� ���$P 	e2D Q%1D"Q ��    � �8�0yA�U�o����bZ3���K�BMÓL$$K����-T0 k� ���$P 	e2D Q%1D"Q ��    � �8�0yA�U�s�����cZ3���K�BMÓL$$K����-T0 k� ���$P 	e2D Q%1D"Q ��    � �8�4zA�U�w�����dZ3���K�BMÓL$$K����-T0 k� ���$P 	e2D Q%1D"Q ��    � �8�8zA�V�{������dZ3���K�BMÒL$$K����.T0 k� ���#KP 	e2D Q%1D"Q ��    � �8�8{A�V�����<�eZ3���K�BMÒL$$K����.T0 k� ���#KP 	e2D Q%1D"Q ��    � �8�<{A�V̃����<�eZ3���K�BMÒL$$K����.T0 k� ���#KP 	e2D Q%1D"Q ��    � �8�@|A�V̇����<�fZ3���K�BMǒL$$K����.T0 k� ���#KP 	e2D Q%1D"Q ��    � �8�@|A�V̋����<�fZ3���K�BMǒL$$K����.T0 k� ���#KP 	e2D Q%1D"Q ��    � �8�D|A�V̏����<�gZ3���K�BMǒL$$K����.T0 k� ���#[P 	e2D Q%1D"Q ��    � �8�H}A�W̓����<�gZ3���K�BMǒL($K����.T0 k� ���#[P 	e2D Q%1D"Q ��    � �8�H}A�W̗����<�hZ3���K��BMǒL($K����.T0 k� ���#[P 	e2D Q%1D"Q ��    � �8�L~A�W̛����<�hZ3���K��BMǑL($K����/T0 k� ���#[P 	e2D Q%1D"Q ��    � �8�L~A�W̟�L��<�iZ3���K��BMǑL($K����/T0 k� ���#[P 	e2D Q%1D"Q ��    � �8�P~A�W̣�L��<�iZ3���K��BMǑL($K����/T0 k� ���#kP 	e2D Q%1D"Q ��    � �8�PA�W̣�L��<�jZ3���K��BMǑL($K����/T0 k� ���#kP 	e2D Q%1D"Q ��    � �8�TA�W̧�L��<�jZ3���K��BMǑL($K����/T0 k� ���#kP 	e2D Q%1D"Q ��    � �8�X�A�X̫�L��<�kZ3���K��BMˑL($K����/T0 k� ���#kP 	e2D Q%1D"Q ��    � �8�XA�X̯�L��<�kZ3���K��BMˑL($K����/T0 k� ���#kP 	e2D Q%1D"Q ��    � �8�\A�X̳�L��L�lZ3���K��BMˑL($K����/T0 k� ���#{P 	e2D Q%1D"Q ��    � �8�\A�X̳�L��L�lZ3���K��BMːL($K����/T0 k� ���#{P 	e2D Q%1D"Q ��    � �8�`A�X̷�L��L�mZ3��|K��BMːL($K����0T0 k� ���#{P 	e2D Q%1D"Q ��    � �8�`~A�X̻�L��L|mZ3��|K��BMːL($K����0T0 k� ���#{P 	e2D Q%1D"Q ��    � �8�d~A�X̿�L��LxnZ3��|K��BMːL($K����0T0 k� ���#{P 	e2D Q%1D"Q ��    � �8�d~A�X̿�L� LtnZ3��|K��BMːL,$K����0T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�h~A�Y���\�LlnZ3��|K��BMːL,$K����0T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�h}A�Y���\�LhoZ3��|K��BMːL,$K����0T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�l}A�Y���\�LdoZ3��|K��BMːL,$K����0T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�l}A�Y���\�L`pZ3��|K��BMːL,$K����0T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�p}A�Y���\�LXpZ3��|K��BMːL,$K����0T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�p|A�Y���\�LTpZ3��|K��BMϏL,$K����0T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�t|A�Y���\�LPqZ3��|K��BMϏL,$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�t|A�Y���\�	LLqZ3��|L�BMϏL,$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�t|A�Y���\�
LHqZ3��|L�BMϏL,$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�x|A�Z���\�LDrZ3��xL�BMϏL,$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�x{A�Z���\�L<rZ3��xL�BMϏL,$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8�|{A�Z���l�L8rZ3��xL�BMϏL,$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}|{A�Z���l�L4sZ3��xL�BMϏL,$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}|{A�Z���l�L0sZ3��xL�BMϏL,$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}�{A�Z���l�L,sZ3��xL�BMϏL,$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}�{A�Z���l�L(tZ3��xL�BMϏL0$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}�zA�Z���l�L$tZ3��xL�BMώL0$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}�zA�Z���l�L tZ3��xL�BMώL0$K����1T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��zA�Z���l�LuZ3��xL�BMώL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��zA�[���l�LuZ3��tL�BMώL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��yA�[���l�LuZ3��tL�BMӎL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��yA�[���l�LvZ3��tL�BMӎL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8��yA�[���|�LvZ3��tL�BMӎL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}�xA�[���|�LvZ3��pL�BMӎL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}�xA�[���|� LwZ3��pL�BMӎL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}�wA�[���|�"LwZ3��pL�BMӎL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}�wA�[���|�#L wZ3��pL�BMӎL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8}�vA�[��ܴ%K�wZ3��pL�BMӎL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8=�uL��[��ܴ&K�xZ3��lL�BMӎL0$K����2T0 k� ���#�P 	e2D Q%1D"Q ��    � �8=�uL��[��ܴ(K�xZ3��lL�BMӎL0$K����2T0 k� ���$P 	e2D Q%1D"Q ��    � �8=�tL��[��ܴ)K�xZ3��lL�BMӎL0$K����2T0 k� ���$P 	e2D Q%1D"Q ��    � �8=�sL��\��ܴ+K�xZ3��lL�BMӍL0$K����2T0 k� ���$P 	e2D Q%1D"Q ��    � �8=�rL��\��ܴ,K�yZ3��lL�BMӍL0$K����2T0 k� ���$P 	e2D Q%1D"Q ��    � �8=�rL��\��ܰ.K�xZ3��lL�BMӍL0$K����3T0 k� ���$P 	e2D Q%1D"Q ��    � �8=�qL��\��ܰ/K�xZ3��hL�BMӍL0$K����3T0 k� ���#;P 	e2D Q%1D"Q ��    � �8=�pL��\��ܰ1;�wZ3��hL�BMӍL0$K����3T0 k� ���#;P 	e2D Q%1D"Q ��    � �8=�oL��\��ܰ2;�wZ3��hL�BMӍL4$K����3T0 k� ���#;P 	e2D Q%1D"Q ��    � �8=�oL��\��ܰ3;�vZ3��hL�BMӍL4$K����3T0 k� ���#;P 	e2D Q%1D"Q ��    � �8=�nM�\�#�ܰ5;�vZ3��hL�BM׍L4$K����3T0 k� ���#;P 	e2D Q%1D"Q ��    � �8=�mM�\�#�ܰ6;�uZ3��dL�BM׍L4$K����3T0 k� ���#[P 	e2D Q%1D"Q ��    � �8=�mM�\�'��7;�uZ3��dL�BM׍L4$K����3T0 k� ���#[P 	e2D Q%1D"Q ��    � �8=�lM�\�+��9��tZ3��dL�BM׍L4$K����3T0 k� ���#[P 	e2D Q%1D"Q ��    � �8=�kM�\M/��:��tZ3��dL�BM׍L4$K����3T0 k� ���#[P 	e2D Q%1D"Q ��    � �8=�kM�\M/��;��sZ3��dL�BM׍L4$K����3T0 k� ���#[P 	e2D Q%1D"Q ��    � �8=�jM�\M3��<��rZ3��dL�BM׍L4$K����3T0 k� ���#kP 	e2D Q%1D"Q ��    � �8=�iM�\M7��=��rZ3��dL�BM׍L4$K����3T0 k� ���#kP 	e2D Q%1D"Q ��    � �8=�iM�]M;��?[�qZ3��`L�BM׍L4$K����3T0 k� ���#kP 	e2D Q%1D"Q ��    � �8M�hL��]M;��@[�pZ3��`L�BM׍L4$K����3T0 k� ���#kP 	e2D Q%1D"Q ��    � �8M�hL��]M?��A[�pZ3��`L�BM׍L4$K����3T0 k� ���#kP 	e2D Q%1D"Q ��    � �8M�gL��]MC��B[�oZ3��`L�BM׍L4$K����3T0 k� ���#{P 	e2D Q%1D"Q ��    � �8M�gL��]MC��C[�nZ3��`L�BM׍L4$K����3T0 k� ���#{P 	e2D Q%1D"Q ��    � �8M�fL��]MG��D[�nZ3��`L�BM׌L4$K����4T0 k� ���#{P 	e2D Q%1D"Q ��    � �8M�eL��]MG��E[�mZ3��`L�BM׌L4$K����4T0 k� ���#{P 	e2D Q%1D"Q ��    � �8M�eL��]]K��F[�mZ3��`L�BM׌L4$K����4T0 k� ���#{P 	e2D Q%1D"Q ��    � �8M�dL��]]O��G[�lZ3��`L�BM׌L4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�dL��]]O��H[�lZ3��`L�BM׌L4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��   � �8M�cA�]]S��I[�lZ3��`L�BM׌L4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�cA�]]S��J[�lZ3��`L�BM׌L4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�bA�\�W��K[�lZ3��`L�BM׌L4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�bA�\�[��L[�lZ3��`L�BM׌L4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�aA�\�[��Mk�kZ3��`L�BM׌L4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�aA�\�_��Nk�kZ3��`L�BM׌L4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�`A�[�_��Ok�kZ3��`L�BM׌L4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�`A�[�c��Pk�kZ3��`L�BMیL4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��   � �8M�_A�[�c��Qk�jZ3��`L�BMیL4$K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�_A�[�g��Rk�jZ3��\L�BMیL4%K����4T0 k� ���#�P 	e2D Q%1D"Q ��   � �8M�^A�[�g��Rk�jZ3��\L�BMیL4%K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�^A�Z�k��Sk�jZ3��\L�BMیL4%K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8M�^A�Z�k��Tk�jZ3��\L�BMیL4%K����4T0 k� ���#�P 	e2D Q%1D"Q ��    � �8as�D`T��7����H_s�
�@_�S�I!�����!�C�T0 k� ����	e2D Q%1D"Q  ��U    ��� �a{�DTTS�4����T_s�
�P_�O�I!�����!�C�T0 k� ����	e2D Q%1D"Q  ��U    ��� �a�DLTS�3����X_s�
�X_�O�I$!�����!�C�T0 k� ����	e2D Q%1D"Q  ��U    ��� �a��DDTS�2����\_s�
�`_�K�I$!�����!�C�T0 k� ����	e2D Q%1D"Q  ��U    ��� �Q��D<TS�1����`	_s�
�h^�K�I$!�����!�C�T0 k� ��
��
	e2D Q%1D"Q  �U    ��� �Q��D0TS�.����h[s�
�x^�G�I$!@����!�C�T0 k� ����	e2D Q%1D"Q  ��O    ��� �Q��I�(TS�-����l[s�
��^�G�B�$!@��Û!�C�T0 k� ����	e2D Q%1D"Q  ��O    ��� �Q��I� TC�,����p[s�
��]�C�B�,!@��˜|C�T0 k� ����	e2D Q%1D"Q  �O    ��� �Q��I�TC�*����x[s�
��Z�C�B�8!@��מ|C�T0 k� 3x�|	e2D Q%1D"Q ��O    ��� �Q��I�TC�)����|[s�
��Y�?�B�<!@��ߟ|C�T0 k� 3x�|	e2D Q%1D"Q ��O    ��� �Q��I�TC�(����|[s�
��W�?�B�D!@���|C�T0 k� 3t�x	e2D Q%1D"Q ��O    ��� �Q��I� T��'���À[��
��V�?�B�L!@���|C�T0 k� 3p�t	e2D Q%1D"Q ��O    ��� �Q��I��TӼ'���ӄ[��
t�U�;�B�P!@���|C�T0 k� 3l�p	e2D Q%1D"Q ��O    ��� �Q��I��TӸ%���ӄ[��t�R�7�B�\!0� ���|C�T0 k� �h�l	e2D Q%1D"Q ��O    ��� �Q��I��TӸ%���Ӏ[��t�Q�7�B�d!0�!��|C�T0 k� �d�h	e2D Q%1D"Q ��O    ��� �A��C��TӸ$����|[��t�O�7�B�h!0�#��|C�T0 k� �`�d	e2D Q%1D"Q	 $�O    ��� �A��C��TӴ$���$�x[��t�Ld3�B�t!0�&��!�C�T0 k� �\�`	e2D Q%1D"Q	 ��O    ��� �A��C��T�#���$�t[��t�Jd/�B�t!0�'��!�C�T0 k� �\�`	e2D Q%1D"Q ��O    ��� �A��C��T�#���$�p[s�t�Id/�B�p!0�)��!�C�T0 k� �X�\	e2D Q%1D"Q ��O    ��� ����C��T�#ã�$�l[s�t�Gd+�B�p!0�*��!�C�T0 k� �X�\	e2D Q%1D"Q ��O    ��� ����C��T�#ß�$�l[s�t�Ed+�B�p!0�,��!�C�T0 k� �X�\	e2D Q%1D"Q ��O    ��� ����C�T�"ß�$�h [s�t�Dd'�B�l!0�.�#�!�C�T0 k� �T�X	e2D Q%1D"Q ��O    ��� ����C�TӨ"Û�$�d![s�d�@d#�B�l!0�1�+�!�C�T0 k� �P�T	e2D Q%1D"Q ��O    ��� �A�C�TӨ!Û�$�`![s�d�>4�B�h!0�3�+�!�C�T0 k� �P�T	e2D Q%1D"Q ��O    ��� �A�C�TӤ!×�$�\"[s�d�<4�B�h! �5�/�!�C�T0 k� �L�P	e2D Q%1D"Q ��O    ��� �A{�I��TӠ!×�$�X#[s�d�;4�B�h! �7�/�|C�T0 k� �L�P	e2D Q%1D"Q ��O    ��� �A{�I��TӜ!Ó�$�X#[s�d�94�B�d! �8�3�|C�T0 k� �H�L	e2D Q%1D"Q ��O    ��� �Aw�I��T� ӓ�$�T$[s�d�74�@dd! �:�3�|C�T0 k� H�L	e2D Q%1D"Q ��O    ��� �Ao�I�|T� Ӌ�$�P%[s�d�34�@d`!��>�7�|C�T0 k� D�H	e2D Q%1D"Q ��O    ��� �Ao�I�xT� Ӈ��L%[s�d�14�@d`!��@�7�|C�T0 k� 4�8	e2D Q%1D"Q ��D    ��� �1k�I�pT�Ӈ��H&[s�d�/4�@d`!� B�7�|C�T0 k� $�(	e2D Q%1D"Q ��D    ��� �1g�I�lTS�Ӄ��D&[s�d�/3��E�\ � D�7�|C�T0 k� � � 	e2D Q%1D"Q ��D    ��� �1c�I�`TS��{��@'[s�d�/3��E�\�H�7�|C�T0 k� �"�"	e2D Q%1D"Q ��D    ��� �1_�I�\TS|�w�c<'Zc�T�.c�E�\�J�7�|C�T0 k� � #�#	e2D Q%1D"Q ��D    ��� �A[�I�XTSx�s�c8(Zc�T�-c�E�\�L�7�|C�T0 k� ��%��%	e2D Q%1D"Q ��D    ��� �A[�I�TTSt�o�c0(Zc�T�-c�A\�N�7�|C�T0 k� �&��&	e2D Q%1D"Q ��D    ��� �AS�I�HTSh�g�c()Zc�T�+c߶A\�N�3�|C�T0 k� �'��'	e2D Q%1D"Q  ,�D    ��� �AS�I�HT�d�`c$*Zc��+c۵AX�O�3�|C�T0 k� �(��(	e2D Q%1D"Q  ��D    ��� �AO�I�HT�`�\c *Zc��*c׳AX�Q�3�|C�T0 k� �)��)	e2D Q%1D"Q  ��D    ��� �AK�I�HT�X�Tc+Zc��*cϱAT\�S�/�|C�T0 k� ��)��)	e2D Q%1D"Q  ��D    ��� �AG�I�DT�P�Ls+Zc��*cǮATX��V�+�|C�T0 k� ��+��+	e2D Q%1D"Q ��D    ��� �AC�I�DT	�L�Ds,Zc��)c��ATX��X�'�|C�T0 k� ��-��-	e2D Q%1D"Q ��D    ��� �QC�I�DT	�H�@s,Zc��)S��ATX��Y�'�|C�T0 k� ��-��-	e2D Q%1D"Q ��D    �   �Q?�I�DT	�D�<r�-Zc��)S��C�T��[�#�|C�T0 k� ¸.��.	e2D Q%1D"Q ��D    �  �Q;�I�DT	�@�4	r�-Zc���(S��C�T��]��|C�T0 k� °/��/	e2D Q%1D"Q ��D    �  �Q7�I�DT	�8�(r�.Zc��(S��C�P ��a��|C�T0 k� ¤0��0	e2D Q%1D"Q ��D    �  �Q7�AQDT	�8�$r�.Zc��(S��C�L ��b��|C�T0 k� 0��0	e2D Q%1D"Q ��D    �  ~Q3�AQDT	�4�r�/Zc��'S��C�H ��d �|C�T0 k� Ҙ0��0	e2D Q%1D"Q ��D    �  {Q3�AQDT	�4�r�/Zc��'S��C�H ��f �|C�T0 k� Ґ1��1	e2D Q%1D"Q ��D    �  xQ/�AQDT	�0���/Zc��'S��C�D ��h �|C�T0 k� ҄1��1	e2D Q%1D"Q ��D    �  uQ+�AQDT�,���0Zc��'ボC�@ ��j �|C�T0 k� �x2�|2	e2D Q%1D"Q ��D    �  rQ+�AQDT�,� ��0Zc��&�{�C�< ��k �|C�T0 k� �p2�t2	e2D Q%1D"Q ��D    �  oa'�AQDT�(����0Z3��&�s�C�8 ��m��|C�T0 k� �h2�l2	e2D Q%1D"Q ��D    �  la'�AQDT�$����1Z3��&�k�C�4 ��o��|C�T0 k� �`3�d3	e2D Q%1D"Q ��D    � 	 ia#�AQDT�����1Z3��%S_�C�, ��r��|C�T0 k� �P3�T3	e2D Q%1D"Q ��D    � 	 fa�C�DT�����2Z3�|%SW�C�( мs��|C�T0 k� �H4�L4	e2D Q%1D"Q  ��D    � 
 c��C�DT�����2Z3�x%SO�C�$!иu��|C�T0 k� �@4�D4	e2D Q%1D"Q  ��D    � 
 `��C�@T�����2Z3�x%SG�C�!дwo��|C�T0 k� �84�<4	e2D Q%1D"Q  ��D    � 
 ]��C�@T�����3Z3�t$S?�C�!�xo��|C�T0 k� �05�45	e2D Q%1D"Q  /�D    �  Z��C�@T����|3Z3�p$S7�C�!�yo��|C�T0 k� �(4�,4	e2D Q%1D"Q  ��D    �  X��C�<T�  ��t3Z3�l$S/�C�!�{o��|C�T0 k� � 3�$3	e2D Q%1D"Q  ��D    �  V��C�8T�� ��d4Z3�d#S�C�!��}o��|C�T0 k� 4�4	e2D Q%1D"Q  ��D    �  S��C�8T�� ��\4Z3�`#S�D�!0�o��|C�T0 k� 4�4	e2D Q%1D"Q  ��D    �  Q��C�4T��!��T5Z3�\#C�D�!0����|C�T0 k�  4�4	e2D Q%1D"Q  ��D    �  N���C�0T��!��L5Z3�X#C�D�!0����|C�T0 k� �5��5	e2D Q%1D"Q  ��D    �  K���C�0T��!��D5Z3�T#B��D�!0���|C�T0 k� �5��5	e2D Q%1D"Q  ��D    �  I���E�,T��!��<5Z3�P"B�D�!0|��|C�T0 k� ��5��5	e2D Q%1D"Q  ��D    �  G��E�(T��"��46Z3�L"B�D�!0x��|C�T0 k� ��6��6	e2D Q%1D"Q  ��D    �  E��E�$T��"��,6Z3�TD"B�D�!0p~��|C�T0 k� ��6��6	e2D Q%1D"Q  ��D    �  C��E� T�"|�$6Z3�T@"BۂD�!0l~��|C�T0 k� ��5��5	e2D Q%1D"Q  ��D    �  A��E�T�"t�7Z3�T<"BӂD�"0d}��|C�T0 k� ��5��5	e2D Q%1D"Q  ��D    �  ?�׶E�T�#l�7Z3�T0!BÀD�"@X|��|C�T0 k� ��5��5	e2D Q%1D"Q  ��D    �  <�ӷE�T�#d�7Z3�T,!���CӨ"@T|��|C�T0 k� ��5��5	e2D Q%1D"Q  ��D    �  :�˸E�U�#`��8Z3�T$!���CӜ"@L{��|C�T0 k� ��5��5	e2D Q%1D"Q  ��D    �  7�ǹE�U�#\��8Z3�T !���CӐ"@Dz���|C�T0 k� ��6��6	e2D Q%1D"Q  ��D    �  5�úE�U�#X
��8Z3�T!���CӀ"@@z���|C�T0 k� ��6��6	e2D Q%1D"Q  ��D    �  3໻E��U�$T	��8Z3�D ���C�t"P8y���|C�T0 k� �6��6	e2D Q%1D"Q  ��D    �  1з�D0�U�$P	��9Z3�D ���C�h"P0x���|C�T0 k� �6��6	e2D Q%1D"Q  ��D    �  /Ч�D0�Vt$H��9Z3�D  �{�C�P"P$w���|C�T0 k� �7��7	e2D Q%1D"Q  ��D    �  ,У�D0�Wl$�D��9Z3�C� �s�C�@"Pw��|C�T0 k� �2��2	e2D Q%1D"Q  ��D    �  *Л�D0�Wd$�D�9Z3�C� �g�C�4"Pv��|C�T0 k� �.��.	e2D Q%1D"Q  ��D    �  (Г�D0�W\%�@�:Z3�C� �_�C�("Pu��|C�T0 k� �,��,	e2D Q%1D"Q  ��D    �  %Џ�D0�XT%�<�:Z3�C�!�W�C�"Pu��|C�T0 k� �*��*	e2D Q%1D"Q  ��D    �  #Ї�D0�YH%�<�:Z3�C�!�O�C�"_�t��|C�T0 k� �x(�|(	e2D Q%1D"Q  �D    �  ��D0�Y@%�8!�:Z3�C�!�C�C�"�t�
|C�T0 k� �l&�p&	e2D Q%1D"Q ��O    �  �w�D0�Z8%�8!�:Z3���!�;�C��"�s�|C�T0 k� �\%�`%	e2D Q%1D"Q ��O    �  �o�D@�Z0&�8!�:Z3���!�3�C��#�s�|C�T0 k� �P#�T#	e2D Q%1D"Q ��O    �  �k�D@�[(&�4!�:Z3���"�'�C��#�r�|C�T0 k� �@!�D!	e2D Q%1D"Q ��O    �  �[�D@�]&�7�!x:Z3�
��"��C��#�r�|C�T0 k� �$�(	e2D Q%1D"Q ��O    �  �S�D@�]�&�7�p:Z3�
Ӱ#��C��#�r�|C�T0 k� ��	e2D Q%1D"Q ��O    � ���K�EP�^�&�7�l;Z3�
Ө#��CҼ#�r��|C�T0 k� ��	e2D Q%1D"Q ��O    � ���G�EP�_��&�3�d;Z3�	Ӡ#���CҰ#�r��|C�T0 k� ��� 	e2D Q%1D"Q ��O    � ���?�EP�_��'�7�\;Z3�	Ӝ$��CҨ#�r�||C�T0 k� ����	e2D Q%1D"Q ��O    � ���7�EP�`��'�7�X;Z3�	Ӕ$��CҜ#�r�||C�T0 k� ����	e2D Q%1D"Q ��O    � ���/�EP�`��'�7�P;Z3�	ӌ$�ߐCҔ#�r�x|C�T0 k� ����	e2D Q%1D"Q ��O    � ���+�EP�a��'�7�H;Z3�ӄ%�בC҈#��r�x|C�T0 k� ����	e2D Q%1D"Q ��O    � ���#�EPxb��'�7�D;Z3��|%�ϒC�#��r�x|C�T0 k� ���	e2D Q%1D"Q ��O    � ����EPpb��'�7�<;Z3��t%�ǓC�t#��r�t|C�T0 k� ���	e2D Q%1D"Q ��O    � ����EPhc�'�;�8;Z3��l&ѿ�C�l#��s�t |C�T0 k� ���	e2D Q%1D"Q ��O    � ����EP`c�(
B;�0;Z3��d&ѳ�C�d#��s�t"|C�T0 k� ����	e2D Q%1D"Q ��O    � ����EPXd�(
B;�(;Z3��\&ѫ�C�X#��s�t#|C�T0 k� �|
��
	e2D Q%1D"Q ��O    � �����EPPe�(
B?�$;Z3��T'ѣ�C�P#�xt�t$|C�T0 k� �l	�p		e2D Q%1D"Q ��O    � �����EPHe�(
B?� <Z3��L'ћ�C�D#�pt�t%|C�T0 k� �`�d	e2D Q%1D"Q ��O    � �����E@@f�(
B?�<Z3��D'я�C�<#�ht�p&|C�T0 k� �P�T	e2D Q%1D"Q ��O    � �����E@4f�("?�<Z3��8'ч�C�0#�du�t'|C�T0 k� �D�H	e2D Q%1D"Q ��O    � �����E@,f�("?�<Z3��0(��C�(#�\u�t(|C�T0 k� �4�8	e2D Q%1D"Q ��O    � �����E@$g�t("?�<Z3��((�w�C� #Tv�t)|C�T0 k� �( �, 	e2D Q%1D"Q ��O    � �����E@g�l)"?�<Z3�� (�k�C�#Lv�t*|C�T0 k� ����	e2D Q%1D"Q ��O    � �����E@g�d)"C� �<Z3��(�c�C�$Dw�t*|C�T0 k� ����	e2D Q%1D"Q ��O    � �����E@h�\)2C� �<Z3��)�[�C� $<w�t+|C�T0 k� �����	e2D Q%1D"Q  ��O    � �����E@h�T)2C� �<Z3��)�O�C��$4x�t,|C�T0 k� ������	e2D Q%1D"Q  ��O    � ����EO�h�H)2C� �<Z3�� )�G�C��$0x�x,|C�T0 k� ������	e2D Q%1D"Q  /�O    � ����EO�h@)2C� �<Z3���)A?�C��$(yx-|C�T0 k� ������	e2D Q%1D"Q  ��O    � ����EO�h8)2C� �<Z3���*A7�C��$ yx-|C�T0 k� ������	e2D Q%1D"Q  ��O    � ����E?�h0)BC� �<Z3���*A+�C��$zx.|C�T0 k� ������	e2D Q%1D"Q  ��O    � ����E?�h$*BG�P�<Z3���*A#�C��$z|.|C�T0 k� ������	e2D Q%1D"Q  ��O    � ����E?�h*BG�P�<Z3���*A�C�${|.|C�T0 k� ������	e2D Q%1D"Q  ��O    � ����E?�g*BG�P�=Z3���*A�C�$/ {�|.|C�T0 k� ������	e2D Q%1D"Q  ��O    � ����E?�g*BK�P�=Z3���+A�C�$.�{�|/|C�T0 k� ������	e2D Q%1D"Q  ��O    � ����CO�g*BK�P�=Z3��+���D�$.�z��/|C�T0 k� �w��{�	e2D Q%1D"Q  ��O    � �|��CO�f �*RK�P�=Z3��+���D�$.�z��/|C�T0 k� �g��k�	e2D Q%1D"Q  ��O    � �x�w�CO�f �*RO�	��=Z3��+��D�$.�z��/|C�T0 k� �[��_�	e2D Q%1D"Q  ��    � �t_o�CO�e �*RO�	��=Z3��,��D�$.�y��/|C�T0 k� �O��S�	e2D Q%1D"Q  ��    � �t_k�CO�e�*RS�	��=Z3��,�ߩDx$.�y��/|C�T0 k� �C��G�	e2D Q%1D"Q  ��     � �t_[�I_�d�*RW�	��=Z3��,�˫Dd$
N�x��.|C�T0 k� �7��;�	e2D Q%1D"Q  ��     � �t_S�I_�d�+R[�	��=Z3��,�ìD\$
N�x��.|C�T0 k� �3��7�	e2D Q%1D"Q  ��     � �s_K�I_|c�+R_�	��=Z3�|-���DT$
N�x�.|C�T0 k� �+��/�	e2D Q%1D"Q  ��     � �r_C�I_tc�+R_�	��=Z3�t-���DH$
N�w�-|C�T0 k� �#��'�	e2D Q%1D"Q  ��     � �q_;�I_pc�+Rc�	��=Z3�l-���D@$
N�w�-|C�T0 k� ����	e2D Q%1D"Q  ��     � �p_3�I_hb�+Rg�	��=Z3�d-���D4$
N�v�,|C�T0 k� ����	e2D Q%1D"Q  ��     � �o_+�Iodb�+Rk�	��=Z3�\-���D,$
N�v�,|C�T0 k� ����	e2D Q%1D"Q  ��     � �no#�Io`b�+Ro�	��=Z3�T-���D $
N�uo�+|C�T0 k� ������	e2D Q%1D"Q  ��     � �mo�IoXb�+Ro�	��=Z3�L.���D$
N�uo�+|C�T0 k� ������	e2D Q%1D"Q  ��     � �lo�IoTb�|+Rs�	��=Z3�D.��D$
Nxto�*|C�T0 k� ������	e2D Q%1D"Q  ��     � �ko�IoPb�t+Rw�	��=Z3�8.�w�D$
Npso�)|C�T0 k� ������	e2D Q%1D"Q  ��     � �j^��I_Hb�d,R{�	�|=Z3�(.�g�D�$
Ndro�(|C�T0 k� ������	e2D Q%1D"Q  ��     � �h^��I_Db�\,R�	�x=Z3� .�_�D�$�`so�'|C�T0 k� ������	e2D Q%1D"Q  ��     � �f^��I_@b�P,R��	�t=Z3�/�W�D�%�\s_�&|C�T0 k� ������	e2D Q%1D"Q  ��     � �d^��I_<b�H,R��	�p=Z3�/�K�D�%�Xt_�&|C�T0 k� ������	e2D Q%1D"Q  ��     � �b^��I_8b�@,R��	�p=Z3�/�C�C��%�Xu_�%|C�T0 k� ������	e2D Q%1D"Q  ��     � �`^��Io4b�8,R��	�l=Z3� /�;�C��%�Tu_�$|C�T0 k� ������	e2D Q%1D"Q  ��     � �^^��Io0b�,,R��	�h=Z3��/�3�C�%�Pv_�$|C�T0 k� ������	e2D Q%1D"Q  ��     � �\^��Io,b�$,R��	�h=Z3���/�+�C�%�Pv_�#|C�T0 k� ������	e2D Q%1D"Q  ��     � �Z^��Io,b�,R��	�d=Z3���0�#�C�%�Lw_�"|C�T0 k� ������	e2D Q%1D"Q  ��     � �XN��Io(b�,R��	�`=Z3���0��C��%�Hw_�!|C�T0 k� ������	e2D Q%1D"Q  ��     � �VN��I_$b�,R��	�`=Z3���0��C��%�Hx_�!|C�T0 k� ������	e2D Q%1D"Q  ��     � �TN��I_$b� ,��	�\=Z3���0��C��%�Dx�| |C�T0 k� �| �� 	e2D Q%1D"Q  ��     � �RN��I_ b��,��	�X=Z3���0��C�|%�@y�| |C�T0 k� �t�x	e2D Q%1D"Q  ��     � �PN��I_ b��,��	�X=Z3��0���C�t%�@y�x|C�T0 k� �l�p	e2D Q%1D"Q  ��     � �NN��I_b��-��	�T=Z3��0���C�h%�<z�x|C�T0 k� �d�h	e2D Q%1D"Q  ��     � �L                                                                                                                                                                            � � �  �  �  f A�  �M����   �      6 \��u� ]��� �  � ^c   � �	    ��i	7     ^���h��    �� �                j  Z�8          ���    ��    0			          Z��        ���B     Z���¶    ����   	               Z�8         �0     ��   0	&
           ���Y   � �  	�Zа    �����ZR�    �f   
            
 Z�8         ��     ��    H
          T��   � �	   �*"N     S��*1.    t�                 t Z�8          � �    ��    @           j1�   � �	    1���     jb���9\    �#�P                *  Z�8          ���    ��   
8          �J ��     E �)F     �J �)F                              ����             
  ��     P5            �    	     Y��q     �k���    �s��                    �        �@     ���   @
%         ���-  $ $       m�3    ��o���    �^                   � �        �  �  ���   H

         ��a� $ $       ��v/G    ��i>�v&�    �� }                           	�     ���   0           %�  $ $       ����     %?��g     q                     A�$         	 �P     ���   	8$          ���  $ $       ���h�    �����`h    � ~                   ���$         
 f@      ���   H

          4�F ��
      ���,�     4���&     � c                  
  ���)              '  ���    		 5                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��yj  ��        ���o     ��yj��o          "                    x                j  �   �   �                             � ;;       ���   ��    ��   1     ��                                      . $        �                         �i���Z�*�� ����v�����������    
   	           
 �   a�y ��^       �$  }� �d  ~  ̄ 0f� �� g  � 0g@ �  b� �D b� ɤ  ]� �� ]����X � �$ d  �D  d@ �� d� �� 0d� �  e  �D e@ D� g  �d �f  �d g  
�\ W  
�� W@ 
�\ W` 
�< X  
�| X  
�\ X@ �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ � }����� ����� � 
�| V� 
�\ X  
�� X  
�| X@���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����8�� �� �  ������  
�fD
��L���"����D" � j  "  B   J jF��   
  �j @ b���
��
���     �j�� (*&�
� �  �  
�  .    ��     ��$  �    Z    ��     ���      ����  ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �&&      �� � �  ���        � �  ���        �        ��        �        ��        �    ��     �C�����         ��                         ��  0 	 ��	�                                      �            	 
    ����             /�& ��"�(��!   �8��               11 Kasparitis  rom v   0:01                                                                       2   5     �=�� �.�� �$c� �4 c� �$J�C<J�3%C1WC4X	C6P4 
C9_ �C:N� �� �1 � �c�c� c�cm u cu mc� c� �cY ca � �C= �C E � C#> �C$= �C&H �C	 � � K � �C � �  C � �!C � �"C � � #C � �$B�I � %B�O �&B�B �'B�J � (B�R �)k� v � *k� �G+"�?G ,"�Q7-"�;7.*�JI/"� �I 0"� �91� �92
� �X 3"N q8 4*GyX  *Ni:6
� �X 7"N q8 8*GyX  *Ni  :"D w(  "S w(  "S w(  "S w �>*'W � *7o                                                                                                                                                                                                                         � R               
     &G <     M P E k  ��        
            ����������������������������������� ���������	�
�����������                                                                                          ��   ��� �� ��������������������������������������������������������  �2, R� B ;���	��@M �@� @��@�@�� �i� ���
���/
                                                                                                                                                                                                                                                                                                        �A���
�p�                                                                                                                                                                                                                                        �  
 " )      
 ��J      �*                             �����������������������������������������������������                                                                   
                                              	                  �  ��eQ �  �  �                              	 
	 
 	 	 	 	 � ��� �� �����������  �������� ���� �������� ��������������������������� ������������������� �������������� �������������������������� ����������   � ������� ������������ �������������������  ��������������������������� �������������         n             
      3  	  = '    �� <�J      �  	                           �������������������������������������������������������                                                                                                                               �  ?� �    ?� � v                            	
  	
 	
 	
 	
 	
 ��������� ������ � ���� �������� � ���� �������������� ��������������������������������������������������������������� ��������������������������������������������� ��  �������������� �������� �������� �������� ������������ ������ ��� ��������                                                                                                                                                                                                                                                                                                               
        �              	
 
                �  }�         �#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" 8 F <                                 � �2� �\                                                                                                                                                                                                                                                                                    !�2"$  )FF                                      m                                                                                                                                                                                                                                                                                                                                                                                                                   5#   Iq� 9#  <#  $#  Cm� �#��� �  ̆ " *R ��� ������q�����q�����                       :        $   �   &  QW  �   y                    �                                                                                                                                                                                                                                                                                                                                      p K K                          !��                                                                                                                                                                                                                            \��   �� � ���      �� B  �� 
� ��� �� �����������  �������� ���� �������� ��������������������������� ������������������� �������������� �������������������������� ����������   � ������� ������������ �������������������  ��������������������������� ���������������������� ������ � ���� �������� � ���� �������������� ��������������������������������������������������������������� ��������������������������������������������� ��  �������������� �������� �������� �������� ������������ ������ ��� ��������             $�˺��˺��̻��̻��̻��̻��̻��̻�����������������������������������ww�wwU�wWU�wuu��uU��wU��wu�wwwuUuwUUUWUUUwUUUuUUUwUUUwUUWwUUwwww��www�wwx�ww�xwxx�w���wxwwwwx�����x�������x��̈������̈��̈����̻��˻��˻��˻��̻��̻��̻�f˻��������������������x˩��˩��˙���wuu�wwU�wwu�www���w���������Y��uUUUUUUUUUuUwWwwwwwx�ww��wx��UxxUwwwwwwwwwwwWwxw�����������x��{�x�̹x���x�̙w�̙��ʘ��ʨ�xň�w���˺��˺��˺��˺��˺��̺��̻��̻��������x����������w���ww��ww��ww�U�z�W�Y�Wu�wwu�wuX�wu��wx��x����wu����x���W���w������x�������x�y�X�����wwwwwuwwwwwwuwwwwww�wwWwww��wu��ww��wxw�wx��w�w�w�w�w����̻��̻���̻���˛̼˛�˼���˹�̼��ww���w���x��ww��ww���w�������x����wx��wxx��wx�xwz�wwz�xux�wwx���x���x���x���W��wW���y����w���wwwwwwwwwwuwwwWwwWuwwWUwwwwwwwwwww���w�W�x�U�x�u�x�w���x�x�������̼̻��̻���˙��˙��˙��˙��˙��̺��w���x������������������������ww���w�������w�x�w���������������wx�wWwx�wuw�������������w�����wwwwxwwwxwww�Wxxx�ww��ww�wwx�wwx������������������������������������̉��̙��̚��̚�˻�̻��̻��˻�����˺��̻���˪��̹��̺���˺��˻�x���������w�����������������������w��wwwwwx�www�ww�wwwx�ww��wxxw�x�����x�������x�������������������������������������������������$    F   '   H   &  ��                       B     �  �����J����'     ��     �� 
 	 � 
 �	  
 	  
 	  
 	  
 	 � 
 	 � 
 	� � 
 
	 � 
 	  
 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �f ��        p���� ��   p���� �$     `d ��     `d �$ ^$ �@          �� �  �� � ��  ��   �   ��  �����    �   ��    �   �$ ^$        ����          � ��� �� � ��� �$ %,  ��% ,      �  ��  ��������2����  g���  �     f ^���       ���      �      ��u����2�������J���� ��      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wenwvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                  8   �   �                    88:���������          �  90 ��  :�  ��  :�  ��  :�  ��  :�  ���������ڡ��ڡ�ّ�ک���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      �������ڡ��ڡ�ّ�ک������������������������������������������ڡ��ڡ�ّ�ک���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  ��  :�  ��  :�  ��8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0         :�  ��  :�  ��  :�  ��  :�  ���������ڡ��ڡ�ّ�ک���                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�������  :�  ��  :�  ��  :�  ��  :�  ��������������������������������������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                        ��  9�  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                  8889���������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5     9   �  �  �  �  	�  9�  9��   0                                                 �  90 ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃���������К������ڡ��ڡ�ّ�ک����  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " �������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک���DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��  �������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک����������ڡ��ڡ�ّ�ک���     	� �� �����3��3��3��33�������������3333333333333333333������������33333333333333333333������������33333333333333333333������������333=3333333333333333�   ��  ��  ��� :�� 3���3:��33����33��33��33��33��33��33��33��333333333333333�333��33���33��33:�3333333333333333333333333333�333333333333333333333333333333333333333333333333333333333333333333333��33��33��33��33��33��33��33����33��33��33��33��33��33��33��33333�333:333333333333333333333333�333��������333333333333333333333333��������333333333333333333333333��������3333333333333333333332�������߭�33��33��33��33��33����33�3	��3 �� �� 
��  �   3333333333333333����������������3333333333333333����������������3333333333333333����������������3333333333333333����������������3?��3:��3��:�� ��� ��  ��  �   wwwwwwwwwwwww}��w}��w���wDDDw��}wwwwwwwwwwww��w���G���M�DDDD��}�wwwwwwwwwwww������������DDDDGw��wwwwwwwwwwww}�ww}�Gw��GwDDGw��wwwwwwwwwwwwwwwwwwwwWwwwUGwwUTwwEUwwwwwwwwwwwwwwwwwwwwwUWUuUDU\TG\wwwwwwwwwwwwwwwwwwwwwuUwGU�GE�Dww��}}�D}}�Gt}���}���t���wDDDwwww��}���}���}������G���G��DwDDwwwwGw��Gw��G}�D���M���M���MDDDtwwww��ww��ww��ww������������DDDDwwwwwwt\www�ww|�Gw��G}�DGtDGGwwwwwww�Dw\�Gw���w�M�G�t�G�wMGDwtGwwwww��Gw�Dww�GwwDwwwGwwwwwwwwwwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "" "  """ ""   "! " ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ ""   "! " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                            " ""   "" !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                          �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                                                                                                                                                                                                                              �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �        �� ۼ�����wp���vvp�ww�             �                                ��  �                               ��  ��  ���                                                                                                                                                                                                 
���	���̜̽�˽�̈ۻ��ۻ�۽��˲"������"���" ��"                "   "   "                 ���       �   �  �  ����           �  ��� ݼ� w�� m}� ggp wz�����""H�""T�B"UJ�"UJ�@T�DT�TUJ�  ��.�                           5J� �J� �˻ �˰ ʘ� ̪ ˲"�" ""�"" �  ��                /���"/�  ��                    �                                                                            �               �  �  ��  �   �   �                         ���                                                                                                                                                                                         � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �                                                                                                                                                                                                        ۻ� ۽� ��� H�DH�D�DP�E X�T H�P H�@ Ȥ� ̻� ˘ �� "*� �/�""/""/���                       ��  ۼ� ݻ� w�� b}ذgvz�w������ɨ�ͨ���ڋ��٭���ۻݻ� �   �          �   �   .   ."  ""  ""  ,   �   
            "  "  ""  "�   �           �   ��  �      �                                     �  �  �  ��  �  �  �  ��  �             �   �   �             � � "            � "�",�"+� ",                       "  .���"    �     �                              �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                                 �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                         �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                                                                                                                                                                                                                                  �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �      �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                                                                                                                                                                                                                                      �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �   �   �"  ""  !� �� ��  �               �   ������  ��   �   �   �                                      �������  ���    �                                                                                                                                                                                                                                      �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �      �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                                                                                                                                                                                                                                      �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �      �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                                                                                                                                                                                                                                            �  ��� ��� ��� �ݪ�                       �   �    �z� 
�� ������������ ˍ� ��� ���������ˉ����� ؤ ݺD��D�؄��P �ܰ�͈��������
�� ْ �" ��"   ��                    ˚ �ȩ ݋� �۰ ˽  �˰ �˹ ̻� ˼� ��� ��D DUD TD3 D30 K�� ۻ� �ɠ ݊� �� �" �""/�!� �� /  /�� �                                         �  ��  �� ��  ���"!�����                            �  �� Ș ��  ��  �     �!� �                                                                                                                                                                                                                                       5    1  !  �� :�� � :� � :� �X     ����11��������XXXX ����111111��������31XXXX :� � :�0�
�0�	P:�
� �:� �� 
Z�  ��  ��                                                                                                                 �� ��� � � � � �� �8 ��P 
� 	 
1 	 1  �	0	�� �� 9�1 �X  �               ��������S��08�1��5� ��        ��������X8XU85858585�������X ���                                                                                                                                                                                    D@ D�D D@  �D�JJN�J��J��J��J��JJD�N�                    �   �       
    �  ��	���������                                                                                                                                                                                                                                                                                                                                                                                                                                                                               "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""��������������������""""������DDH�D��""""������D�H�H""""�������HH�H�H""""����������D�H""""������A�DA����""""�����AD�DH����""""����������D�����������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD���������������������3333DDDD����DHHDD�H����3333DDDDAHAH�H�H�D�H����3333DDDD�H������D������3333DDDD�H���DD������3333DDDD����A��A�DHD�����3333DDDD�����AA�HDD����3333DDDD���������D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""��ݙ��ٙ�ݙ��ٙݙ�ٙ�""""������MDAD��M��""""�ٙ����A�IAA""""��������A��A�A""""�������A�MAA""""�������A��A�A""""������������""""�������A��A�M""""������DD������"""$���4���4���4���4�ݙ4�ٙ4�������ݙ�ٙݙ�ٙ�333DDD���������љ��ݙ��ݙ���3333DDDDM��ݑ�A�DID����3333DDDDADA�A�A��MD����3333DDDD�A�A�A�A��MD����3333DDDDADA�A�A��MD����3333DDDD�A�AAD�DM�D����3333DDDDDD������A��DM����3333DDDD�M�M�A�AD��M����3333DDDD������D�DDM���ٙ3333DDDDݙ�4ٙ�4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  � � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�DDqwqqAtDGDwwww3333DDDD �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�wUU4uUU4UUU4UUU4UUU4UUU43334DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=""""������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����DDD�II x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx������������������333DDD w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xwwDAIAIAIA�I�I����3333DDDD  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(I�A������D�D����3333DDDD �  + � � � � � � � � � � � ��� � ��� � � � � � � � � � � � ��� � ��� �� ����(+((�""""UUUUUZ�A��A�A ` m � W � � � � ��� � ����� � ��� � � � � � ��� � ����� � ��� � ����(W(�m(`""""������������ M   a �B � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ���	B�(a((M""""�������DJD� � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�UQUDQJUDD�UZ��3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(��A���JJJ�DD�����3333DDDD 5 6  X � �F � � � � � ����� � � ������ ��� � � ����� � � � � ��	F ��(X((6(5AU4�E4E4E4DDU4UUU43334DDDD x �  l � �G � � � � � � � � � � � � ������� �� � � � � � � � � � � � ��	G ��l((�x""""�ٙ����A�IAA w w x y�������H���������������������������������H������yxww""""������������  � + w�������I�J�K�L�M�N�O � � � � � � � � � � � � � � � � � � � ��O�N�M�L�K�J�I������w(+�(�������ݙ�ٙݙ�ٙ�333DDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,�A�A�A�A��MD����3333DDDD +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+�M�M�A�AD��M����3333DDDD 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5""""����������������ݪ�� =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=""""������A�DA����M     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( """"������������������������ � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � ������������������ݪ���3333DDDD � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � �AAD�M���D�����3333DDDD ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`ݪ�4ڪ�4���4���4���4���43334DDDD M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M""""������A��AA � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�""""����DDD�II � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�����������������333DDD 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5ADA�A�A��ID����3333DDDD x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xI�A������D�D����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""��ww��ww�www�ww|www�ww|� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""wwwwwwGGqqqqD � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4ww|4ww�4w|�4��w��w�ww�wwwwwww|333DDDww��w|��w���|������w���w3333DDDD�ww��w|�ww��w|��w��w|��w3333DDDD�qD�qwwqwwqwwwDwwwww3333DDDDGGwwGwwwwtDDwwww3333DDDDqGwDwwGwwGwwtGwwwww3333DDDDDDqwqqqwAwtDGwwww3333DDDDDwGwqqwqDwtGwwww3333DDDDtwwqwwDwDDGwwwww3333DDDDwwwwwwwwwwwwwww|www�ww|�3333DDDDw��4|��4���4���4���4���43334DDDD"""UUUUUUUUUUUUUUUUUU""""UUUwUUWqUUwUWqUwWq""""wqqwQuQ""""UUUUUUQUAQQAA""""wwwwDDDwGGG""""wwwwwwwqqDqG""""wwwwwGDDGGG""""wwwwqqqAqAqAqA""""wwwwwwqAqwAwG""""wwwwwwDDwwwwww"""$www4www4www4wwu4wwU4wuU4UUUUUWUUwUWqUwWq333DDDwqwuwUuU3333DDDDwUQuUQUUQUUQUUUDUUWw3333DDDDDqTGqwwwwwwqwwwwwwww3333DDDDDGGwwGGGDDtGwwww3333DDDDqGqqqqwwDwtwwww3333DDDDqGqqwDDwtwwww3333DDDDqAqAAADDtGwwww3333DDDDwGwGwAwADwtGwwww3333DDDDtwwqwwDuDDGUwwuU3333DDDDwUU4uUU4UUU4UUU4UUU4UUU43334DDDD"""������������������""""�������������������""""��������DH�H�""""�������A�D�AI�A""""�������A��AA""""�������A��A�A""""������AD�H�""""������H�H�H�H�""""������D""""�����AADD�����"""$���4���4���4���4���4���4������������������333DDD��������������������3333DDDDH�H�H��H��I�D�����3333DDDDI�A�AAD��DH�����3333DDDDD�H�����D��H����3333DDDD�A�AAD�DDH�����3333DDDDH�����AD��A����3333DDDDH������D���3333DDDDDD���D��D����3333DDDD������ADHDDH����3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""���w���w��ww��ww�www�www""""www�wwx�ww�wx�w��x���""""�����ADDA�qq""""wwwwqwqqqD""""wwwwwwDqGq""""wwwwwwwGAD""""wwwwqqDGDDwwq""""wwwwwwwGwwDGwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4wwx4ww�4wx�4��������w��w�ww�ww333DDDwwwwwwwxwww�wwx�ww��wx��3333DDDD�����������������t���w3333DDDDAq�AAADDwDwwww3333DDDDAqDqGqGwDtGwwww3333DDDDAAAqGqGwDtGwwww3333DDDDGwDwGqGwDtGwwww3333DDDDwwAwwqqwDtDwwww3333DDDDwwwGwwGwwGwwDwwwwwww3333DDDDwwwwwwwwwwwwwwwxwww�wwx�3333DDDDw��4x��4���4���4���4���43334DDDD"""����������������""""�UU�UUUUUUUQUUUUUQ""""U��Q��������U��U""""UUQUQUQDUQ""""��������A�A���""""��������������""""������IADDA�AI""""������IDDI����""""������������������������""""������������������������"""$���4���4���4���4��4��4�U�UUUUUUUUUUQ333DDDUU�UQ�U��Q������3333DDDD�UU�UQUUUQUU�UQ�3333DDDD����������DD����3333DDDD��A�AAD�DD����3333DDDD�����I�I�DD����3333DDDDADIA��II�I�DD����3333DDDD=�� �.�� �$c� �4 c� �$J�C<J�3%C1WC4X	C6P4 
C9_ �C:N� �� �1 � �c�c� c�cm u cu mc� c� �cY ca � �C= �C E � C#> �C$= �C&H �C	 � � K � �C � �  C � �!C � �"C � � #C � �$B�I � %B�O �&B�B �'B�J � (B�R �)k� v � *k� �G+"�?G ,"�Q7-"�;7.*�JI/"� �I 0"� �91� �92
� �X 3"N q8 4*GyX  *Ni:6
� �X 7"N q8 8*GyX  *Ni  :"D w(  "S w(  "S w(  "S w �>*'W � *7o333DDDIBIBIBBBB$B�"")�3333DDDDAADA�A�ID������3333DDDDADA�IA��A��ID������3333DDDD���������I�DDI����3333DDDDDI��������DD�����3333DDDD���������I�DDI����3333DDDDDI����DD�����3333DDDDADAI�I�I�D�����3333DDDDDD��I���I��I��I��D���"3333DDDD"4�"4"4D"4DB"4"""43334DDDD"""������������������""""������������������������""""��������������������""""������DDH�D��""""������D�H�H""""�������HH�H�H��������������������������������""""�����AD�DH����""""����������D�������������������������������������������������������������������3333DDDD���������������������3333DDDD�������������� � � � � � � � � � � � � � � � � ����H������D������3333DDDD�H���DD������3333DDDD����������������p�q����f�g�y�z�������������������D���H�������3333DDDD���4���4���4���4���4���43334DDDD����������������������¤����������������""""���ݙ��ݙ��ݝ�����ݙ��ٙ""""ݙ��ٙ�ٙ�ݙ��ٙ�ݙ��ٙ�������������� �$��0�X�^�[�]�W�J�U�U��d�"�e����""""�����ADAI�I�""""��������DD������������������������.�\�\�R�\�]��K�b�(��������"""$���4���4���4���4���4���4�������������ݙ�ٙ333DDD��������������'��4�[�J�_�N�\��d� �e�������ݙ��ٙ������������������3333DDDD��A��A�I�D��DI�����3333DDDD����������������8�J�\�Y�J�[�R�]�R�\��d� �e����������D��DI������3333DDDD������������������������3333DDDD��������������������������������"""������������������""""����������A��������������������������������������""""������DHDH""""�������HA�A�A��������������������������������""""������DD�H�""""������H�DDH����������������������������������������������������D�����3333DDDDA�A�OO��O�D����3333DDDD���������������������������������AADOOOD��O����3333DDDD�A�AO�O�DO��O334CDDDD��������������������������������A���O�O�O�DD������3333DDDD���4���4���4���4���4���43334DDDD��������������������������������""""wwwwwqDDDG""""wwwwwqGAGGGG��������������������������������""""wwwwwwDGqGq""""wwwwwqGqGqGqGq��������������������������������"""$www444DD4ww4w4JJJJ�J����333DDD��������������������������������DJJJJJJJ�J�J����3333DDDD�������������D������3333DDDD��������������������������������J������DD����3333DDDDJ�������A��DJ����3333DDDD��������������������������������"""������������������""""��������������������������������������������������������""""�����������""""�����ADIA������������������������������������""""������������������������""""��������������������������� � � � � � � ������������������ � � � � � ��������������������������3333DDDD������������������������3333DDDD���@��"�(��!�����������������:�@�9���#��D�������M�DM�D����3333DDDD��A�������DD����3333DDDD��ȡɡʡˡ̡͡Τ�����������������������������������������������3333DDDD���4���4���4���4���4���43334DDDD��ϡСѡҡӡԡդ����������������B�.�;���$��""""���������������������""""������MDDA�����������������������������������""""��������A��AA""""�����DDD�M�""""�������M��DM���������""""���������������"""$���4���4���4���4���4���4wwwwwwwwwwwwwwwwww333DDDwwwwwwwwwwwwwwwwwwwwwwww3333DDDDwwwwwwwwwwwwwwwwwtwwww3333DDDDAqwAAADDwDwwww3333DDDDADAwAwAwtGDwwww3333DDDDtqwAAADDwDwwww3333DDDDDqGqqwwwqwtGwwwww3333DDDDDGwAwwwwDDtDwwww3333DDDDwwwGwwGwwGwwDwwwwwww3333DDDDwwwwwwwwwwwwwwwwwwwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""�������������������""""������ADDA����""""���������������""""�������A�IAA""""�������A��A�A""""��������A��A�A""""����DDD�II""""�������DD�""""�������I��DI���������"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDD�A���AAA�DD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�A�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDL��ALLDD�L����3333DDDDL�A������D�D����3333DDDD���L��L��L��D�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""������������������������""""������������������������""""�����������""""�����ADIA����""""�����DDD����""""��������I���I�����������""""������������������������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD������������������������3333DDDD����������������������3333DDDD�DD�M�D�������3333DDDDD�������M�DM�D����3333DDDD��A�������DD����3333DDDD����M���M���M�����������3333DDDD������������������������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            