GST@�                                                            \     �                                               �   �   ��                  � �e 
�	 J�����������x���z���        �h     #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"  ""B�j"B �����
�"    B�jl �   B ��
  ��                                                                              ����������������������������������      ��    bb QQb  114 44c c   c      		 

       	   
       ��G �   ( (                 nhp ))1         888�����������������������������������������������������������������������������������������������������������������������������o  b  o   1  +    '           �                  	  7  V  	                  �            := �����������������������������������������������������������������������������                                �X  X       4�   @  #   }   �                                                                                'w w  )n)h1p  �    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    I�;-�B޻� ltG4�f|,��!p;�[	���X��FZ3�T0 k� ����U2G�$'1e1�t B ��    � %��I�<-�B��� ltG4�g|,��!p;�[	���X��GZ3�T0 k� ����U2G�$'1e1�t B ��    � $��I�=-�B��� ltG4�g|,� "p;�[	���X��HZ3�T0 k� �'��+�U2G�$'1e1�t B  �    � #��I�>-�B��� ltG4�g|,�"pK�[	���X
��IZ3�T0 k� �7��;�U2G�$'1e1�t B ��    � "��I�?�B��� ltG4�g|,�#pK�[	.���\	��JZ3�T0 k� �C��G�U2G�$'1e1�t B ��/    � !��I�@�B��� ltG4�f|,�#pK�[	.���\��JZ3�T0 k� �S��W�U2G�$'1e1�t B ��/    �  ��F�A�B��� ltG4�f|,�$pK�[	.���\��KZ3�T0 k� �_��c�U2G�$'1e1�t B ��/    � ��F�B�B��� ltG4�f|,�$pK�[	.���`��LZ3�T0 k� �k��o�U2G�$'1e1�t B ��/    � ��F�C�B��� ltG4�f|,� %pK�[	.���`��MZ3�T0 k� �{���U2G�$'1e1�t B ��/    � ��F�D�B��� ltG4�f|,�$%pK�[ ���d��NZ3�T0 k� ������U2G�$'1e1�t B ��/    � ��F�E�E��� ltG4�f|,�,&p[�[ ���h��OZ3�T0 k� ������U2G�$'1e1�t B ��/    � ��E��F�E��� ltG4�e|,�0&p[�[ ���h��OZ3�T0 k� ������U2G�$'1e1�t B ��/    � ��E��G�E��� ltG4�e|,�4&p[�[ ���l��PZ3�T0 k� ������U2G�$'1e1�t B ��/    � ��E��H��E��� tG4�e|,�8'p[�[ ���p��QZ3�T0 k� ������U2G�$'1e1�t B ��/    � ��E��I��E��� tG4�e|,�@'p[�[����t ��RZ3�T0 k� ������U2G�$'1e1�t B ��/    � ��E��J��E��� tG[�e|,�D(p[�[����w���SZ3�T0 k� ������U2G�$'1e1�t B  ��/    �   B��K��E�� tG[�e|,�H(p[�[����{���SZ3�T0 k� ������U2G�$'1e1�t B  ��/   �  B��L��E�� tG[�e|,�P)p[�[�������TZ3�T0 k� ������U2G�$'1e1�t B  -�/    �  B��M�#�B��LtG[�e|,�T)p[�[��������UZ3�T0 k� ����U2G�$'1e1�t B  ��/    �  B��N�#�B��LtG[�e|,�X)p[�[������ UZ3�T0 k� ����U2G�$'1e1�t B  ��/    �  B��O�'�B��LtG��e|,�`*p[�[������ VZ3�T0 k� ���#�U2G�$'1e1�t B  ��/    �  B��P�+�B��LtG��e|,�d*p[�[�����WZ3�T0 k� �+��/�U2G�$'1e1�t B  ��/    �  B��Q�/�B�'�LtG��e|, �l*p[�[�����XZ3�T0 k� �7��;�U2G�$'1e1�t B ��/    �  B��R�3�B�+��tG��e|, �p+p[�[�����XZ3�T0 k� �G��K�U2G�$'1e1�t B ��/    �  B��R7�B�3��tG��e|, �x+p[�[�����YZ3�T0 k� �S��W�U2G�$'1e1�t B ��/    �  B��S7�B�;��tG��e|/���+p[�[����ZZ3�T0 k� �[��_�U2G�$'1e1�t B ��"   �  B��T?�@C��tG��e|/���,p[�[�����ZZ3�T0 k� �c��g�U2G�$'1e1�t B ��"    �  B��UC�@G��tG��e|/���,p[�[�����[Z3�T0 k� �k��o�U2G�$'1e1�t B ��"    � 
  B��VG�@O��tF��e|/���-p[�[�����[Z3�T0 k� �s��w�U2G�$'1e1�t B ��"    � 	 !B��WK�@W��tF��e|/���-p[�[�#����\Z3�T0 k� �{���U2G�$'1e1�t B ��"    �  "B��WO�@_��tFK�e|/���-p[�[�'����]Z3�T0 k� �����U2G�$'1e1�t B ��"   �  #B� XS�@g��tEK�e|/���-p[�[�+���� ]Z3�T0 k� ������U2G�$'1e1�t B ��"    �  $B�Y[�@k��tEK�e|/���.p[�[�3����$^Z3�T0 k� ������U2G�$'1e1�t B ��"    �  %B�Z�_�@s��tDK�e|/���.p[�[�7����(^Z3�T0 k� ������U2G�$'1e1�t B ��"    �  &B�Z�c�@{��tDK�e|/���.p[�[�;����,_Z3�T0 k� ������U2G�$'1e1�t B ��"    �  'B�[�k�@���tCK�e|/���/p[�[�C�����0_Z3�T0 k� ������U2G�$'1e1�t B  ��"    �  (B�\�o�@���tBK�e|/���/p[�[�G�����8`Z3�T0 k� ������U2G�$'1e1�t B  ��"    �  )B�]�s�@���tBK�d|/���0p[�[�O����<aZ3�T0 k� ������U2G�$'1e1�t B  ��"    �  *B� ]�{�@����tA��d|/���0p[�[�S����@aZ3�T0 k� ������U2G�$'1e1�t B  ��"    �   +B�$^�| @����t@��d|/���1p[�[�[����DbZ3�T0 k� ������U2G�$'1e1�t B  /�"    ��� ,B�,_݄@����t?��c|/���1p[�[�c����HbZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� -B�0_݈@����t?��c|/���2p[�[�g����PcZ3�T0 k� �˿�ϿU2G�$'1e1�t B  ��"    ��� .B�4`ݐ@����t>��c|/�� 2p[�[�o����TcZ3�T0 k� �Ӿ�׾U2G�$'1e1�t B  ��"    ��� /B�<aݔE���t=��b|/��3p[�[�w����XdZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� 0B�@aݜE���t<��b|/��3p[�[�w���\dZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� 1B�HbݠE���t;��a|/��4p[�[�{���deZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� 2B�Lb�E���t9��a!�/��4p[�[�����heZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� 3B�Tc�E���t8��`!�/��$5p[�[������peZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� 4B�\d�E���t7��`!�/��,6p[�[��� ��tfZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� 5B�`d�E���t6��_!�/��46p[�[ϗ� ��|fZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� 6B�he��E���t5��^!�/��<7p[�[ϟ� ���gZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� 7B�pe��E���t4��^!�/��D8p[�[ϧ� ���gZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� 8B�xf��E���t2��]!�/��L8p[�[ϯ� ���gZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� 9B܀f��E���t1��\!�/��T9p[�[Ϸ� #���gZ3�T0 k� ������U2G�$'1e1�t B  ��"    ��� :B܄g��E���t0��\!�/��\:p[�[Ͽ��+���gZ3�T0 k� �����U2G�$'1e1�t B  ��"    ��� ;B܌g��E���t/��[!�/��d;p[�[����3���gZ3�T0 k� ����U2G�$'1e1�t B  ��"    ��� <Bܔh��E���t.��[!�/��l;p[�[����7���hZ3�T0 k� ����U2G�$'1e1�t B  ��"    ��� =Bܜi��E����t-��Z|/��p<p[�[����?�ЬhZ3�T0 k� ����U2G�$'1e1�t B  ��"    ��� >Bܤi��E���t,� Y|/��x=p[�[����G�аhZ3�T0 k� ����U2G�$'1e1�t B  �"    ��� >Bܬj��E���t*� Y|/�M�>p[�[����O�иhZ3�T0 k� 0���U2G�$'1e1�t B  ��/    ��� >Bܴj�E���t)�X|/�M�?p[�[����S�мgZ3�T0 k� 0���U2G�$'1e1�t B ��/    ��� >B��j�E���t(�X|/�M�@p[�[����[���gZ3�T0 k� 0���U2G�$'1e1�t B ��/    ��� >B��k�E���t'�W|/�M�Ap[�[���_���gZ3�T0 k� 0���U2G�$'1e1�t B ��/    ��� >B��k�D���t&�V|/�M�Bp[�[���g���gZ3�T0 k� 0��#�U2G�$'1e1�t B ��/    ��� >B��l� D�#��t%�V|/� ��Cp[�[�� o���gZ3�T0 k� ���#�U2G�$'1e1�t B ��/    ��� >B��l�(D�+��t$�U|/� ��Dp[�[�� s���gZ3�T0 k� ���#�U2G�$'1e1�t B ��/    ��� >B��m�0D�3��t"�T|/� ��Ep[�[�'� {���fZ3�T0 k� ���#�U2G�$'1e1�t B ��/   ��� >B��m�8D�7��t!�S|/� ��Fp[�[�/� ���fZ3� T0 k� ���#�U2G�$'1e1�t B ��/    ��� >B��n@D�?��t �R!�/� ��Gp[�[�;� ����fZ3� T0 k� �#��'�U2G�$'1e1�t B ��/    ��� >B� nHD�G��t�R!�/� ��Gp[�[�C� ����eZ3��T0 k� �#��'�U2G�$'1e1�t B ��/    ��� >B�oPD�K��t� Q!�/� ��Hp[�[�K� ����eZ3��T0 k� �#��'�U2G�$'1e1�t B ��/    ��� >B�oXD�K��t�$P!�/� ��ISK�[�W�����eZ3��T0 k� �#��'�U2G�$'1e1�t B ��/    ��� >B�o`D�O��t�(O!�/� ��JSK�[�_�����dZ3��T0 k� �'��+�U2G�$'1e1�t B ��/    ��� >B�$pd E�W��t�,N!�/� ��KSK�[�g�����dZ3��T0 k� �'��+�U2G�$'1e1�t B ��/    ��� >B�,pl E�[�	�t�0M!�/� ��KSK�[�s�����cZ3��T0 k� @'��+�U2G�$'1e1�t B ��/    ��� >B�4qw�E�c�	�t�4L!�/� ��LSK�[�{����� cZ3��T0 k� @'��+�U2G�$'1e1�t B ��/    ��� >B�<q�E�g�	�t�4K!�/� ��MSK�[�������(bZ3��T0 k� @+��/�U2G�$'1e1�t B ��/    ��� >B�Dq��E�o�	�t|8J!�/� ��NSK�[�������,bZ3��T0 k� @+��/�U2G�$'1e1�t B ��/    ��� >B�Lr��E�s�	�t|<I!�/� ��NSK�[������4aZ3��T0 k� @+��/�U2G�$'1e1�t B ��/    ��� >B�Trޗ�E�{�	�t|@G|/� ��OSK�[����ñ�<`Z3��T0 k�  +��/�U2G�$'1e1�t B ��/    ��� >B�\rޟ�E��	�t|DF|/� ��PU�[����Ǳ�D`Z3��T0 k�  /��3�U2G�$'1e1�t B ��/    ��� >B�hsާ�Ep��	�t|DE|/� � QU�[����˰�H_Z3��T0 k�  /��3�U2G�$'1e1�t B ��/    ��� >B�psޯ�Ep��	�t�HD|/� �QU�[����ϰ�P^Z3��T0 k�  /��3�U2G�$'1e1�t B ��/    ��� >B�xs޷�Ep��	�t�LB|/� �RU�[����ׯ�X^Z3��T0 k�  /��3�U2G�$'1e1�t B ��/    ��� >B̀t޿�Ep��	�t�PA|/� �SU�[����ۯ�`]Z3��T0 k� 0/��3�U2G�$'1e1�t B ��/    ��� >B͈t���Ep��	�t�P@|/� �SU�[����߯�d\Z3��T0 k� 03��7�U2G�$'1e1�t B ��/    ��� >B͐t���Ep��	�t�T>|/� �TU�[������l[Z3��T0 k� 03��7�U2G�$'1e1�t B ��/    ��� >B͘u���Ep��	�t
�X=|/� �UU�[������tZZ3��T0 k� 03��7�U2G�$'1e1�t B ��/    ��� >B͠u���Ep��	�t
�\;|/� � UU�[������|ZZ3��T0 k� 03��7�U2G�$'1e1�t B ��/    ��� >Bͬu���Ep��	�t	�\:|/� �$V@�[������YZ3��T0 k� �7��;�U2G�$'1e1�t B ��/    ��� >Bʹv���Ep��	�t	�`8|/� �(V@�[�����XZ3��T0 k� �7��;�U2G�$'1e1�t B ��/    ��� >Bͼv���Ep��	�t�d7|/� �,W@�[�����WZ3��T0 k� �7��;�U2G�$'1e1�t B ��/    ��� >B��v���Ep��	�t�d5|/� �0X@�[������VZ3��T0 k� �7��;�U2G�$'1e1�t B ��/    ��� >B��w��Ep��	�t�h4|/� �4X@�[�#�����UZ3��T0 k� �;��?�U2G�$'1e1�t B ��/    ��� >B��w��Ep��	�t�l2|/� �8YB��[�+�����TZ3��T0 k� �;��?�U2G�$'1e1�t B ��/   ��� >B��w��E`Ƿ	�t�l0|/� �<YB��[�3�����SZ3��T0 k� �;��?�U2G�$'1e1�t B ��/    ��� >B��w��E`˷	�t�p/|/� �@ZB��[�;�����RZ3��T0 k� �;��?�U2G�$'1e1�t B ��/    ��� >B��x�#�E`ϸ	�t�p-|/� �DZB��[�C����QZ3��T0 k� �?��C�U2G�$'1e1�t B ��/    ��� >B��x�+�E`Ϲ	�t�t+|/� �H[B��[�K����PZ3��T0 k� �?��C�U2G�$'1e1�t B ��/    ��� >B� x�3�E`ӹ	�t�x*|/� �L\B��[�S����OZ3��T0 k� �?��C�U2G�$'1e1�t B ��/    ��� >B�y�;�E`׺	�t�x(|/� �P\B��[�W����NZ3��T0 k� �?��C�U2G�$'1e1�t B ��/    ��� >B�y�C�E`ۻ	�t�|&|/� �T]B��[�_����MZ3��T0 k� �?��C�U2G�$'1e1�t B ��/    ��� >B�y�K�E`ۼ	�t�|$|/� �X]B��[�g�����LZ3��T0 k�  C��G�U2G�$'1e1�t B ��/    ��� ?B� y�S�E`߽	�t��"|/� �\^B��[�k�����KZ3��T0 k�  C��G�U2G�$'1e1�t B  ��/    ��� ?B�(z�[�EP��t�� |/� �`^B��[�s�����JZ3��T0 k�  C��G�U2G�$'1e1�t B  ��/    ��� ?B�4z�_�EP��t��|/� �d_B��[�w�����IZ3��T0 k�  C��G�U2G�$'1e1�t B  -�/    ��� ?B�<z�g�EP��t��|/� �d_B��[�{�����HZ3��T0 k�  G��K�U2G�$'1e1�t B  ��/    ��� @B�Dz�o�EP���t��|/� �h_B��[������GZ3��T0 k� �G��K�U2G�$'1e1�t B  ��/    ��� @B�L{�w�EP���t��|/� �l`B��[ч�����FZ3��T0 k� �G��K�U2G�$'1e1�t B  ��/    ��� @B�T{��EP��Lt��|/� �p`B��[ы�����EZ3��T0 k� �G��K�U2G�$'1e1�t B  ��/    ��� @B�\{���EP��Lt�|/� �taB��[я�����DZ3��T0 k� �K��O�U2G�$'1e1�t B ��/    ��� AB�d{���E@��Lt�|/� �taB��[ѓ����� CZ3��T0 k� �K��O�U2G�$'1e1�t B ��/    ��� AB�p{���E@��Lt�|/� �xbB��[ї�����(BZ3��T0 k� �K��O�U2G�$'1e1�t B ��/    ��� AB�x|��E@��Lp�|/� �|bB��[ћ�����,AZ3��T0 k� �K��O�U2G�$'1e1�t B ��/    ��� AB��|��E@��Lp�|/� ��cB��[ћ����4@Z3��T0 k�  O��S�U2G�$'1e1�t B ��/    ��� BB��|��E@��Lp�|/� ��cB��[џ����<?Z3��T0 k�  O��S�U2G�$'1e1�t B ��/    ��� BB��|��C���Lp�|/� ��cB�[џ����D>Z3��T0 k�  O��S�U2G�$'1e1�t B ��/    ��� BB��}��C���Lp�|/� ��dB�[ѣ����H<Z3��T0 k�  O��S�U2G�$'1e1�t B ��/    ��� BB��}��C���Lpܬ|/� ��dB�[ѣ����P;Z3��T0 k�  O��S�U2G�$'1e1�t B ��/    ��� BB��}��C���Lpܰ|/� ��eB�[�����X:Z3��T0 k� �S��W�U2G�$'1e1�t B ��/    ��� CB��}��C���Lpܴ	|/� ��eB� [�����\9Z3��T0 k� �S��W�U2G�$'1e1�t B ��/    ��� CB��}��C���Lpܸ|/� ��eB�([��Pߪ�d8Z3��T0 k� �S��W�U2G�$'1e1�t B ��/    ��� CB��}��C���Lpܼ|/� ��fB�0[��P۪�l7Z3��T0 k� �S��W�U2G�$'1e1�t B ��/    ��� CB��~��C���Lp|�|/� ��fB�8[��Pש�t6Z3��T0 k� �W��[�U2G�$'1e1�t B ��/    ��� DB��~���C���Lp|�|/� ��fB�@[��Pө�x5Z3��T0 k� �W��[�U2G�$'1e1�t B  ��/    ��� DB��~���C���Lp|�|/� ��gB�L[� Pϩ�3Z3��T0 k� �W��[�U2G�$'1e1�t B  ��/    ��� DB��~���C���Lp|�|/� ��gB�T[1�P˩�2Z3��T0 k�  W��[�U2G�$'1e1�t B  ��/    ��� DB��~���C���Lp|��|/� ��hB�\[1�PǨ�1Z3��T0 k�  [��_�U2G�$'1e1�t B  ��/    ��� EB����C���Lp|��|/� ��hB�d[1�P���0Z3��T0 k�  [��_�U2G�$'1e1�t B  /�/    ��� EB� ��C���Lp|��|/� ��hB�p[1�P���/Z3��T0 k�  [��_�U2G�$'1e1�t B  ��/    ��� EB���C���Lp���|/� ��iB�x[1�P���.Z3��T0 k�  [��_�U2G�$'1e1�t B  ��/    ��� EB���C���Lp���|/� ��iB܀[1�г��,Z3��T0 k� �_��c�U2G�$'1e1�t B  ��/    ��� EB��#�C���Lp���|/� ��iB܈[1�Ы��+Z3��T0 k� �_��c�U2G�$'1e1�t B  ��/    ��� EB� �+�C��� p���|/� ��iBܔ[1�Ч��*Z3��T0 k� �_��c�U2G�$'1e1�t B  ��/    ��� EB�(��3�C��� p���|/� ��jBܜ[1�У��)Z��T0 k� �_��c�U2G�$'1e1�t B  ��/    ��� EB�4�;�C��� p|��|/� ��jBܤ[1�Л���(Z��T0 k� �_��c�U2G�$'1e1�t B  ��/    ��� EB�<�C�C��� p|��|/� ��jB��[1�����&Z��T0 k� �c��g�U2G�$'1e1�t B  ��/    ��� CB�D�K�C��� p|��|/� ��kB��[1�����%Z��T0 k� �g��k�U2G�$'1e1�t B  ��)    ��� AB�L�S�C��� p|��|/� ��kB��[A�����$Z��T0 k� �c��g�U2G�$'1e1�t B  ��)    ��� ?E�T~�[�C��� p|��|/� ��kB��[A�����#Z��T0 k� �c��g�U2G�$'1e1�t B  ��)    ��� =E�\~�_�C��� p|��|/� ��kB��[A����"Z3��T0 k� �_��c�U2G�$'1e1�t B  ��)    ��� ;E�d~�g�C��� pl��|/� ��lB��[A��{�� Z3��T0 k� �W��[�U2G�$'1e1�t B  ��)    ��� 9E�p~�o�C��� pl��|/� ��lB��[A��w��Z3��T0 k� �S��W�U2G�$'1e1�t B  ��)    ��� 7E�x}	o�C��� pm�|/� ��lB��[A��o��Z3��T0 k� �O��S�U2G�$'1e1�t B  ��)    ��� 5E��}	k�C��� pm�|/� ��lB��[A��k� Z3��T0 k� �G��K�U2G�$'1e1�t B  ��)    ��� 3E��}	k�C��� pm�|/� ��lB� [A��g�	�Z3��T0 k� �C��G�U2G�$'1e1�t B  ��)    ��� 1E��}	k�C��� pm�|/� ��lB�[A��c�	�Z3��T0 k� �?��C�U2G�$'1e1�t B  ��)    ��� /E��}	k�C��� pm�|/� ��lB�[A��[�	�Z3��T0 k� �;��?�U2G�$'1e1�t B  ��)    ��� -E��|	 k�C��� pm�|/� ��lB�[A|�W�	�Z3��T0 k� �3��7�U2G�$'1e1�t B  ��)    ��� +E��|	 k�C��� pm�|/� ��lB� [Qx�S�	�Z3��T0 k� �/��3�U2G�$'1e1�t B  ��)    ��� )E��|	 k�C��� pm�|/� ��lB�,[Qt�O�	� Z3��T0 k� �+��/�U2G�$'1e1�t B  ��)    ��� 'E��{	 k�C��� pm�|/��lB�4[Qp�K�
$Z3��T0 k� �'��+�U2G�$'1e1�t B  ��)    ��� %E��{	 k�C��� pm�|/��lB�<[Ql�C�
,Z3��T0 k� �#��'�U2G�$'1e1�t B  ��)    ��� #E��{	k�C��� pm�|/��lB�H[Qh�?�
0Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� !E��z	k�C��� p]�|/��lB�P[Qd�;�
4Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E��z	k�C��� p]�|/��lB�X[Q`�7�
8Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E��z	k�C��� p]�|/�^�lB�`[Q\�3�	�<Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E��y	k�C��� p]�|/�^�lB�l[QT�/�	�@Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E��y	 k�C��� p]�|/�^�lB�t[QP�'�	�@b���T0 k� ����U2G�$'1e1�t B  ��)    ��� E� x	 k�C��� p]�|/�^�lB�|[�L�#�	�Db���T0 k� ����U2G�$'1e1�t B  ��)    ��� E�x	 k�C��� p]�|/�^�lB̈́[�D��	�Hb���T0 k� ������U2G�$'1e1�t B  ��)    ��� E�w	 k�C��� p]�|/�^�lB͐[�@ ��
Lb���T0 k� ������U2G�$'1e1�t B  ��)    ��� E�v	 k�C��� p]�|/���lB͘[�8 ��
Lb���T0 k� �����U2G�$'1e1�t B  ��)    ��� 
E� v�k�C��� p]�|/���lB͠[�4 ��
Pb���T0 k� ����U2G�$'1e1�t B  ��)    ��� E�(u�o�C��� p]�|/���lBͨ[�, ��
Pb���T0 k� ����U2G�$'1e1�t B  �)    ��� E�0t�o�C����p��|/���l@�[Q+���
Tb���T0 k� ����U2G�$'1e1�t B  �)    ��� E�4s�o�C����p��|/���l@�[Q#���CTb���T0 k� ����U2G�$'1e1�t B  ��)    ��� E�<s�o�C����p��|/���l@�[Q���CXb���T0 k� �ߋ��U2G�$'1e1�t B  ��)    ��� E�Dr�o�C����p��|/���l@�[Q����C\b���T0 k� �ۋ�ߋU2G�$'1e1�t B  ��)    ��� E�Lq�o�EЇ��t���|/���l@�[Q����C\Z3��T0 k� �׊�ۊU2G�$'1e1�t B  ��)   ��� E�Tp�o�EЃ��t���|/���l@�[Q����C`Z3��T0 k� �׊�ۊU2G�$'1e1�t B  ��)    ��� C@Xo�o�EЃ��t���|/���l@�[Q����C`Z3��T0 k� �Ӊ�׉U2G�$'1e1�t B  ��)    ��� C@`m�o�E���x���|/���l@�[Q���CdZ3��T0 k� �ω�ӉU2G�$'1e1�t B  ��)    ��� C@hl�o�E���x���|/���l@�[P����CdZ3��T0 k� �ˈ�ψU2G�$'1e1�t B  ��)    ��� C@lk�o�E�{��|��|/���l@ [P����CdZ3��T0 k� �ǈ�ˈU2G�$'1e1�t B  ��)    ��� C@tj�o�E�{��|��|/���l@[P����ChZ3��T0 k� �Ç�ǇU2G�$'1e1�t B  ��)    ��� C@|i�o�E�w�����|/���l@[P����ChZ3��T0 k� ����ÇU2G�$'1e1�t B  ��)    ��� C@�g�o�E�s�����|/���l@[P����ClZ3��T0 k� ����ÇU2G�$'1e1�t B  ��)    ��� C@�f�o�E�o�����|/���l@$[P���ߑClZ3��T0 k� ������U2G�$'1e1�t B  ��)    ��� C@�d�o�C�k�����|/���l@,[P���ۑCpZ3��T0 k� ������U2G�$'1e1�t B  ��)    ��� C@�c�o�C�g�����|/���l@4[P���אCpbs��T0 k� ������U2G�$'1e1�t B  ��)    ��� C@�a�o�C�c�����|/���l@<[P���אCtbs��T0 k� ������U2G�$'1e1�t B  ��)    ��� C@�`�o�C�c����ߝ|/���l@D[P���ӐCtbs��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�^�o�C�_����ۛ|/���l@P[P���ϏCtbs��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�]�o�E�[����ۙ|/���l@X[P���ˏCxbs��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�[�o�E�W����ח|/���l@`[P���ˏCx
bs��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�Y o�E�S���ו|/���l@h[P���ǎC|
bs��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�X o�E�G���ӓ|/���l@p[P���ÎC|
bs��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�V o�E�?�̬ӑ|/���l@x[P���ÍC|
bs��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�T o�C�3�̰ӏ|/���l@�[P�����C�
bs��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�S o�C�'�̴ύ|/���l@�[P�����C�
bs��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�Q �o�C��̸ϋ|/���l@�[P�����C�	Z3��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�O �o�C��̼ψ|/���l@�[P�����C�	Z3��T0 k� ������U2G�$'1e1�t B  ��)    ��� CP�M �o�C����ˆ|/���l@�[P�����C�	Z3��T0 k� ������U2G�$'1e1�t B  ��)    ��� C`�L �o�C�����ˇ|/���l@�[P�����C�	Z3��T0 k� ������U2G�$'1e1�t B  ��)    ��� C`�J �o�C������ˇ|/���l@�[P�����C�	Z3��T0 k� ������U2G�$'1e1�t B  ��)    ��� C`�H �o�C�����ˈ|/���l@�[P�����C�	Z3��T0 k� ������U2G�$'1e1�t B  ��)    ��� C`�F o�C�����ˈ|/���l@�[P�����C�	Z3��T0 k� ������U2G�$'1e1�t B  ��)    ��� C`�D o�C�۩���ˉ|/���l@�[P�����C�Z3��T0 k� ������U2G�$'1e1�t B  ��)    ��� C`�C o�C�ϩ���ˉ|/���l@�[P�����C�Z3��T0 k� ������U2G�$'1e1�t B  ��)    ��� C`�A o�C�ǩ���ˊ|/���l@�[P�����C�Z3��T0 k� ������U2G�$'1e1�t B  ��)    ��� E� ? o�C߿����ϊ|/���l@�[P�����C�Z3��T0 k� ���U2G�$'1e1�t B  ��)    ��� E�=Po�C߷����ϋ|/���l@�[P����C�Z3��T0 k� ���U2G�$'1e1�t B  ��)    ��� E�;Po�C߯�� �ϋ|/���l@�[P{����C�Z3��T0 k� �{�U2G�$'1e1�t B  ��)    ��� E�9Po�Cߣ��ό|/���l@�[Pw����C�Z3��T0 k� �{�U2G�$'1e1�t B  ��)    ��� E�7Po�Cߛ��ӌ|/���l@[Ps����C�Z3��T0 k� �w~�{~U2G�$'1e1�t B  ��)    ��� E�5Pk�Cߓ��Ӎ|/���l@[Po����C�Z3��T0 k� �w~�{~U2G�$'1e1�t B  ��)    ��� E�4�k�Cߋ��׍|/���l@[Po����C�Z3��T0 k� �s~�w~U2G�$'1e1�t B  ��)    ��� E�2�k�C߃� �׍|/���l@ [Pk����C�Z3��T0 k� �s}�w}U2G�$'1e1�t B  ��)    ��� E� 0�g�C�{�(�ێ|/���l@([Pg����C�Z3��T0 k� �o~�s~U2G�$'1e1�t B  ��)    ��� E�$.�g�C�s�0�ߎ|/���l@0[Pc����C�Z3��T0 k� �o}�s}U2G�$'1e1�t B  ��)    ��� E�$,�c�C�o��8�ߏ|/���l@8[Pc����C�Z3��T0 k� �k}�o}U2G�$'1e1�t B  ��)    ��� E�(*�c�C�g��@��|/���l@@[P_����C�Z3��T0 k� �k}�o}U2G�$'1e1�t B  ��)    ��� E�,(�_�E__��H��|/���l@H[P[����C�Z3��T0 k� �g}�k}U2G�$'1e1�t B  ��)    ��� C�0&_�E_W��P��|/���l@P[PW����C�Z3��T0 k� �g}�k}U2G�$'1e1�t B  ��)    ��� C�0$[�E_O��T��|/���l@X[PW����C�Z3��T0 k� �c}�g}U2G�$'1e1�t B  ��)    ��� C�4"[�E_G��\��|/���l@`[PS����C�Z3��T0 k� �c}�g}U2G�$'1e1�t B  ��)    ��� C�4 W�E_?��d��|/���l@h[PO����C�Z3��T0 k� �_}�c}U2G�$'1e1�t B  ��)    ��� C�8W�E_7��l���|/���l@p[PO���C�Z3��T0 k� �_}�c}U2G�$'1e1�t B  ��)    ��� C�8S�E_/��t���|/���l@x[PK���C�Z3��T0 k� �_}�c}U2G�$'1e1�t B  ��)   ��� C�8S�E_'��|���|/���l@�[PG���C�Z3��T0 k� �[|�_|U2G�$'1e1�t B  ��)    ��� C�8S�E_�݄ ��|/���l@�[PG��{�C�Z3��T0 k� �[}�_}U2G�$'1e1�t B  ��)    ��� C�<O�E_�݈ ��|/���l@�[PC��{�C�Z3��T0 k� �W}�[}U2G�$'1e1�t B  ��)    ��� C�<O�A_�ݐ ��|/���l@�[PC��w�C�Z3��T0 k� �W|�[|U2G�$'1e1�t B  ��)   ��� C�<K�A_�ݛ���|/���l@�[P?��w�C�Z3��T0 k� �W|�[|U2G�$'1e1�t B  ��)    ��� C�<K�A^��ݣ���|/���l@�[P;��w�C�Z3��T0 k� �S{�W{U2G�$'1e1�t B  ��)    ��� C�<G�A^��ݫ���|/���l@�[P;��s�C�Z3��T0 k� �S|�W|U2G�$'1e1�t B  ��)    ��� C�<G�A^�ݳ���|/���l@�[P7��s�C�Z3��T0 k� �S|�W|U2G�$'1e1�t B  ��)    ��� L�<	 G�A^�ݷ��#�|/���l@�[P7��s�C�Z3��T0 k� �O{�S{U2G�$'1e1�t B  ��)    ��� L�< C�A^ߣݿ��+�|/���l@�[P3��o�C�Z3��T0 k� �O{�S{U2G�$'1e1�t B  ��)    ��� L�@ C�A^ۣ����/�|/���l@�[P3��o�C�Z3��T0 k� �K{�O{U2G�$'1e1�t B  ��)    ��� L�@ ?�A^ӣ����7�|/���l@�[P/��o�C�Z3��T0 k� �K{�O{U2G�$'1e1�t B  ��)    ��� L�@ ?�A^ˣ����;�|/���l@�[P+��k�C�Z3��T0 k� �K{�O{U2G�$'1e1�t B  ��)    ��� L�@  ?�A^ã����?�|/���l@�[P+��k�C�Z3��T0 k� �G{�K{U2G�$'1e1�t B  ��)    ��� L�C� ;�A^������G�|/���l@�[P'��k�C�Z3��T0 k� �Gz�KzU2G�$'1e1�t B  ��)    ��� MC� ;�A^������K�|/���l@�[P'��g�C�Z3��T0 k� �Gz�KzU2G�$'1e1�t B  ��)   ��� MC� ;�A^������S�|/���l@�[P#��g�C�Z3��T0 k� �Gz�KzU2G�$'1e1�t B  ��)    ��� MC� 7�A^������[�|/���l@[P#��g�C�Z3��T0 k� �Cz�GzU2G�$'1e1�t B  ��)   ��� MC� 7�A^������_�|/���l@[P��c�C�Z3��T0 k� �Cz�GzU2G�$'1e1�t B  ��)   ��� MC� 7�A^�����g�|/���l@[P��c�C�Z3��T0 k� �Cz�GzU2G�$'1e1�t B  ��)    ��� MG� 3�A^�����k�|/���l@[P��c�C�Z3��T0 k� �?y�CyU2G�$'1e1�t B  ��)    ��� MG� 3�A^�����s�|/���l@$[P��_�C�Z3��T0 k� �?y�CyU2G�$'1e1�t B  ��)    ��� MG� 3�A^�����{�|/���l@,[P��_�C�Z3��T0 k� �?y�CyU2G�$'1e1�t B  ��)   ��� MG� /�A^���#����|/���l@4[P��_�C�Z3��T0 k� �;y�?yU2G�$'1e1�t B  ��)    ��� L�G� /�A^��+����|/���l@<[P��_�C�Z3��T0 k� �;y�?yU2G�$'1e1�t B  ��)    ��� L�G� /�A^{��3����|/���l@@[P��[�C�Z3��T0 k� �;z�?zU2G�$'1e1�t B  ��)    ��� L�G� +�A^s��7����|/���l@H[P��[�C�Z3��T0 k� �;z�?zU2G�$'1e1�t B  ��)    ��� L�G� +�A^o��?����|/���l@P[P��[�C�Z3��T0 k� �7z�;zU2G�$'1e1�t B  ��)    ��� L�G� +�A^k��G����|/���l@X[P��[�C�Z3��T0 k� �7z�;zU2G�$'1e1�t B  ��)    ��� L�G� +�A^c�~K����|/���l@`[P��W�C�Z3��T0 k� �7z�;zU2G�$'1e1�t B  ��)    ��� L�G� '�A^_�~S����|/���l@h[P��W�C�Z3��T0 k� �7{�;{U2G�$'1e1�t B  ��)    ��� L�K� '�A^[�~[����|/���l@p[P��W�C�Z3��T0 k� �3{�7{U2G�$'1e1�t B  ��)    ��� L�K� '�A^S�~_��Ú|/���l@x[P��W�C�Z3��T0 k� �3{�7{U2G�$'1e1�t B  ��)    ��� C�K� '�A^O�~g��˛|/���l@�[P��S�C�Z3��T0 k� �3{�7{U2G�$'1e1�t B  ��)    ��� C�K� #�LK�~k��ӛ|/���l@�[P��S�C�Z3��T0 k� �3|�7|U2G�$'1e1�t B  ��)    ��� C�K� #�LG�~s��ۛ|/���l@�[P��S�C�Z3��T0 k� �/|�3|U2G�$'1e1�t B  ��)    ��� C�K� #�LC�~w��ߛ|/���l@�[P��S�C�Z3��T0 k� �/|�3|U2G�$'1e1�t B  ��)    ��� C�K� #�L;�~���|/���l@�[P��O�C�Z3��T0 k� �/|�3|U2G�$'1e1�t B  ��)    ��� L�K� �L7�~����|/���l@�[_���O�C�Z3��T0 k� �/|�3|U2G�$'1e1�t B  ��)    ��� L�K� �L3�~����|/���l@�[_���O�C�Z3��T0 k� �+}�/}U2G�$'1e1�t B  ��)    ��� L�K� �L3�������|/���l@�[_���O�C�Z3��T0 k� �+}�/}U2G�$'1e1�t B  ��)    ��� L�K� �L3�������|/���l@�[_���K�C�Z3��T0 k� �+}�/}U2G�$'1e1�t B  ��)    ��� L�K� �L7�������|/���l@�[_���K�C�Z3��T0 k� �+}�/}U2G�$'1e1�t B  ��)    ��� L�K� �L7�������|/���l@�[_���K�C�Z3��T0 k� �+}�/}U2G�$'1e1�t B  ��)    ��� MK� �L7�������|/���l@�[_���K�C�Z3��T0 k� �'~�+~U2G�$'1e1�t B  ��)    ��� MK� �L;�������|/���l@�[_���K�C�Z3��T0 k� �'~�+~U2G�$'1e1�t B  ��)    ��� MK� �L;�������|/���l@�[_���G�C�Z3��T0 k� �'~�+~U2G�$'1e1�t B  ��)    ��� MK� �L;������|/���l@�[_���G�C�Z3��T0 k� �'~�+~U2G�$'1e1�t B  ��)    ��� MK� �L.?������|/���l@�[_���G�C�Z3��T0 k� �'~�+~U2G�$'1e1�t B  ��)    ��� MK��L.?������|/���l@�[_���G�C�Z3��T0 k� �#~�'~U2G�$'1e1�t B  ��)    ��� MK��L.?������|/���l@�[_���G�C�Z3��T0 k� �#�'U2G�$'1e1�t B  ��)    ��� MK��L.C������|/���l@[_���G�C�Z3��T0 k� �#�'U2G�$'1e1�t B  ��)    ��� MK��L.C������|/���l@[_���C�C�Z3��T0 k� �#�'U2G�$'1e1�t B  ��)    ��� L�K��L.C������|/���l@[_���C�C�Z3��T0 k� �#�'U2G�$'1e1�t B  ��)    ��� L�K��L.C������|/���l@[_���C�C�Z3��T0 k� �#�'U2G�$'1e1�t B  ��)    ��� L�K��L.G������|/���l@ [_���C�C�Z3��T0 k� ��#U2G�$'1e1�t B  ��)    ��� L�K��L.G������|/���l@([_���C�C�Z3��T0 k� ���#�U2G�$'1e1�t B  ��)    ��� L�K��L.G������|/���l@,[_���C�C�Z3��T0 k� ���#�U2G�$'1e1�t B  ��)    ��� L�K��L.K������|/���l@4[_���?�C�Z3��T0 k� ���#�U2G�$'1e1�t B  ��)    ��� L�K��L.K������|/���l@<[_���?�C�Z3��T0 k� ���#�U2G�$'1e1�t B  ��)    ��� L�K��L.K������|/���l@D[_���?�C�Z3��T0 k� ���#�U2G�$'1e1�t B  ��)    ��� L�K��L.K������|/���l@L[_���?�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�K��L.O������|/���l@P[_���?�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�K��L.O������|/���l@X[_���?�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�K��L.O������|/���l@`[_���?�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�K��L.O������|/���l@h[_���;�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�K��L.S�����|/���l@l[_���;�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�K��L.S�����|/���l@t[_���;�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�G��L.S�����|/���l@|[_���;�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�G��L.S�����|/���l@�[_���;�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�G� �L.S����#�|/���l@�[_���;�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�C� �L.W����#�|/���l@�[_���;�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�C� �L.W����#�|/���l@�[_���7�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�?� �L.W����#�|/���l@�[_���7�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�?� �L.W����'�|/���l@�[_���7�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�;� �L.W��#��'�|/���l@�[_���7�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�;� �L.[��'��'�|/���l@�[_���7�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�7� �L.[��+��'�|/���l@�[_���7�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�3� �L.[��+��+�|/���l@�[_���7�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�3� �L.[��/��+�|/���l@�[_���7�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�/� �L.[��3��+�|/���l@�[_���7�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�+� �L._�7��+�|/���l@�[_���3�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�'� �L._�7��/�|/���l@�[_���3�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�'� �L._�;��/�|/���l@�[_���3�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�#� �L._�?��/�|/���l@�[_���3�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�� �L._�?��/�|/���l@�[_���3�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�� �L.c�C��3�|/���l@�[_���3�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�� �L.c��G��3�|/���l@ [_���3�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�� �L.c��G��3�|/���l@[_���3�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�� �Lc��K��3�|/���l@[_���3�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�� �Lc��S��7�|/���l@[_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C��� �Lg��W��7�|/���l@ [_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C��� �Lg��[��7�|/���l@([_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�� �Lg��[��;�|/���l@,[_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C��/��A^g��_��;�|/���l@4[_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C��/��A^g��c��?�|/���l@<[_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�ߕ/��A^g��g��?�|/���l@@[_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�۔/��A^g��k��?�|/���l@H[_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� C�ӓ/��A^k��o��C�|/���l@P[_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�ϒ/��A^k��s��C�!�/���l@T[_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�Ǒ/��A^k��w��C�!�/���l@\[_���/�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� Eп�/��A^k����G�!�/���l@d[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� Eл�/��A^k����G�!�/���l@h[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� Eг�/��A^k����G�!�/���l@p[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� EЫ�/��A^k����K�!�/���l@x[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� EУ�/��A^o����K�!�/���l@|[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E���/��A^o����K�!�/���l@�[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E���/��A^o����O�!�/���l@�[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E���/��A^o����O�!�/���l@�[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E���/��A^o�����O�!�/���l@�[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E����A^o�����S�|/���l@�[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�w���A^o�����S�|/���l@�[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�o���A^o�����S�|/���l@�[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�g���A^s�����W�|/���l@�[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�_���A^s�����W�|/���l@�[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�W���A^s�����W�|/���l@�[_���+�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�O���A^s�����[�|/���l@�[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�G���A^s�����[�|/���l@�[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�?�_��A^s�����[�|/���l@�[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�7�_��A^s��۾�[�|/���l@�[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�/�_��A^s�߽�_�|/���l@�[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�'�_��A^s���_�!�/���l@�[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E��_��A^w���_�!�/���l@�[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E��_��A^w���_�!�/���l@�[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E��_��A^w����c�!�/���l@�[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E����A^w�	����c�!�/���l@�[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E����A^w�	���c�!�/���l@[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E�����A^w�	���c�!�/���l@[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� E����A^w�	���g�!�/���l@[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� F���A^w�	���g�!�/���l@[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� F���A^w�	���g�!�/���l@[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� F���A^w�
 ��g�!�/���l@$[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� Fۇ��A^{�
 ��k�|/���l@([_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� F׈��A^{�
 ��k�|/���l@0[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� Fψ��A^{�
 #��k�|/���l@4[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� Fˉ��A^{�
 '��k�|/���l@<[_���'�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)    ��� D�Ǌ��A^{�	�+��k�|/���l@@[_���#�C�Z3��T0 k� ����U2G�$'1e1�t B  ��)   ��� Cޘ#�I�01�4#	�?��(ݠ_C�Q>���p,�(bs�T0 k� �x\�|\U2G�$'1e1�t B  ��    � 7�8Cތ�I�,1�4#	�7��(ݘ_C�R>���l-�$bs�T0 k� �p\�t\U2G�$'1e1�t B  ��    � 7�8Cބ�I�,1�0$	�3��(�_C�R>��d-�bs�T0 k� �lW�pWU2G�$'1e1�t B  ��    � 7�8C�|�I�(2�0$	�/��(�_C�S>��`.�bs�T0 k� �dS�hSU2G�$'1e1�t B  ��    � 7�8C�t��I�$2�,%	�+��(�_C�T>��X.�bs�T0 k� �\P�`PU2G�$'1e1�t B  ��    � 7�8C�h ���I�$2�,&	�'��(�x_C�|U>��P/�bs�T0 k� �TN�XNU2G�$'1e1�t B  ��    � 7�8C�X ��I�2�$'	���(�h_C�lV>��D/� bs�T0 k� �DM�HMU2G�$'1e1�t B  ��    � 7�8C�P �ߑE^3�$(	���$�`_C�dW>��<0�bs�T0 k� �<L�@LU2G�$'1e1�t B  ��    � 7�8C�H �בE^3� )	���$�X_C�\X>��40�bs�T0 k� �4J�8JU2G�$'1e1�t B  ��    � 7�8C�@ �ϐE^3� *	���$�P_C�TY>��,1�bs�T0 k� �,I�0IU2G�$'1e1�t B  ��    � 7�8C�8 �ǐE^3�+	���$�H_C�LY>��$1�Z3�T0 k� �$I�(IU2G�$'1e1�t B  ��    � 7�8C�0 ﻐE^3�+	���$�@_C�@Z>��1�Z3�T0 k� �I� IU2G�$'1e1�t B  ��    � 7�8A^$ ﳏE^3�,	��� �8_C�8[>��2�Z3�T0 k� � I�$IU2G�$'1e1�t B  ��    � 7�8A^ EN4�.	��� �(^C�(\>��3�Z3�T0 k� �H� HU2G�$'1e1�t B  ��    � 7�8A^ EN 4�0	��� � ^C� ]>���3�Z3�T0 k� �H� HU2G�$'1e1�t B  ��    � 7�8A^ ���EM�4�1	��� �]C�^>���3�Z3�T0 k� �G�GU2G�$'1e1�t B  ��    � 7�8A]� ���EM�4�2	��� ]C�^>����4�Z3�T0 k� �F�FU2G�$'1e1�t B  ��    � 7�8A]� ���EM�3�3	��� \C�_>����4�Z3�T0 k� �E�EU2G�$'1e1�t B  ��    � 7�8A]� �w�EM�3�4	����  \C� `>����4�Z3�T0 k� ��E� EU2G�$'1e1�t B  ��    � 7�8A]� �o�EM�3� 5	���� �[C��`>����5�Z3�T0 k� ��D��DU2G�$'1e1�t B  ��    � 7�8A]� �_�EM�3��7	���� �ZD�b>����5� b��T0 k� ��C��CU2G�$'1e1�t B  ��    � 7�8A]� �W�E=�2��9	���� �YD�b>��Ѹ6� b��T0 k� ��B��BU2G�$'1e1�t B  ��    � 7�8A]� �O�E=�2��:	���� �XD�c>��Ѱ6� b��T0 k� ��A��AU2G�$'1e1�t B  ��    � 7�8A]� �G�E=�1��;	�����WD�c>��Ѩ6x b��T0 k� ��@��@U2G�$'1e1�t B  ��    � 7�8A]� �?�E=�1��<	�����VD�d>��Ѡ7p b��T0 k� ��=��=U2G�$'1e1�t B  �    � 7�9A]� +�E=�0��>������TD�e>��ѐ7` b��T0 k� ��5��5U2G�$'1e1�t B  ��    � 7�:A]� #�E=�/��?������SD�f>��ш8�X!b��T0 k� ��2��2U2G�$'1e1�t B  ��    � 7�;A]� �E=�.��@������SD�f>��р8�P!b��T0 k� � .�.U2G�$'1e1�t B  ��    � 7�<A]� �E=�.��A������RD�g>���x8�H!b��T0 k� �+�+U2G�$'1e1�t B ��    � 7�=A]� �E=�-��B������QD�gN���p9�@!Z3�T0 k� �'�'U2G�$'1e1�t B ��    � 7�>A]���E=�,��C������QD�hN���h9�8!Z3�T0 k� �#� #U2G�$'1e1�t B ��    � 7�?I�����E-�+��C������QD|hN���`9�0!Z3�T0 k� �$ �( U2G�$'1e1�t B ��    � 7�@I�{��E-�)�C���|��QDliN���L:� !Z3�T0 k� �4�8U2G�$'1e1�t B ��    � 7�AI�w�ߊE-�(�C���|��PE]djΏ��D:�"Z3�T0 k� �@�DU2G�$'1e1�t B ��    � 7�BI�s�׉E-�'�C���| ��PE]\j΋��<:�"Z3�T0 k� �H�LU2G�$'1e1�t B ��    � 7�CI�k�ωE-�&	��CL� | �|PE]Tk΋��4:�"Z3�T0 k� �P�TU2G�$'1e1�t B  ��    � 6�DI�c���E-�$	��CL�| �pPE]@l·��$;��"Z3�T0 k� �d�hU2G�$'1e1�t B  ��    � 5�CI�_���E-�#	��CL�|$�hPE]8lރ��;��"Z3�T0 k� �`�dU2G�$'1e1�t B  ��     � 4�BI�[�^��E-�"	��CL�|$
�`OE]0mރ��<��"Z3�T0 k� �P�TU2G�$'1e1�t B  ��     � 3�AI�S�^��E-�!	��CL�|$	�XOE](m���<��"Z3�T0 k� �D�HU2G�$'1e1�t B  ��     � 2�@I�O�^��E-�	̘C<�|(�TOE] n���<��"Z3�T0 k� �8�<U2G�$'1e1�t B  ��     � 1�?E�G�^��E�	̐C<�|(�HOE]o^{���=��#Z3�T0 k� �,�0U2G�$'1e1�t B  ��     � 0�>E�C�^��E�	̐C<�|(�@OE]o^{���=��#Z3�T0 k� �$�(U2G�$'1e1�t B  ��     � /�=E�?�^{�E�	̌C<�|,�8NEL�p^{���=�#Z3�T0 k� �� U2G�$'1e1�t B  ��     � .�<E�;�^s�E�	��C<�|,�4NEL�p^w���=�#Z3�T0 k� ��U2G�$'1e1�t B  ��     � -�;E�3�^k�E�	��C��|,�,NEL�p^w���=�#Z3�T0 k� ��U2G�$'1e1�t B  ��     � ,�:E�+�^W�B��	��C��	|,� NEL�q^w���>�#Z3�T0 k� ��U2G�$'1e1�t B  ��     � +�9E�#�NO�B��	��C��|0�NE��q^w��>�#Z3�T0 k� ��U2G�$'1e1�t B  ��     � *�8E� NG�B��	̀C��|0�NE��r^w��>�#Z3�T0 k� ��� U2G�$'1e1�t B  ��     � )�8E� N?�B��	�|C��|0�ME��r^w��>�$Z3�T0 k� ��
��
U2G�$'1e1�t B  ��     � (�8E� N7�B��	�|C̴|0�MEܸr^w��>x$Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E� N/�B��	�xC̴|0�MEܰr�w�0�=l$Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E�� N�B��	�xC̬|0��MEܜs�w�0�=\$Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��N�B��	�xC̨|0��MEܔs�w�0|=T$Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��N�B��	�tC̨|0��LE܌t�w�0t=L$Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��N�B��	�tC̤|0��LE܄t�w�0l=D$Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��M��B��	�tC̠|0��LE�xt�w�0d<<$Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��=�B��
	�tC̜|0��KE�pt�w��\<4$Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��=�B��	�tC̘|0��JE�`u�w��L<$%Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��=ۉB��	�tC̔|0��IE�XuNw��D;%Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��=ӉB��	�tCܐ|0��IE�PvNw��<;%Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��=ˊB��	�tC܌|0��HE�DuNw��0;A%Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��=ÊB��	�tC܈|0��GE�<tNw��(:A%Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��=��B͸�tC�|"|0�FE�,s w��9@�&Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��=��B���tC�x#|0�ED<$r w��9@�&Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��	=��B���tC�t$|0�DD<r w��8@�&Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��
=��B���tC�p&|0�CD<q w�� 8@�&Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��=��B�� �tC�l'|0�BD<p {���7@�'Z3�T0 k� ����U2G�$'1e1�t B  ��     � (�8E��-��B���\tCL`*|0	�@E��o�{���6@�'Z3�T0 k� ��"��"U2G�$'1e1�t B  ��     � (�8E�x-��B���\tCL\+�,	�?E��n����5@�(Z3�T0 k� ��#��#U2G�$'1e1�t B  ��     � (�8E�t-{�B���\tCLX,�,
�>E��m����4@�(Z3�T0 k� ��$��$U2G�$'1e1�t B  ��     � (�8Fl-w�B���\tCLP.�,
�<E��k�����40�(Z3�T0 k� ��$��$U2G�$'1e1�t B  ��     � (�8F`-k�B���tCLH1�,
�:A��i�����20�)Z3�T0 k� ��%��%U2G�$'1e1�t B  ��     � (�8F\-c�B���tC�@2�,
�9A��g�����10�*Z3�T0 k� ��&��&U2G�$'1e1�t B  ��     � (�8FX-_�B��tC�<4�,�8A��f�����00�*Z3�T0 k� ��&��&U2G�$'1e1�t B  ��     � (�8FT-[�B��tC�45�,�6A��e����/0�+Z3�T0 k� ��%��%U2G�$'1e1�t B  �     � (�?H�L�S�B��tC�(8�(�4E��c����-0t,Z3�T0 k� ��"��"U2G�$'1e1�t B ��    � (�FH�H�O�B�� �tC�$:�(�3E��b����+0p-Z3�T0 k� �� �� U2G�$'1e1�t B ��    � (�MH�H�K�B�'� �tC�;�(۔1E��a����*0h.Z3�T0 k� ����U2G�$'1e1�t B ��    � (�SH�D �G�B�+� �tD�=�(۔0E��a����)0`/Z3�T0 k� ����U2G�$'1e1�t B ��    � (�YH�@!�C�B�3� �tD�>�,۔.E��`	���(0X/Z3�T0 k� ����U2G�$'1e1�t B ��    � (�_H�<#�?�B�;� �tD�@�,۔-F�_	���'0T0Z3�T0 k� ����U2G�$'1e1�t B ��    � (�eH�8$�;�B�?�LtD�B�,۔,F�^	���% L1Z3�T0 k� ��� U2G�$'1e1�t B ��    � (�kH�0'�7�B�O�LtE��E|,��)F�]	��x# @3Z3�T0 k� ��U2G�$'1e1�t B ��    � (�qH�,(�3�B�S�LtE��G|,��(F�]	��t! <4Z3�T0 k� �$�(U2G�$'1e1�t B ��    � (�wH�()�3�B�[�LtF��J|,��&F�\	.��p  45Z3�T0 k� �0�4U2G�$'1e1�t B ��    � (�|I(*�/�B�c�LtF��M|,��%F�\	.���l 06Z3�T0 k� �@�DU2G�$'1e1�t B ��    � (��I$,�+�B�g�LtF��O|,��$E��[	.���h (7Z3�T0 k� �L�PU2G�$'1e1�t B ��    � (��I -M+�B�o�LtG��R|,
��"E��[	.���h $8Z3�T0 k� �X�\U2G�$'1e1�t B ��    � (��I.M'�B�s�\tG��R|,	��!E��[	.���d  9Z3�T0 k� �h�lU2G�$'1e1�t B �    � (��I/M#�B�{�\tG4�T|,	�� E��[	���` :Z3�T0 k� �t�xU2G�$'1e1�t B ��    � (��I1M#�Bރ�\tG4�V|,��E��[	���` <Z3�T0 k� ��
��
U2G�$'1e1�t B ��    � (��I2M�Bއ�\tG4�Y|,��p+�[	���\=Z3�T0 k� ����U2G�$'1e1�t B ��    � (��I3M�Bޏ�\tG4�Y|,��p+�[	���\>Z3�T0 k� ����U2G�$'1e1�t B ��    � (��I4-�Bޗ�\tG4�Z|,��p+�[	���X?Z3�T0 k� ����U2G�$'1e1�t B ��    � (��I5-�Bޛ�\tG4�\|,��p+�[	.���X@Z3�T0 k� ����U2G�$'1e1�t B ��    � (��I6-�Bޣ� �tG4�^|,��p+�[	.���XAZ3�T0 k� ����U2G�$'1e1�t B ��    � (��I7-�Bާ� �tG4�_|,��p;�[	.���X�BZ3�T0 k� ����U2G�$'1e1�t B ��    � (��I 8-�Bޯ� �tG4�a|,��p;�[	.���X� CZ3�T0 k� �� �� U2G�$'1e1�t B ��    � (��I 9-�B޷� �tG4�c|,�� p;�[	.���X��DZ3�T0 k� ������U2G�$'1e1�t B ��    � '��I�:-�B޷� �tG4�d|,�� p;�[	���X��EZ3�T0 k� �����U2G�$'1e1�t B ��    � &��                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \���H ]�!�!� � ���4�  M `      ���    ������    
��$              
��           ���   
  ���  (	 
          ��o�   � � 
	   ����%    ��o����%           	            %	��          p�     ���   0	%
 
         ��>    
	   ��Z(    ���>��D�     C   	            ��           �P     ���   (	G  
          ��Ѵ   � �     
�    ��a 	P7    ���              ��           �Pb  �  ��� 0
		H         ��1�   � �
     .���.    ��7o���1    ��-              O ��             ��    ���   8'
         ���  ��	      B��R    �����R           
               ���]               �  ���    0 3             lW�        V��e�     lW���e�                       
 b 6         �      ��@   0
 	          [x�         j ���     [x� �oM      A                  j 5          K�     ��A   (
          ��c�    	     ~��    ��d��    ����               �� 6         ��     ��@   8�
         ��(O    	     ����q    �����
      ��a               	    �         	 ��     ��H  (
           ��  $ �     � ��     �� ���       ^                   	   �         
 �0     ��@   P

B         �����     � ���    ��� ��l       C                      ���                 ��@    8		 1                   ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��wt  ��        ���bc    ��j���m     ��a                   x                j  �    	   �                         ��    ��        ���      ��  ��           "                                                �                         ������ 
����� ����� � ������� 	 
               
 �   > �t H��T       3� �[� �$ `c` �� @d  �d d� �D �^@ �� _����J ����X � �d ]  ۄ ]  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0� ���� � �� �R� � }`���� � 
�\ W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����   ������  ������  
�fD
��L���"����D" � j  "  B   J jF�"  ""B�j"B ����
��"    B�j l �  B �
� �  �  
� ����  ��     ���      ��    ��     ���      ����  ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �)G      �� �T ��        �tT ���        �        ��        �        ��        �      ��    t�� q�        ��                         I:   +��                                    �                 ���� 	          	���� 	���%��  �� ��               25 Vincent Damphousse   4:37                                                                        1  1      �C
2� �HC. �@C4 �(C8 �DK �d K �0 � �/ � �	c� �0 
c� � �c~' c�/ �J� � �J� � �B� � � B� � �  � �	C � �C! � � C% �9"� �9 "� �)� �)
� �d"� �d "� �T"� �T*� �9"� �9 "� �)� �) 
� �  !"E � � "" | #"E �?$"* |_ "2 |?&"* |_ "2 | � ("  | )"J �?*"  |W !� |?,"* |_ "2 |  "G �O  "I �/ 0"& |?1"* |_ "2 |_ "2 |X  *KPP 5*ChX 6*GpX  *KP_ 8*Gg_  *KG:
�  ~ ;"Q � � <"O z � !� r � !� r. " �                                                                                                                                                                                                                         �� R        �     @ 
        B     P P E ]  ��        	            �������������������������������������� ���������	�
��������                                                                                          ��    ���   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, 5    :� i���@q���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ?    1    ��  $>�J      ,�  	                           ������������������������������������������������������                                                                     	                                                                    �    ��  �                    �      �          	     ������������������������ ���� � �  ���� ��������������� �������������������� ������������������������������ ������������� �������������������������������������������� ��  ����������� �������� ������ ����� ����� �� ���������������                           	                 �  L�J      ]                             ������������������������������������������������������                                                                                                                                             Q  4��              �          ��                 	 	 �� ��  ���� ������������ ������������� ��� �� ���� ����� ����� � �������������� ������� ��������� �� ������������  ������� ��������� �� ��  ������ ����������������������� ��� �����������������  � ����� ���������������������� �� �������� ����                                                                                                                                                                                                                                               
                                                   	                            �             


           �   }�                                                                             N�            ������������   /   ����������������������������  +	�����������������������������������������������������ww�ww333wwwwwwww�ww�ww�ww�ww333wwww > D 6                                 � RO� �\                                                                                                                                                                                                                                                                                         )n)h1p  �        m            l                  e      f      m                        ��                                                                                                                                                                                                                                                                                                                                                                              � � �  � ��  � ��  � 2��  � #��  EZm0  �N ������"�����.���������������������ؤ�����q                      �� [           �   & AG� �   �                 �                                                                                                                                                                                                                                                                                                                                      p I I   �      ��               !�� !��                                                                                                                                                                                                                        Y    �� �� Ѱ��      �� M      ������������������������ ���� � �  ���� ��������������� �������������������� ������������������������������ ������������� �������������������������������������������� ��  ����������� �������� ������ ����� ����� �� ��������������� �� ��  ���� ������������ ������������� ��� �� ���� ����� ����� � �������������� ������� ��������� �� ������������  ������� ��������� �� ��  ������ ����������������������� ��� �����������������  � ����� ���������������������� �� �������� ����               ���������������������������������������������������f��ff�fff�ff���������l�ff�ffffl��ff˼fllf������l��̼�ʗ���˹�ffjz�fkyl�l��fƨ�����������������������̼��̉������������������������������f���f�fff�ff�ffl�ff�flfl�l��xl�wwl���l̻�����˺��fl����l�xx��w��̻���l�f�f�ƻ�fl�����ffl�ffffffff���f���̚���ffflffflfffffffffflfffff������������������������l���l������f����������������������������l��lf��f�fff�f��l˪���ww��w�����flflffffffff�̼̙��fww��w��fx�̻�llffff�ffff���fl���f�l�l�˶����fffl��fflfll����ff��ff��lfl�lf��l���l�����������l�������l�������ʼ�j˚��̩��ʨ��ɘ���xxxȈ��ɉ�x���̇�̺������www��ww��xw���x��xk�����������wx��������������x����l�ƈ��Ƈ���w��Ɨ��̩z�̩yf̪�f�������������������������������̙i���ɖ�yɌ��ˌȉ̚ə̩���ə��Ɉ����x�̹x�̹�����������ƺ�������������������ˈ������˙������̫��̺�������˪�������������̸��̗�����̇��̇�����������������������̈���xx����x���w���ɉ��̨���k���̛̻�������������l��Ʀl�Ɗl�l���̻�lk��̺�f̩�l��f�ɫ�ˉ�lɊ�˙���ʚ���˙�˫̼���ɬ�̚��̼�����̼���̬������̼�����˻������������f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff���m�    A      +     ��                       M     �  ���������J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��       p���� ��     .T  �h  � >     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@      
g� ��   
g� �$ ^$  �� � ��� �� � ��� M� ���� �       �  ��   "���� e�����  g���         f ^�         �� ���      "      �������2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                                 � UP��f\�j�             �UUU] ���ff��������            U_� � �Uff�̪�������                �   �U�l�����fl                       �P  �     �   �j �̪ Pʪ \j��j����j��j����������̪�����P��P ��� ��������l�����UU�� �� ��U��̪����������jU��� \�] \�]U\�P���P������������j����ƪ�]�ʪ  ]�   l  ��� ��P ��[ ��[ l  ��  U   ����\j� Pƪ �ƪ �j     U��� ��] ���_��l����l����j�����������U�� U�� ���Uf��̪����������PU\�P \�P \�UU������f��������  \  ���ƪ��j��j���������������   mP  ��  ��P �l� �l� ��� �P            �                    P�j���f  U    �                ����������ffU���UU            �������ffl� �U]U_�             �f����UPU�                      P                    �          wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                               �   �   
                                       
   �  
   �  
   
   
    �   
�            ����        �   
    �   
    �  
   �  
   �      
   �  
   �  
   �  
   �                   ����   
   
   
   
   
   
   
   
   
   
�  

  
 � 
 
 
  �
  

   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        "! "   "      ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                   " ""   """! "   "      ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       "! "   "      ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        �  ��� ��� }�� wݪ �� 	�� �� �ͼ ��� ��� ̘� �ͻ +���"�8"8  8� �� �U��EU��3 ̻�"̰""�" ��" �"                             �   ��� �˹��˚���ڍ�̽���ͽ��ͽ���ݼ��л�� ��D �UT EUT UU0 C3  2"  ""  -�  ��  ��  �   � ��"/ �" � ���    �        �   ��  ��  ��  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                            � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                     �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                 �   ��  �   ��  ��  �  �  �   �                        �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                             � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                    0  300 11   10      �   �   �� �����  �    �   �   ,   "   "                   ���ۼ����� 9��C��UTDD�D33��0��  "��
/� � �, �"  �"   �   ˻ڛ��Ȱ��  ��  ��  TJ  EJ  DT  4E  �P  ��  �   /   ��  ��� �                                     � 	�� �� �˙	���
������                Ͱ  ˻  ˻  ۻ  ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                       �  ��                    �����                         �     �                                                                                                                                                                                   ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                      ��  ��  ��� ���                                                                                                                                                                                                   �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �           �   �     �   �                                         �     �                                      � ����ݼ� ����                                                                                                                                                                 �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��       �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �        � ��                    ���� �                                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   ��  ��  ��  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ��� ���                                                                                                                                                                                             	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                                  �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������            �   �   ��� ������ �   �      �       �                        �   ��  ���  � �    �                                ����                  �   �� �       �  �  ��  �   �   �   �                                    �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������                                ��  ��  ���  �  �  �   �   ��  �                            �   ���                            �   �                                                                                                                1    1   "    �   �   �� �����  �    �   �   ,   "   "                   ���ۼ����� 9��C��UTDD�D33��0��  "��
/� � �, �"  �"   �   ˻ڛ��Ȱ��  ��  ��  TJ  EJ  DT  4E  �P  ��  �   /   ��  ��� �                                     � 	�� �� �˙	���
������                Ͱ  ˻  ˻  ۻ  ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                       ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                                          �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""����������""""��������AD�I�""""��������AA�A�""""��������AI�I�""""����DD�I�""""��������DD""""�������IAA�I�""""�������������A��A��"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��������D�D�����3333DDDDM����D��D����3333DDDDA�A�A�D��M�D�����3333DDDDM�M�M�M��M�D����3333DDDD��A�M�M���M�����3333DDDDMDD�����D��D����3333DDDD��D��A�MD������3333DDDDA��A��A�AMMDDM����3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
2� �HC. �@C4 �(C8 �DK �d K �0 � �/ � �	c� �/ 
c� � �c~' c�/ �J� � �J� � �B� � � B� � �  � �	C � �C! � � C% �9"� �9 "� �)� �)
� �d"� �d "� �T"� �T*� �9"� �9 "� �)� �) 
� �  !"E � � "" | #"E �?$"* |_ "2 |?&"* |_ "2 | � ("  | )"J �?*"  |W !� |?,"* |_ "2 |  "G �O  "I �/ 0"& |?1"* |_ "2 |_ "2 |X  *KPP 5*ChX 6*GpX  *KP_ 8*Gg_  *KG:
�  ~ ;"Q � � <"O z � !� r � !� r. " �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������ �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������"��<�Z�K�V�N�G�T��6�K�H�K�G�[� � � � � � �7�=�6�����������������������������������������#��.�K�T�O�Y��<�G�\�G�X�J� � � � � � � � �7�=�6����������������������������������������� ��?�O�T�I�K�T�Z��.�G�S�V�N�U�[�Y�Y�K� � �7�=�6�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������7�=�6� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                