GST@�                                                           Zq     Z�                                               *            q            � h� ����J����������    ����        Ȁ      #    ����                                d8<n    �  ?    4�����  �
fD�
�L���"����D"� j   " B   J  jF�"    "�j* ,  �����
�"     �j@ �    ��
                                                                                  ����������������������������������      ��    ?o= 00 5o4 8 1  +     '       � 
   
           �	� 47� V� �	�                 Y 
         ::�����������������������������������������������������������������������������������������������������������������������������oo    og     +      '            ��                     	  7  V  	                  �            :8 �����������������������������������������������������������������������������                                D   N           @  &   q   �                                                                                 'w w  Y
  �    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E N �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ���E�.D�����	���c��C�z�_�E����3���|+�T0 k� �K��O�U8D"!%�0d    ��7 
   ��� ����E�.D�����	Ë�c��C�y�c�E����2���|+�T0 k� �O��S�U8D"!%�0d    ��7 
   ��� ����E�-D������	Ë�c��C�y�g�E����2��|+�T0 k� �S��W�U8D"!%�0d    ��7 
   ��� ��åE -D������	Ë�c��C�x�k�E����1��|+�T0 k� �W��[�U8D"!%�0d    ��7 
   ��� ��ϧE�,E������	Ë�c��C�v�k�E�#���1��|+�T0 k� �[��_�U8D"!%�0d    �7 
   ��� ��רE�,E������%���c��C�u�o�E�'���0��|+�T0 k� �[��_�U8D"!%�0d    ��7 
   ��� ��۩E� +E������%���c��C�t�o�E�/���0�#�|+�T0 k� �W��[�U8D"!%�0d    ��7 
   ��� ���E�,+E������%���c��C�t�s�E�3�� /�+�|+�T0 k� �W��[�U8D"!%�0d    ��7 
   ��� ���E�4+E������%���c��C�s�s�E�;��/�3�|+�T0 k� �W��[�U8D"!%�0d    ��7 
   ��� ���E�<+E������%���c��C�r�s�E�C��/�;�|+�T0 k� �O��S�U8D"!%�0d    ��7 
   ��� ���E�D+E������%���c��C�q�w�ErG��.�?�|+�T0 k� �O��S�U8D"!%�0d    ��7 
   ��� ����E�L*Eq�����%���c��C�p�w�ErO�� .�G�|+�T0 k� �K��O�U8D"!%�0d    ��7 
   ��� ����E�T*Eq��t�%���c��C�o�{�ErS��(.�O�|+�T0 k� �K��O�U8D"!%�0d    ��7 
   ��� ���E�\*Er�t�%���c��C�n�{�Er[��0-�W�|+�T0 k� �G��K�U8D"!%�0d    ��' 
   ��� ��D�h*Er�t�%���c��C�l�{�Er_��8-�_�|+�T0 k� �G��K�U8D"!%�0d    ��' 
   ��� ��D�p+Er�t�%���c��C k��Erg��@-�g�|+�T0 k� �K��O�U8D"!%�0d    ��' 
   ��� ��D�x+Er�t�%Û�c��Cj��Erk��H,�o�|+�T0 k� �K��O�U8D"!%�0d    ��'    ��� �#�Dр+Er���%ß�c��Ci��Ers��P,�w�|+�T0 k� �K��O�U8D"!%�0d    ��'    ��� �/�Dє+Er#���%ã�c��E�gӃ�Er��`+͇�|+�T0 k� �O��S�U8D"!%�0d    ��'    ��� �7�Dќ,Er'���%ã�c��E� fӃ�Er���d+͏�|+�T0 k� �O��S�U8D"!%�0d    ��'    ��� ��?�DѤ,Er+���%ã�c��E�$dӇ�Er���l+͗�|+�T0 k� �O��S�U8D"!%�0d    ��'    ��� ��G�DѰ,Er/���%ç�c��E�,cӇ�Eb���t+͟�|+�T0 k� �O��S�U8D"!%�0d    ��'    ��� ��O�DѸ-Eb3��#�%ç�c��E�4bӇ�Eb���|*ͧ�|+�T0 k� �S��W�U8D"!%�0d    ��'    ��� ��W�D��-Eb7��#�%ç�c��E�8aӋ�Eb����*ͯ�|+�T0 k� �S��W�U8D"!%�0d    ��'    ��� ��_�D��.Eb;�t'�%ç�c��E�@`Ӌ�Eb����*ͻ�|+�T0 k� �S��W�U8D"!%�0d    ��'    ��� ��g�D��.Eb?�t+�%���c��E�H^Ӌ�Eb����)�ÿ|+�T0 k� �S��W�U8D"!%�0d    ��'    ��� ��o�D��/EbC�t+�%���c��E�L]ӏ�Eb����)�˿|+�T0 k� �W��[�U8D"!%�0d    ��'    ��� ��w�D��/P�G�t/�%���c��E�T\ӏ�Eb��Τ)�ӿ|+�T0 k� �W��[�U8D"!%�0d    ��    ��� 	�D��0P�K�t3�%���c��E�X[ӏ�Eb��ά)�ۿ|+�T0 k� �W��[�U8D"!%�0d    ��    ��� 	��D��1P�O��3�%���c��E�`Yӓ�Eb��δ(��|+�T0 k� �[��_�U8D"!%�0d    ��    ��� 	��E� 1P�S��7�%���c��E�hXӓ�Eb��μ(��|+�T0 k� �[��_�U8D"!%�0d    ��    ��� 	��E�3P�[��7�%���c��E�tUӓ�ER����(���|+�T0 k� �[��_�U8D"!%�0d    ��    ��� 	��E�3P�_��;�%���c��E�xTӓ�ER����'��|+�T0 k� �_��c�U8D"!%�0d    �    ��� 	!��E�$4P�c��;�%���c��E��Sӗ�ER����'��|+�T0 k� �_��c�U8D"!%�0d    �    ��� 	!��E�05P�g��;�%ë�c��E��Qӗ�ER�� �' �|+�T0 k� �_��c�U8D"!%�0d    ��    ��� 	!��E�85P�k��;�%ë�c��E��Pӗ�ER�� �' #�|+�T0 k� �_��c�U8D"!%�0d    ��7    ��� 	!��E�@6P�o��;�%ë�c��E��Oӗ�E��� �& +�|+�T0 k� �c��g�U8D"!%�0d    ��7    ��� 	!��BBH6P�o��?�%ë�c��@��Mӗ�E��� �& 3�|+�T0 k� �c��g�U8D"!%�0d    ��7    ���  ��BBP7P�s��?�%ë�c��@��Lӗ�E���  & ;�|+�T0 k� �c��g�U8D"!%�0d    ��7    ���  ��BBX8P�w��?�%ë�c��@��Kӗ�E��� & C�|+�T0 k� �c��g�U8D"!%�0d    ��7    ���  ��BB`8P�{��;�%ë�c��@��Jӗ�E��� % K�|+�T0 k� �c��g�U8D"!%�0d    ��7    ���  ��BBh9P���;�%ë�c��@��Iӗ�E��� % S�|+�T0 k� �c��g�U8D"!%�0d    ��7    ���  ��BBp:P���;�%ë�c��@��Hӛ�E��� % [�|+�T0 k� �g��k�U8D"!%�0d    ��7    ���  ��BBx:P����;�%ë�c��@��Fӛ�A��� $% c�|+�T0 k� �g��k�U8D"!%�0d    ��7    ���  ��BB�;A����;����c��@��Eӛ�A��� (% g�|+�T0 k� �g��k�U8D"!%�0d    ��G    ���  ��BB�;A����;����c��@��D��A��� 0$ o�|+�T0 k� �k��o�U8D"!%�0d    ��G    ���  ��BB�<A����;����c��@��C��A��� 4$ w�|+�T0 k� �o��s�U8D"!%�0d    ��G    ���  ��BB�<A����;����c��@��B��A��� <$ �|+�T0 k� �s��w�U8D"!%�0d    �G    ���  ��BB�=A����;����c��@��A��A��� @$ ��|+�T0 k� �w��{�U8D"!%�0d    ��O    ���  ��BB�=A����;�3��c��@��@��A��� H$ ��|+�T0 k� �{���U8D"!%�0d   ��O    ���  �BB�>A����;�3��c��@��?��A��  L$ ��|+�T0 k� �����U8D"!%�0d   ��O    ���  �BB�>A����;�3��c��@��>��A�� T# ��!�+�T0 k� Ã����U8D"!%�0d   ��O    ���  �BB�?A����;�3��c��@��=��A�� X# ��!�+�T0 k� Ç����U8D"!%�0d   ��O    ���  �BB�?A�� �;�3��c��@��<S��A�� `# ��!�+�T0 k� Ë����U8D"!%�0d   ��O    ���  �BB�@A�� �;�3��c��@��;S��A�� d# ��!�+�T0 k� ӏ����U8D"!%�0d   �O    ���  �BB�@A���;����c��@��:S��A�� l# ��!�+�T0 k� ӓ����U8D"!%�0d   ��O    ���  �BB�AA���7����c��@��9S��A�� p" ��!�+�T0 k� ӗ����U8D"!%�0d   ��O    ���  #�BB�AA���7����c��@��8S��A�� t" ��!�+�T0 k� ӛ����U8D"!%�0d   ��O    ���  '�BB�BA���7����c��@��7��A�� |" ǿ!�+�T0 k� ӟ����U8D"!%�0d  	 ��O    ���  +�BB�BA���7����c��@� 6��A�� �" ˿!�+�T0 k� �����U8D"!%�0d  	 ��/    ���  /�BB�CEb��7����c��@�5��A�� �" Ͽ!�+�T0 k� �����U8D"!%�0d  
 ��/    ���  3�BB�CEb�T7�ë�c��@�5��A�� �" ׿!�+�T0 k� �����U8D"!%�0d   ��/    ���  7�BB�DEb�T7�ë�c��@�4��A��	 �" ۿ|+�T0 k� �����U8D"!%�0d   $�/    ���  ;�BB�DEb�T7�ë�c��@�3#��A��	 �! �|+�T0 k� �����U8D"!%�0d   ��U    ���  ?�BC DEb�T7�ë����@�2#��A��
 �! �|+�T0 k� �����U8D"!%�0d   ��U   ���  C�BCEEb�T7�ë����@�1#��A�� �! �|+�T0 k� �����U8D"!%�0d   ��U    ���  G�BCEEb�T7�ë����@�1#��A�� �! �|+�T0 k� �����U8D"!%�0d   �U    ���  K�BCFEb�	T7�ë����@�0#��A�� �! ��|+�T0 k� �����U8D"!%�0d   ��O    ���  O�BCFEb�
T7�ë����@� /#��A�� �! ��|+�T0 k� �����U8D"!%�0d   ��O    ���  O�BCFEb�
T7�ë����@�$.3��A�� �! ��|+�T0 k� �����U8D"!%�0d   ��O    ���  S�BC GA��T7�������@�(-3��A�� �  �|+�T0 k� ����U8D"!%�0d   ��O    ���  W�BC(GA��T7�������@�(.3��A�  �  �|+�T0 k� s��w�U8D"!%�0d   ��O 