GST@�                                                           �j�                                                       ���   @                   ����e ��	 ʴ����������P���z���        �h     #    z���                                d8<n    �  ?     �J����  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    $�j� � �$  ��
  ��                                                                              ����������������������������������      ��    bb QQb  114 44c c   c      		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������=o  0  4g  1                      �                         �  �  �  �                  �  
          8 �����������������������������������������������������������������������������                                D   $           @  &   r   �                                                                                 'w w  )n)n1n  
�    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E $ �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    B�xQ�xB���N$R�|$ ��BϐE��41��b3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B��RҀB���N$R�|$ ��BϔE��41��c3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B��R҄B���N$R�|$ �BϘE��31��c3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B��SB�ð�$R� |$ '�BϜE� 21�� d3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B��TB�ǰ�(R�$|$ /�BϠE�11��(e3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B��TB�ϰ�(R�(|$ 7�BϤE�11��0e3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B��U B�װ�(R�(|$ ?�BϬE�01�8f3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B��V¤B�߰�,R�,|$ G�BϰC�/1�@g3�T0 k� �� �� %�@c  I%1t'2Q  ��    �   �BдW¬B���,R�0|$ O�BϴC�.1�Hg3�T0 k� �� �� %�@c  I%1t'2Q  ��    �   �BмW´B���,R�4|$ W�BϸC� -1�Ph3�T0 k� �� �� %�@c  I%1t'2Q  ��    �   �B��X¸B����0R�8|$ c�B��C�$,1�Xh3�T0 k� �� �� %�@c  I%1t'2Q  ��    �   �B��Y��B����4R�<|$ �k�B��C�(+1�`i3�T0 k� ������%�@c  I%1t'2Q  ��    �   �B��Z��B���8R�D|$ �{�B��C�4)1#�pj3�T0 k� ������%�@c  I%1t'2Q  ��    �   �B��Z��B���<R�H|$ ���B��E38(1#��xk3�T0 k� ������%�@c  I%1t'2Q  ��    �   �B��[��B���<R�P|$ ���B��E3<'1#���k3�T0 k� ������%�@c  I%1t'2Q  ��    �   �B��\��B�'��@R�T|$ ���B��E3@$1#���l3�T0 k� ������%�@c  I%1t'2Q  ��    �   �B��\��B�/��DR�X|$ ���B��E3D!1'���l3�T0 k� ������%�@c  I%1t'2Q  ��    �   �B� ]��B�;��HR�\|$ ���B��E3H1'���l3�T0 k� ������%�@c  I%1t'2Q  ��    �   �B�]��B�C��LR�d|$ ���B��C3L1'���m3�T0 k� �����%�@c  I%1t'2Q  ��    �   �B�^��B�K��PR�h|$ ���B� C3P1'���m3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B�^��B�S��TR�p|$ ���B�C3P1'���m3�T0 k� ����%�@c  I%1t'2Q  �    �   �B�_��B�[��XR�t|$ �ǼB�C3T1+���m3�T0 k� �+��/�%�@c  I%1t'2Q ��    �   �B�$`� B�g��\R�x|$ �ϼB�C3X1+���m3�T0 k� �?��C�%�@c  I%1t'2Q ��    �   �B�,`�B�o��`Rހ|$ �ۼB� C3\1+���m3�T0 k� �S��W�%�@c  I%1t'2Q ��    �   �B�4a�Ew��hRވ |$ ��B�(C3`1+���n3�T0 k� �g��k�%�@c  I%1t'2Q ��    �   �B�<a�E��lRތ |$ ��B�0C3d1+���n3�T0 k� �{���%�@c  I%1t'2Q ��    �   �B�Db�E���pRޔ |$ ��E�8C3h	1+���n3�T0 k� ������%�@c  I%1t'2Q ��    �   �B�Lb	E���tRޘ |$ ���E�@C3l1/���nC�T0 k� ������%�@c  I%1t'2Q $�    �   �B�Pc	E���|Rޠ |$ ��E�HC3l1/���mC�T0 k� ������%�@c  I%1t'2Q ��    �   �B�Xc	 E���΀Rި |$ ��E�PC3p1/�� mC�T0 k� ������%�@c  I%1t'2Q ��    �   �B�`d	$E���ΈRޯ�|$ ��E�XC3t 1/��mC�T0 k� ������%�@c  I%1t'2Q ��    �   �B�hd	,E���ΌR���|$ ��E�`C3{�1/��mC�T0 k� ������%�@c  I%1t'2Q ��    �   �B�pe	0E���ΔR���|$ �'�E�hC3{�1/��mC�T0 k� ������%�@c  I%1t'2Q ��    �   �B�xe	4E�ǰΘR���|$ �/�D�pC3{�1/�� mC�T0 k� ������%�@c  I%1t'2Q ��    �   �B��e	8e�ϰΠR���|$ �7�D�xC3�13��(lC� T0 k� ������%�@c  I%1t'2Q ��    �   �B��f	<e�װޤR���|$ �?�DЀC3��13��0lC� T0 k� ������%�@c  I%1t'2Q ��    �   �B��f	@e��ެR���|$ �G�DЈC3��13��<lC� T0 k� ������%�@c  I%1t'2Q ��    �   B��g	De��޴R���|$ �O�DАC3��13�sDkC� T0 k� ������%�@c  I%1t'2Q ��    �   B��g	He��޸R���|$ �W�DИC3��13�sLkC� T0 k� ������%�@c  I%1t'2Q ��    �   B��h	Pe����R���|$ �g�DШC3��13�s\jC� T0 k� ������%�@c  I%1t'2Q ��    �   B��h	Te����R��|$ �o�DаEÓ�17�sdjC� T0 k� ������%�@c  I%1t'2Q ��    �   B��i	Xe����R��|$ �w�E��EÓ�17�sliC� T0 k� ������%�@c  I%1t'2Q ��    �   B��i	Xe����Q��|$ ��E��E×�17�sphC� T0 k� ������%�@c  I%1t'2Q ��    �   B��j	\e�#���Q��|$ ���E��E×�17�sxhC� T0 k� ������%�@c  I%1t'2Q ��    �   B��j	`e�+���Q��|$ ���E�� E×�17�s�gC��T0 k� ������%�@c  I%1t'2Q ��    �   B��j	de�/���Q�'�|$ ���E��!EÛ�17�s�fC��T0 k� ������%�@c  I%1t'2Q ��    �   B��k�he�7���P�/�|$ �E��"EÛ�A7���eC��T0 k� ������%�@c  I%1t'2Q ��    �   B��k�le�?�� P7�|$ �E��#EÛ�A7���dC��T0 k� ������%�@c  I%1t'2Q ��    �   B��l�te�O��OG�|$ ¯�E��$Eß�A;���bC��T0 k� ������%�@c  I%1t'2Q  -�    �   �B�l�xe�S��OO�|$ ³�E� %C���A;���aC��T0 k� ������%�@c  I%1t'2Q  ��    �   �B�m�|e�[��NW�|$ ·�Eq&C���A;���`C��T0 k� ������%�@c  I%1t'2Q  ��    �   �B�mӀe�c��$M_�|$ ¿�Eq'C���A;�s�_C��T0 k� ������%�@c  I%1t'2Q  ��    �   �B�m��e�g��,Mc�|$ ���Eq(C���A;�s�^C��T0 k� ������%�@c  I%1t'2Q  ��    �   �B�$n��e�o��4Lk�|$ ���Eq )C���A;�s�]C��T0 k� ������%�@c  I%1t'2Q ��    �   �B�4n��e�{��@K{�|$ ���Eq,+Eß�;�s�ZC��T0 k� ������%�@c  I%1t'2Q ��    �   �B�8o��
e��HJ��|$ ���Eq4-Eß�?�s�YC��T0 k� ������%�@c  I%1t'2Q ��    �   �B�@o��
e��PJ���|$ ���Eq<.Eß�?�s�WC��T0 k� ������%�@c  I%1t'2Q ��    �   �B�HoÔ	e��XI���|$ ���Eq@/Eß�?�s�VC��T0 k� ������%�@c  I%1t'2Q ��    �   �B�PpÔ	e��`I���|$ ���EqH0Eß�?�s�Ts��T0 k� ������%�@c  I%1t'2Q �    �   �B�`pÜ	e��pG��|$ ���EqT3EÛ�?�s�Qs��T0 k� ������%�@c  I%1t'2Q ��    �   �B�hpàe��tG��|$ ���Eq\5Eӛ�?�s�Ps��T0 k� ������%�@c  I%1t'2Q ��    �   �B�pqӤe��|F��|$ ���Eqd6Eӗ��?�d Ns��T0 k� ������%�@c  I%1t'2Q ��    �   �B��qӬE����D��|$ ���Eap9Eӗ��C�dKs��T0 k� ������%�@c  I%1t'2Q ��    �   �B��rӰE����D��|$ ���Eat;Eӓ��C�dIs��T0 k� ������%�@c  I%1t'2Q  ��    �   �B��rӴE�ø�C��|$ ���Ea|<Eӏ��C�dHs��T0 k� ������%�@c  I%1t'2Q  ��    �   �B��rӸE�˸�B��|$ ���Ea�>Eӏ��G�dFs��T0 k� ������%�@c  I%1t'2Q  ��    �   �B��r�E�Ϲ�A���|$ ���Ea�@EӋ��G�dDs��T0 k� ������%�@c  I%1t'2Q  ��    �   �B��s��E�ۺ�@���|$ ���Ea�CEӇ��K�d$As��T0 k� ������%�@c  I%1t'2Q  /�    �   �B��s��E����?���|$ ���Ea�ECレ�O�4(?���T0 k� ������%�@c  I%1t'2Q  ��    �   �E��t��E����>���|$ ���Ea�FC���S�4,>���T0 k� ������%�@c  I%1t'2Q  ��    �   �E��t��E����=	���|$ ���Ea�HC�{��S�40<���T0 k� ������%�@c  I%1t'2Q  ��    �   �E��t��Er����=	��|$ ���Ea�JC�{��W�40:���T0 k� ������%�@c  I%1t'2Q  ��    �   �E��u��Es���;	��|$ 2��Ea�ME�s��[�d87���T0 k� ������%�@c  I%1t'2Q  ��    �   �E��u��Es���:	��|$ 2��Ea�OE�o��_�d85���T0 k� ������%�@c  I%1t'2Q  ��   �   �E��u��Es���9
 �!�$ 2��Ea�QE�k��c�d<3���T0 k� ������%�@c  I%1t'2Q  ��    �   �E��v�� Es�� 8
 #�!�$ 2��EQ�TE�c��k�d@/���T0 k� ������%�@c  I%1t'2Q  ��   �   �E�v�� Es#��7
 '�!�$ 2��EQ�VE�_��o�d@-���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�v���Es'��6
 +�!�$ 2��EQ�XE�[��s�d@+���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�v���Es/�p5p/�!�$ B��EQ�YE�W��w�dD*���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�$w���Es;�p 3p7�!�$ B��EQ�]E�K���d@*���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�,w���Es?�p(2p?�!�$ B��EQ�^E�G����d@+���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�4w���EsC�p01pC�!�$ B��EQ�`E�C����T<+���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�Dw���EcO�p</pK�!�$ B��EQ�cE�7����T8,���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�Lw��EcS�pD.pO�|$ B��EQ�eE�3����T8,���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�Tw��EcW�pH,pS�|$ B��EQ�fE�+���T4-���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�\w��Ec_�pP+pW�|$ B��EA�hE�'���T0-���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�lw��Ecg�p\)p_�|$ B��EA�jD3���T,.���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�tw��Eck�p`(pc�|$ R��EA�lD3���T(.���T0 k� ������%�@c  I%1t'2Q  ��    �   �E�|w��Eco�ph&`g�|$ R��EA�mD3����$/���T0 k� �����%�@c  I%1t'2Q  ��    �   �E��w��Eco�`l%`k�|$ R��EA�nD3���� /���T0 k� �{���%�@c  I%1t'2Q  ��    �   �E��v��Ecw�`x"`s�|$ R��EA�pD2�����0c��T0 k� �w��{�%�@c  I%1t'2Q  ��    �   �E��v��Ecw�`|!`s�|$ R��EA�qD2������0c��T0 k� �s��w�%�@c  I%1t'2Q  �    �   �E��v��Ts�`� `w�!�$ R��EA�rD2�����0c��T0 k� �o��s�%�@c  I%1t'2Q  ��    �   �E��u��Tk�`�`{�!�$ R��EA�tD2�����1c��T0 k� �_��c�%�@c  I%1t'2Q �    �   �E��t��Tg�`�`�!�$ R��EA�uD2߂���� 1S��T0 k� �S��W�%�@c  I%1t'2Q ��    �   �E��t��Tg�`�`�!�$ R��E��uD2ׁ�����2S��T0 k� �K��O�%�@c  I%1t'2Q ��    �   �E��s��Tc�`�`��!�$ b��E��vDBӀ�����2S��T0 k� �C��G�%�@c  I%1t'2Q ��    �   �E��s��T_�`�`��!�$ b��E��wDBˁ����2S��T0 k� �;��?�%�@c  I%1t'2Q ��    �   �E��q��TW�`�`��!�$ b��E��xDB������3S��T0 k� �+��/�%�@c  I%1t'2Q ��    �   �E��p��T#W��P��!�$ b��EєxDB������3S��T0 k� �#��'�%�@c  I%1t'2Q ��    �   �E��p��T#S��P��!�$ b��EѐyDB���#���4c��T0 k� ����%�@c  I%1t'2Q ��    �   �E��o��T#O��P��|$ R��EѐzE⫂�+���4c��T0 k� ����%�@c  I%1t'2Q ��    �   �E��m��T#K��P��|$ R{�Eф{E⛃�;���4c��T0 k� ��� %�@c  I%1t'2Q ��    �   �E��l��T#G��
���|$ Rs�Eр{EⓄ�C���4c��T0 k� ����%�@c  I%1t'2Q ��    �   �E� k��T#C��	���|$ Ro�E�||E⏄�C��5c��T0 k� ����%�@c  I%1t'2Q ��    �   �E�j��T3C�����|$ Rk�E�x|E⇅�G��5c�T0 k� ����%�@c  I%1t'2Q ��    �   �E�i��T3?�����|$ Rg�E�t}E���K��5c�T0 k� ����%�@c  I%1t'2Q ��    �   }E�g��T3;�	�����|$ R[�E�h~E�o��S��4c{�T0 k� ����%�@c  I%1t'2Q ��    �   yE�f��T37�	�� ���|$ RW�E�d~E�k��W��4Sw�T0 k� ����%�@c  I%1t'2Q	 ��    �   uE�e��T33�	������|$ �S�E�\}E�c��[��4Sw�T0 k� ����%�@c  I%1t'2Q	 ��    �   rE� d��T33�	������|$ �O�E�X}E�[��_�	��4Ss�T0 k� ����%�@c  I%1t'2Q	 ��    �   oE� c��T3/�	�����|$ �K�E�P}E�S��c�	��4Ss�T0 k� ����%�@c  I%1t'2Q	 ��    �   lE�$b��T3/�	����{�|$ �C�D1L}E�K��k�	�|4So�T0 k� ����%�@c  I%1t'2Q	 ��    �   iE�(a��T3+�	����{�|$ �?�D1H|E�G��o�	�t4So�T0 k� �� �� %�@c  I%1t'2Q	 ��    �   fE�,`��T3'�	����w�|$ �;�D1@|E�?��s�	�l4Sk�T0 k� ��#��#%�@c  I%1t'2Q	 ��    �   cE�0^��T3#�	����s�|$ �/�D14|E�3��{�	�d4Sg�T0 k� �|'��'%�@c  I%1t'2Q	 ��    �   `E�0]��T3#�	����o�|$ �'�EQ,{E�+����	�\4Sg�T0 k� �t*�x*%�@c  I%1t'2Q	 ��    �  ]E�4\��T3�	���Pk�|$ �#�EQ({E�#����	�X4Sc�T0 k� �h,�l,%�@c  I%1t'2Q	 ��    �  ZE�4[��T3�	���Pg�|$ ��EQ {D�����	�T4Sc�T0 k� �`.�d.%�@c  I%1t'2Q	 ��    �  WE�4Z��T3�	���Pc�|$ ��EQ{D�����	�L4S_�T0 k� �X1�\1%�@c  I%1t'2Q	 ��    �  TC�8Y��T3�	���P_�|$ ��EQ{D�����	�H4S_�T0 k� �P3�T3%�@c  I%1t'2Q	 ��    �  QC�8X��T3�	���P[�|$ ��E�zD������D4S_�T0 k� �H6�L6%�@c  I%1t'2Q	 ��    �  NC�8W��T3�	���PW�|$ ���E�zD������@4S[�T0 k� �@8�D8%�@c  I%1t'2Q	 ��    �  KC�8V��T3�	���PS�|$ ���E��zD�������<3S[�T0 k� �8:�<:%�@c  I%1t'2Q ��    �  HC�8U��T3�	���PO�|$ ���E��zD�������83SW�T0 k� �,=�0=%�@c  I%1t'2Q ��    � 	 EC�8T��T3�	���@K�|$ ���E��yD������43sW�T0 k� �$?�(?%�@c  I%1t'2Q ��    � 
 BC�8S��T3�	���@G�|$ ���E��yD������03sS�T0 k� �B� B%�@c  I%1t'2Q ��    �  ?C�8S��T3�	���@C�|$ ���E��yD������,2sS�T0 k� �D�D%�@c  I%1t'2Q ��    �  <C�4R��T3�	���@;�|$ ���E��yD������(2sO�T0 k� �F�F%�@c  I%1t'2Q ��    �  9C�4P��T3�	����3�|$ ���E��xD�ס���� 1�K�T0 k� ��K� K%�@c  I%1t'2Q ��    �  6C�0O��T3�	����/�|$ ��D0�xD�ӣ����0�G�T0 k� ��N��N%�@c  I%1t'2Q ��    �  3C�0N��T2��	����'�|$ ��D0�xD�Ϥ���0�C�T0 k� ��P��P%�@c  I%1t'2Q ��    �  0C�0N��T2��	����#�|$ ��D0�wD�Ǧ���/�?�T0 k� ��R��R%�@c  I%1t'2Q ��    �  -C�,M��T2��	�����|$ ��D0�wD�ç���.�?�T0 k� ��U��U%�@c  I%1t'2Q ��    �  +C�,L��T2��	�����|$ ��D0�wD������-�?�T0 k� ��W��W%�@c  I%1t'2Q ��    �  )C�(K��T2��	�����|$ ��EP�wD�����-�;�T0 k� ��Y��Y%�@c  I%1t'2Q ��    �  'C�$K��T2��`����|$ ��EP�vD�����,�7�T0 k� ��\��\%�@c  I%1t'2Q ��    �  %C�$J��T2��`����|$ ��EP�vD�����+�7�T0 k� ��^��^%�@c  I%1t'2Q ��    �  "C� I��T2��`����|$ �EP�vD����� *�7�T0 k� ��a��a%�@c  I%1t'2Q ��    �   C�H��T2��`�����|$ w�EPxvD������ )�3�T0 k� ��c��c%�@c  I%1t'2Q ��    �  C�H��T2��`�����|$ o�EPpvD����'�� (�/�T0 k� ��e��e%�@c  I%1t'2Q  �    �  C�G��T2��P����|$ Qg�EPluD����/���(�+�T0 k� ��h��h%�@c  I%1t'2Q  ,�    �  DF��T2��P���|$ Q[�APduD����3���'�'�T0 k� ��j��j%�@c  I%1t'2Q  ��    �  DF��T2��P���|$ QS�AP\uD����;���&�#�T0 k� ��m��m%�@c  I%1t'2Q  ��    �  DE��T2��P��߅|$ QK�APXuD����C���&��T0 k� �xo�|o%�@c  I%1t'2Q  ��    �  DD��T2��P��ۅ|$ QC�APPuD����G���%��T0 k� �pq�tq%�@c  I%1t'2Q ��    �  D D��T2��P��ӆ|$ Q7�APHtD����O���$��T0 k� �ht�lt%�@c  I%1t'2Q ��    �  D�C��T2��P��φ|$ /�I�DtD����S���$��T0 k� �`v�dv%�@c  I%1t'2Q ��    �  D�C��T2��P��ˇ|$ '�I�<tD����[���#��T0 k� �Xx�\x%�@c  I%1t'2Q ��    �  D�B��T2��P��Ǉ|$ �I�8tD����_���#��T0 k� �P{�T{%�@c  I%1t'2Q ��    �  AS�A��T2��P����|$ �I�0tD����g���#��T0 k� �H}�L}%�@c  I%1t'2Q ��    �  AS�A��T2��P����|$ �I�,tD����k���#���T0 k� �@��D�%�@c  I%1t'2Q ��    �  AS�@��T2��P����|$ �E�$tD���o���"���T0 k� �4��8�%�@c  I%1t'2Q ��    �  AS�@��T2��P����|$ ��E�tD���s���"���T0 k� �,��0�%�@c  I%1t'2Q )�    �  AS�?��T2��P����|$ ��E�tD�{��{��"���T0 k� 1$��(�%�@c  I%1t'2Q ��    �  E��?��T2��P����|$ �E�tD�w����"���T0 k� 1�� �%�@c  I%1t'2Q ��    �  E��>��T2��P����|$ �E�sD�w�Ã��"���T0 k� 1���%�@c  I%1t'2Q ��    �  E��>��T2��P����|$ �E�sD�s�Ç��"���T0 k� 1���%�@c  I%1t'2Q ��    �  E��=��T2��P����|$ ۳E��sD�o�Ë��"���T0 k� 1���%�@c  I%1t'2Q ��    �  E��=��T2��P����|$ ӲE��sD�o�Ë���"���T0 k� ���� �%�@c  I%1t'2Q ��    �  E��<��T2��P����|$ ϲE��rD�k�Ï���#���T0 k� �����%�@c  I%1t'2Q ��    �  EӼ<�T2��P����|$  ǱE��rD�g�Ó���#���T0 k� �����%�@c  I%1t'2Q ��    �  EӸ;�T2��P����|$  ��E��rD�g�×���#⿿T0 k� ����%�@c  I%1t'2Q  ��    �  AS�;�T2��P����|$  ��E��rD�c�Ӕ ��#ⷽT0 k� ��~��~%�@c  I%1t'2Q  ��    �  AS�:�T2��P����|$  ��E��qD�c�Ә��#⳼T0 k� ��~��~%�@c  I%1t'2Q  ��    �  AS�:�T2��P���|$  ��E��qD�_�Ә��#⫺T0 k� ��}��}%�@c  I%1t'2Q  ��    �  AS�9�T2��P��{�|$  ��E��qD�[�Ӝ��#⧹T0 k� ��}��}%�@c  I%1t'2Q  /�    �  AS�9�T2��P��w�|$  ��E��qD�[�Ӝ��#⟷T0 k� �|��|%�@c  I%1t'2Q  ��    �  AS�8�T2��P��s�|$  ��E��pEaW����#⛶T0 k� �{��{%�@c  I%1t'2Q  ��    �  AS�8�T2��P��o�|$  ��E��pEaS����#⓵T0 k� @�{��{%�@c  I%1t'2Q  ��    �  AS�7��T2��P��k�|$  ��F�pEaS����#⏳T0 k� @�z��z%�@c  I%1t'2Q  ��    �  AS�7��T2��P��g�|$  ��F�pEaO����#⇲T0 k� @�z��z%�@c  I%1t'2Q  ��    �  AS�7��T2��P��c�|$  ��F�pEaK����#⃰T0 k� @�y��y%�@c  I%1t'2Q  ��    �  AS�6��T2��P��_�|$  �F�oL1K��	�#��T0 k� @�y��y%�@c  I%1t'2Q  ��    �  AS�6��T2��P��[�|$  w�F�oL1G��
�#�w�T0 k� ��x��x%�@c  I%1t'2Q  ��    �  AS�5��T2��P��[�|$  s�F�oL1G���#�s�T0 k� �xw�|w%�@c  I%1t'2Q  ��    �  AS�5��T2��P��W�|$  o�F�pL1C���#�k�T0 k� �pw�tw%�@c  I%1t'2Q  ��    �  AS�5��T2��P��S�|$  g�F�pL1?���$�g�T0 k� �hv�lv%�@c  I%1t'2Q  ��    �  AS|4��T2��P��O�|$  c�F�pL1?���$�_�T0 k� �`v�dv%�@c  I%1t'2Q  ��    �  ASx4D�T2��P��K�|$  _�E��pL1;���$�[�T0 k� �Xu�\u%�@c  I%1t'2Q  ��    �  ASt4D�T2��P��K�|$  [�E��pL1;���$�S�T0 k� �Pu�Tu%�@c  I%1t'2Q  ��    �  ASp3D�T2��P��G�|$  S�E��pL17���$�O�T0 k� �Ht�Lt%�@c  I%1t'2Q  ��    �  ASl3D�T2��P��C�|$  O�E��pL17���$�G�T0 k� �@s�Ds%�@c  I%1t'2Q  ��    �  ASl2D�T2��P��?�|$  K�E��qLA3���$�C�T0 k� �8s�<s%�@c  I%1t'2Q  ��    �  ASh2D�T2��P��?�|$  G�E��qLA0��$�;�T0 k� �0r�4r%�@c  I%1t'2Q  ��    �  ASd2D�T2��P��;�|$  C�E�|qLA,�|$�7�T0 k� �(r�,r%�@c  I%1t'2Q  ��    �  AS`1D�T2��P��7�|$  ;�E�|qLA,�x$�/�T0 k� � q�$q%�@c  I%1t'2Q  ��    �  AS`1D�T2��P��3�|$  7�E�|qLA(�t$�+�T0 k� �q�q%�@c  I%1t'2Q  ��    �  AS\1D�T2��P��3�|$  3�E�|qLA(�p$�'�T0 k� �p�p%�@c  I%1t'2Q  ��    �  ASX0D�T2��P��/�|$  /�E�xqLA$�l$��T0 k� �o�o%�@c  I%1t'2Q  ��    �  ASX0D�T2��P��+�|$  +�E�xqLA$
�h$��T0 k� � o�o%�@c  I%1t'2Q  ��    �  AST0D�T2��P��+�|$  '�E�xqLA #�d$��T0 k� ��n��n%�@c  I%1t'2Q  ��    �  ASP0D�T2��P��'�|$  #�@oxqLA #�`$��T0 k� ��n��n%�@c  I%1t'2Q  ��    �  ASL/D�T2��P��'�|$  �@oxqLA#�"X$��T0 k� ��m��m%�@c  I%1t'2Q  ��    �  ASL/D�T2��P��#�|$  �@otqLA#�"T$��T0 k� ��m��m%�@c  I%1t'2Q  ��    �  ASH/D�T2��P���|$  �@otqLA#�"P$���T0 k� ��l��l%�@c  I%1t'2Q  ��   �  ASH.D�T2�P���|$  �@otqLA#�"L$���T0 k� ��l��l%�@c  I%1t'2Q  ��    �  ASD.D�T2�P���|$  �@otqLA#�"H$��T0 k� ��k��k%�@c  I%1t'2Q  ��    �  AS@.D�T2�P���|$  �@otqLA#�"D$��T0 k� ��j��j%�@c  I%1t'2Q  ��    �  AS@.D�T2{�P���|$  �@oprLA#�"@$��T0 k� ��j��j%�@c  I%1t'2Q  ��    �  AS<-D�T2{�P���|$  �@oprLA#�"@%�ۈT0 k� ��g��g%�@c  I%1t'2Q  ��    �  AS<-D�T2{�P���|$ /��@oprLA#�"<%�ׇT0 k� ��e��e%�@c  I%1t'2Q  ��    �  AS8-D�T2{�P���|$ ��@oprLA#�"8%�υT0 k� ��d��d%�@c  I%1t'2Q  ��    �  AS4-D�TBw�P���|$ ��@oprLA#�"4%�˄T0 k� ��d��d%�@c  I%1t'2Q  ��    �  AS4,D�TBw�P���|$ ��@oprLA#�"0%�˄T0 k� ��c��c%�@c  I%1t'2Q  ��    �  AS0,D�TBw�P���|$ �@olrLA#�",%�˃T0 k� ��b��b%�@c  I%1t'2Q  ��    �  AS0,D�TBw�P���|$ �@olrLA#�"(%1˃T0 k� ��b��b%�@c  I%1t'2Q  ��    �  AS,,D�TBs�P���|$ �@olrLA#� "$%1˂T0 k� ��b��b%�@c  I%1t'2Q  ��    �  AS,+D�TBs�P���|$ _�@olrLA #� " %1˂T0 k� ��b��b%�@c  I%1t'2Q  ��    �  AS(+D�TBs�P���|$ _�@olrLA!#�!" %1ˁT0 k� ��b��b%�@c  I%1t'2Q  ��    �  AS(+D�TBs�P����|$ _�@olrLA"#�!"%1ˁT0 k� ��b��b%�@c  I%1t'2Q  ��    �  AS$+D�TBo�P����|$ _ߣK�lrLA##�""%1ˀT0 k� ��f��f%�@c  I%1t'2Q  ��    �  AS$*D�URo�P���|$ _ۣK�hrLA $#�""%�ˀT0 k� �xi�|i%�@c  I%1t'2Q  ��    �  AS *D�URo�P���|$ OףK�hrLA %#�#"%��T0 k� �tk�xk%�@c  I%1t'2Q  ��    �  AS *D�URo�P���|$ OӣK�hrLA &#�#"%��T0 k� �pl�tl%�@c  I%1t'2Q  ��    �  AS*D�URo�P���|$ OˣK�hrL@�'#�#"%��~T0 k� �hm�lm%�@c  I%1t'2Q  ��    �  AS*D�URk�P��|$ OǣK�hrL@�(#�$"%��~T0 k� �hn�ln%�@c  I%1t'2Q  ��   �  AS)D�URk�P��|$ OãK�hrL@�)#�$"%��}T0 k� �ho�lo%�@c  I%1t'2Q  ��    �  AS)D�URk�P��|$ ?��K�hrL@�*#�%"%��}T0 k� �ho�lo%�@c  I%1t'2Q  ��    �  AS)D�URk�P��|$ ?��K�drL@�+#�%" %��|T0 k� �do�ho%�@c  I%1t'2Q  ��    �  AS)D�URk�P��|$ ?��K�drL@�,#�&!�%��|T0 k� �do�ho%�@c  I%1t'2Q  ��    �  AS)D�ARg�P��|$ ?��K�drL@�,#�&!�%��{T0 k� �do�ho%�@c  I%1t'2Q  ��    �  AS(D�ARg�P��|$ ?��K�drL@�-#�&!�%��{T0 k� �do�ho%�@c  I%1t'2Q  ��    �  AS(D�ARg�P��|$ ?��K�drL@�.#�'!�%��{T0 k� �`o�do%�@c  I%1t'2Q  ��    �  AS(D�ARg�P{��|$ ?��K�drL0�/#�'!�%��zT0 k� �`o�do%�@c  I%1t'2Q  ��    �  AS(D�ARg�P{��|$ ?��K�drL0�0#�(!�%��zT0 k� �`o�do%�@c  I%1t'2Q  ��    �  AS(D�ARc�P{��|$ ?��K�drL0�1#�(!�%��yT0 k� �`o�do%�@c  I%1t'2Q  ��    �  AS(D�ARc�P{��|$ ?��K�`rL0�1#�(!�%��yT0 k� �`o�do%�@c  I%1t'2Q  ��    �  AS'D�ARc�P{��|$ O��K�`rL0�2#�)!�%��xT0 k� �`o�do%�@c  I%1t'2Q  ��    �  AS'D�ARc�P{�ߛ|$ O��K�`rL0�3#�)!�%��xT0 k� �`o�do%�@c  I%1t'2Q  ��    �  AS'D�ARc�P{�ߛ|$ O��K�`sD0�4#�)!�%��xT0 k� �`p�dp%�@c  I%1t'2Q  ��    �  AS'D�ARc�P{�ߛ|$ O��K�`sD0�5#�*!�&��wT0 k� �`p�dp%�@c  I%1t'2Q  ��    �  AS 'D�AR_�P{�ۛ|$ O��K�`sD0�5�*!�&��wT0 k� �\p�`p%�@c  I%1t'2Q  ��    �  AS 'D�AR_�P{�ۛ|$ O��K�`sD0�6�*!�&��vT0 k� �\p�`p%�@c  I%1t'2Q  ��    �  AS &D�AR_�P{�ۛ|$ O��K�`sD0�7�+�&��vT0 k� �\p�`p%�@c  I%1t'2Q  ��    �  AR�&D�AR_�P{�ל|$ O�K�`sD0�8�+�&��vT0 k� �\p�`p%�@c  I%1t'2Q  ��    �  AR�&D�AR_�P{�ל|$ O{�K�`sD0�9�+�&��uT0 k� �\q�`q%�@c  I%1t'2Q  ��    �  AR�&D�AR_�P{�ל|$ Ow�K�\sD0�:�,�&��uT0 k� �\q�`q%�@c  I%1t'2Q  ��    �  AR�&D�AR_�Pw�Ӝ|$ ?s�K�\sD0�;�,�&��uT0 k� �\q�`q%�@c  I%1t'2Q  ��    �  AR�&D�AR[�Pw�Ӝ|$ ?o�K�\sD0�<�,�&��tT0 k� �\q�`q%�@c  I%1t'2Q  ��    �  AR�&D�AR[�Pw�Ӝ|$ ?o�K�\sD0�=�-��&��tT0 k� �\q�`q%�@c  I%1t'2Q  ��    �  AR�%D�AR[�Pw�Ϝ|$ ?k�K�\sD0�>�-��&��tT0 k� �\q�`q%�@c  I%1t'2Q  ��    �  AR�%D�AR[�Pw�Ϝ|$ ?g�K�\sD@�?�-��&��sT0 k� �Xq�\q%�@c  I%1t'2Q  ��    �  AR�%D�AR[�Pw�Ϝ|$ ?c�K�\sD@�@�.��&��sT0 k� �Xq�\q%�@c  I%1t'2Q  ��    �  AR�%D�AR[�Pw�ϝ|$ ?c�K�\sD@�A�.��&��sT0 k� �Xq�\q%�@c  I%1t'2Q  ��    �  AR�%D�AR[�Pw�˝|$ ?_�K�\sD@�B�.��&��rT0 k� �Xq�\q%�@c  I%1t'2Q  ��    �  AR�%D�ARW�Pw�˝|$ ?[�K�\sD@�C�.�&��rT0 k� �Xq�\q%�@c  I%1t'2Q  ��    �  AR�%D�ARW�Pw�˝|$ ?[�K�\sD@�E�/�&��rT0 k� �Xq�\q%�@c  I%1t'2Q  ��    �  AR�%D�ARW�Pw�˝|$ /W�K�\sD@�F�/�& �rT0 k� �Xq�\q%�@c  I%1t'2a  ��    �  AR�$D�ARW�Pw�ǝ|$ /S�K�XsD@�G�|/�& SxT0 k� �Xq�\q%�@c  I%1t'2a  ��    �  AR�$D�ARW�Pw�ǝ|$ /S�K�XsI��H�|/A�&�SxT0 k� �Xq�\q%�@c  I%1t'2a  ��    �  AR�$D�ARW�Pw�ǝ|$ /O�K�XsI��I�x0A�&�SxT0 k� �Xq�\q%�@c  I%1t'2a  ��    �  AR�$D�ARW�Pw�ǝ|$ /O�K�XsI��J�t0A�&�SxT0 k� �Xq�\q%�@c  I%1t'2a  ��    �  AR�$D�ARW�Pw�Ý|$ /K�K�XsI��K�p0A�&�SxT0 k� �Xq�\q%�@c  I%1t'2a  ��    �  AR�$D�ARS�Pw�Ý|$ /K�K�XsI��L�p0A�'�SxT0 k� �Xq�\q%�@c  I%1t'2a  ��    �  AR�$D�ARS�Pw�Þ|$ /K�K�XsI��M�l1A�'�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�$D�ARS�Pw�Þ|$ /K�K�XsI��N�h1A�'�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�$D�ARS�Ps���|$ /G�K�XsI��O�d1A�(�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�$D�ARS�Ps���|$ �G�K�XsI��O�`1A�(�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�#D�ARS�Ps���|$ �G�K�XsI��P�\2A�(�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�#D�ARS�Ps���|$ �G�K�XsI��P�X2�|)�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��   �  AR�#D�ARS�Ps���|$ �G�K�XsI��QT2�x)�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�#D�ARS�Ps���|$ �G�K�XsI��RL2�t*�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�#D�ARS�Ps���|$ �G�K�XsI��RH3�p*�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�#D�ARO�Ps���|$ �G�K�TsI��RD3�h+�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�#D�ARO�Ps���|$ �G�K�TsI��S@3�d,�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�#D�ARO�Ps���|$ �K�K�TsI��S83�\,�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�#D�ARO�Ps���|$ �K�K�TsI��S43�X-�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�#D�ARO�Ps���|$ �K�K�TsI��T04�P.�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�#D�ARO�Ps���|$ �K�K�TsI��T(4�L/�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�"D�ARO�Ps���|$ O�K�TsI��T$4�H/�SxT0 k� �Tq�Xq%�@c  I%1t'2a  ��    �  AR�"D�ARO�Ps���|$ O�K�TsI��T4�@0�SxT0 k� �Pq�Tq%�@c  I%1t'2a  ��    �  AR�"D�ARO�Ps���|$ S�@oTsI��T4�81�SxT0 k� �Xm�\m%�@c  I%1t'2a  ��    �  AR�"D�ARO�Ps���|$ S�@oTsI��T5�42�SxT0 k� �\j�`j%�@c  I%1t'2a  ��    �  AR�"D�ARO�Ps���|$ S�@oTsI��T5�,3�SxT0 k� �`h�dh%�@c  I%1t'2a  ��    �  AR�"D�ARK�Ps���|$ W�@oTsI��T5�(4�SxT0 k� �df�hf%�@c  I%1t'2a  ��    �  AR�"D�ARK�Ps���|$ [�@oTtA��T 5� 5�SxT0 k� �he�le%�@c  I%1t'2a  ��    �  AR�"D�ARK�Ps���|$ [�@oTtA��T�5�6�SxT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�"D�ARK�Ps���!�$ _�@oTtA��T�5�7�SxT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�"D�ARK�Ps���!�$ _�@oTtA��T�6�8�SxT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�"D�ARK�Ps���!�$ c�@oTtA��T�6�9�SxT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�"D�ARK�Ps���!�$ g�@oTtA��T�6� :�SxT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�"D�ARK�Ps���!�$ h @oTtA��T�6��;�SxT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARK�Ps���!�$ h@oTtA��T��6��<�SxT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARK�Ps���!�$ l@oPtA��T��6��=�SxT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARK�Ps���!�$ p@oPtA��T��7��>�SxT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARK�Po���!�$ �t	@oPtAP�T�7��A�SxT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARK�Po���!�$ �x@oPtAP�T�7	p�B�SyT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARK�Po���|$ �x@oPtAP�T�7	p�CQSzT0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���|$ �|@oPtAP�T�7	p�DQS{T0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���|$ ��@oPtAP�T�7	p�DQS|T0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���|$ ��@oPtAP�U�8	p�DQS}T0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���|$ ��@oPtAP�U�8	��DQS~T0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���|$ ��@oPtAP�V�x8	��DQST0 k� �hd�ld%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���|$ ��@oPtAP�V�p8	��DQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���|$ ό@oPtAP�V�h8	��DQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���|$ ό@oPtAP�W�`8	��DQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���|$ ϐ@oPtAP�W�X8@�DQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���|$ ϐ@oPtAP�W�P9@�DQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR�!D�ARG�Po���!�$ ϔ @oPtAP�W�H9@�EQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARG�Po���!�$ ϔ!@oPtAP�W�@9@�EQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARG�Po���!�$ Ϙ#@oPtAP�X�89@�EQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARG�Po���!�$ Ϙ$@oPtAP�X�09@�EQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARG�Po���!�$ Ϝ%@oPtAP�X�(9@�FQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARG�Po���!�$ Ϝ'@oPtAP�X�90�FQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARG�Po���!�$ Ϡ(@oPtAP�X90�FQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARG�Po���!�$ Ϡ*@oPtAP�X90�GQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARG�Po���!�$ Ϥ+@oPtAP�X:0�GQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���!�$ Ϥ,@oPtAP�X�:0�HQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���!�$ Ϩ.@oPtAP�X�:0|HQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ Ϩ/@oPtAP�X�:0xIQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ Ϭ0@oPtAP�X�:0tJQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ Ϭ2@oPtAP�X�:�pJQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ϰ3@oPtAP�X�:�lKQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ϰ4@oPtAP�X�:�hLQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ϴ5@oLtAP�X�:�dLQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ϴ6@oLtL�X�;�dMQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ϴ8@oLtL�X�;�`NQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ϸ9@oLtL�X�;�\NQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ϸ:@oLtL�X�;�XOQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ϼ;@oLtL�X�;�TPQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ϼ<@oLtL�XA�;�TPQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ϼ=@oLtL�XA�;�PQQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ��>@oLtL�XA�;�LQQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ��?@oLtL�XA|<�HRQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR� D�ARC�Po���|$ ��@@oLtL�XAt<�HSQS�T0 k� �dd�hd%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��AK�LtL�X�l<�DSQS�T0 k� �\h�`h%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��BK�LtL�X�d<�@TQS�T0 k� �Xk�\k%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��CK�LtL�X�\<�<TQS�T0 k� �Tm�Xm%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��DK�LtL�X�T<�<UQS�T0 k� �Pn�Tn%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��EK�LtL �X�L=�8UQS�T0 k� �Lo�Po%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��FK�LtL �X�D=�4VQS�T0 k� �Lp�Pp%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��GK�LtL �X�<=�4VQS�T0 k� �Lq�Pq%�@c  I%1t'2a  ��   �  AR�D�ARC�Po���|$ ��HK�LtL �X�8=�0WQS�T0 k� �Lq�Pq%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��IK�LtL �X�0=�,WQS�T0 k� �Lq�Pq%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��JK�LtL �X�(>�,XQS�T0 k� �Lq�Pq%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��KK�LtL �X�$>�(XQS�T0 k� �Lq�Pq%�@c  I%1t'2a  ��    �  AR�D�ARC�Po���|$ ��KK�LtL �X�>�(YQS�T0 k� �Lq�Pq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��LK�LtL �X�>�$YQS�T0 k� �Lq�Pq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��MK�LtL �X>� ZQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��NK�LtL �X>� ZQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��OK�LtL �X >�[QS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��PK�LtL �X �?�[QS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��PK�LtL �X �?�\QS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��QK�LtL �X �?�\QS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��   �  AR�D�AR?�Po���|$ ��RK�LtL �X �?�\QS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��RK�LtL �X �?�]QS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ /�SK�LtL �X �?�^QS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ /�SK�LtL �X �@�_QS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ /�TK�LtL �X �@�_QS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ /�UK�LtL �X �@�`QS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ /�VK�LtL �X �@�aQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ �VK�LtL �X �@�aQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ �WK�LtL �X �@�bQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ �XK�LtL �X �@�cQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ �YK�LtL �X �@�cQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ �YK�LtL �X �A�dQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��ZK�LtL �X �A�eQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��ZK�LtL �X �A�fQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��[K�LtL �X �A�fQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��[K�LtL �X �A�gQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��[K�LtL �X �A�hQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��\K�LtL �X �A�iQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��\K�LtL �X �A�jQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��]K�LtL �X �A�jQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��]K�LtL �X �B�kQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��]K�LtL �X �B�lQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��^K�LtL �X �B�lQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��^K�LtL �X |B�mQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��_K�LtL �X xB�nQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��_K�LtL �X tB�nQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ ��_K�LtL�X pB�oQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ � _K�LtL�X lB�pQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ _K�LtL�X hB0qQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ `K�LtL�X dB0 qQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ `K�LtL�X `C0 rQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ `K�LtL�X \C0 sQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��   �  AR�D�AR?�Po���|$ aK�LtAP�X XC0 sQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ �aK�LtAP�X TC $sQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ � aK�LtAP�X PC $sQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ �$aK�LtAP�X�PC $rQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ �(aK�LtAP�X�LC (rQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ �,aK�LtAP�X�HC (rQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�0aK�LtAP�X�DC�(rQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�4aK�LtAP�X�@C�,rQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�8aK�LtAP�X�@C�,rQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�<aK�LtAP�X�<D�,qQS�T0 k� �Hq�Lq%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�@a@oLtAP�X�8D�,qQS�T0 k� �Pm�Tm%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 
 Da@oLtAP�X�4D�0qQS�T0 k� �Tj�Xj%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 
 Ha@oLtAP�X�0D�0qQS�T0 k� �Xh�\h%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 
 Ha@oLtAP�X�,D�0qQS�T0 k� �\g�`g%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 
 La@oLtAP�X�(E�4qQS�T0 k� �`f�df%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 
 Pa@oLtAP�X�$E�4qQS�T0 k� �`e�de%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�Pa@oLtAP�X� E�4pQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�Ta@oLtAP�X@F�4pQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�Ta@oLtAP�X@F�8pQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�Xa@oLtAP�X@G�8pQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�Xa@oLtAP�X@G�8pQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 
 Xa@oLtL�X@H�8pQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 
 \a@oLtL�X@H�<pQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 
 \a@oLtL�X@I�<oQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 
 \a@oLtL�X� I�<oQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 
 \a@oLtL�X��J�<oQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�`a@oLtL�X��J�@oQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  AR�D�AR?�Po���|$ 	�`a@oLtL�X��K�@oQS�T0 k� �`d�dd%�@c  I%1t'2a  ��    �  D߰�E��ޤA�	|$ PG�E���E�L% ��0�-3� T0 k� ����%�@c  I%1t'2Q  ��    �   HD߰ �E��ޠB�	|$ PG�E���E�T& ��0�.3� T0 k� ����%�@c  I%1t'2Q  ��    �   JD߰ �E��ޘC�
|$ PG�E���E�\'0��0�.3� T0 k� ����%�@c  I%1t'2Q  ��    �   LD߰!�E��ޔC�
|$ @G�E���E�d(0��1 /3� T0 k� ����%�@c  I%1t'2Q  ��    �   ND߰! E��ސD�
|$ @G�E���E�l)0��1 03� T0 k� �#��'�%�@c  I%1t'2Q  ��    �   PD߰"B��ތE�|$ @G�E���E�p*0��! 13� T0 k� �'��+�%�@c  I%1t'2Q  ��    �   RD߰#B��ވE�|$ @G�E���E�x,0��!23� T0 k� �, �0 %�@c  I%1t'2Q  ��    �   UD�#B��ބF�||$ @G�E���E��-0��!33� T0 k� �4�8%�@c  I%1t'2Q  ��    �   XD�$B���|G�x|$ @G�E���E��.0��!43� T0 k� �<�@%�@c  I%1t'2Q  ��    �   [D�%(B���tH�p|$ 0G�E��E��00��!73� T0 k� �H�L%�@c  I%1t'2Q  ��    �   ^D�&,B���pI�l|$ 0G�E���E��10��!83� T0 k� �P�T%�@c  I%1t'2Q  ��    �   aD�'4B���lI�h|$ 0G�E���E��20��!93� T0 k� �T�X%�@c  I%1t'2Q  ��    �   dD�(8B���hJ�d|$ 0K�E���E��30��!:3� T0 k� �\�`%�@c  I%1t'2Q  ��    �   gD�)@B���dK�`|$ 0K�E���E��30��!;3� T0 k� �`�d%�@c  I%1t'2Q  ��    �   jD��*DB���`K�\|$  `K�E���E��40��!=3� T0 k� �d�h%�@c  I%1t'2Q  ��    �   mD��+LB���\L�X|$  `K�E���E��50��>3� T0 k� �d	�h	%�@c  I%1t'2Q  ��    �   pD��,TB���XL�T|$  `O�E���E��60��?3� T0 k� �h�l%�@c  I%1t'2Q  ��    �   sD��,XB���TM�P|$  `O�E���E��60�� @3� T0 k� �l�p%�@c  I%1t'2Q  ��    �   vD��-`B���PN�L|$  `O�E���E��70��$A3� T0 k� �t�x%�@c  I%1t'2Q  ��    �   yD��0�lB���HO�D|$  S�F��E��80��(D3� T0 k� ����%�@c  I%1t'2Q  ��    �   }D��1�tB���DO�@|$  W�F��B��90���,E3� T0 k� ����%�@c  I%1t'2Q  ��    �   �F�2�|B���@P�<|$  [�F��B��90���4F3� T0 k� ����%�@c  I%1t'2Q  ��    �   �F�3��B���<P�8|$  _�F��B� 90���8G3� T0 k� ����%�@c  I%1t'2Q  ��    �   �F�4��B���<P�4|$  _�F�B�:0���<H3� T0 k� ����%�@c  I%1t'2Q  ��    �   �F�5��B���8Q�0|$ c�F{�B�:0���@I3� T0 k� ����%�@c  I%1t'2Q  ��    �   �F�6��B���4Q�,|$ g�Fw�E�:0���DJ3� T0 k� ����%�@c  I%1t'2Q  ��    �   �E��7��B���4Q�(|$ k�Fw�E�;0���LK3� T0 k� ����%�@c  I%1t'2Q  ��    �   �E��9��B�#��0R�(|$ o�E�s�E�$;0���PL3� T0 k� ����%�@c  I%1t'2Q  ��    �   �E��:��B�'��0R$|$ s�E�s�E�,;0���TM3�T0 k� ��	��	%�@c  I%1t'2Q  ��    �   �E��;��B�+��,R |$ �w�E�o�E�4;0���\N3�T0 k� ����%�@c  I%1t'2Q  ��   �   �E��<��B�/��,R|$ �{�E�l E"<;0���`O3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B��=��B�3��(R|$ ��E�l E"D;0���hP3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B��>��B�7��(R|$ ���B�lE"L;0���lQ3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B� ?��B�;��(R|$ ���B�hE"T;0���tR3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B�@Q�B�?��(R�|$ ���B�hE"\;1��xS3�T0 k� ����%�@c  I%1t'2Q  ��    �   �B�AQ�B�C��$R�|$ ���B�hE"d;1���T3�T0 k� ��� %�@c  I%1t'2Q  ��    �   �B�BQ�B�G��$R�|$ ���B�hE"l;1���U3�T0 k� �	�	%�@c  I%1t'2Q  ��    �   �B�CQ�B�O��$R�|$ ���B�hE�t;1���V3�T0 k� �
�
%�@c  I%1t'2Q  ��    �   �B�DR B�S��$R�|$ ���B�lE�|;1���W3�T0 k� �
�
%�@c  I%1t'2Q  ��    �   �B� ERB�W��$R�|$ ���B�lE��;1���W3�T0 k� � 
�$
%�@c  I%1t'2Q  ��    �   �B�$FRB�[��$R�|$ ���B�lE��:1���X3�T0 k� �(	�,	%�@c  I%1t'2Q  ��    �   �B�,G�B�c��$R�|$ ���B�lE��:1���Y3�T0 k� �0�4%�@c  I%1t'2Q  ��    �   �B�0H�$B�g��$R�
|$ ���B�pE��:1���Z3�T0 k� �8�<%�@c  I%1t'2Q  ��    �   �B�8I�,B�o��$R�
|$ �ǸB�pE��:1���[3�T0 k� �@�D%�@c  I%1t'2Q  ��    �   �B�<J�4B�s��$R�	|$ �˸B�tE��91���\3�T0 k� �H�L%�@c  I%1t'2Q  ��    �   �B�DJ�<B�{��$R�	|$ �ӹB�tE��91���\3�T0 k� �P�T%�@c  I%1t'2Q  ��    �   �B�HK�DB���$R�	|$ �۹B�xE��91���]3�T0 k� �T�X%�@c  I%1t'2Q  ��    �   �B�PL�LBЇ��$R�|$ �߹B�|E��81���^3�T0 k� �\�`%�@c  I%1t'2Q  ��    �   �B�XM�TB����$R�|$ ��B�|	E��81���_3�T0 k� �d�h%�@c  I%1t'2Q  ��    �   �B�\N�\B����$R�|$ ��B��	E��71���_3�T0 k� �l�p%�@c  I%1t'2Q  ��    �   �B�dO�`B����$R�|$ ���B��	E��71���`3�T0 k� �p�t%�@c  I%1t'2Q  ��    �   �B�lO�hB���N$R�|$ ���B��
E��61���a3�T0 k� �x�|%�@c  I%1t'2Q  ��    �   �B�pP�pB���N$R�|$ ��B��
E��51�� a3�T0 k� �|��%�@c  I%1t'2Q  ��    �   �                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \���� ]�'�'� ` � �S         � �n�     � �r�    ����                  >          �p     ���   0
% 
          ����   $/
    ���    ������                       	    �8          �     ���  0
 	         ���I         �0(    ���I �1      ��               	   �         p     ���   8	          �ϻ-           �    �ϻ- �                        �$          ��     ���   8         ��Ԓ           .����    ���@����     2��               
  �$          �     ���   P
	
           �^  ��     B�	��      �^�	��                             ���              �  ���    P              a�8  � �    V �     a�8 K       �             	 Z          ���     ��@  (
I  
          ty       j��@)     ty��@)                  V  Z           �      ��H   8	            XS � � 
	   ~ *X     XS *X                   ]	 Z           �     ��`   P	
           K�%  � �	    ���*      J���8�    .�            R  Z          	 &0�   	  ��` Pw           op�  � �
	   � X�     o�P q    �3o            G Z          
 � �    ��`@  
2	         ����          � T�    ���� T�    �                  	 d�p P _               ��B   0
	 	               ��      �                                                                           �                               ��        ���          ��                                                                 �                          dO8  ��        ��ب      dO8�ب          "                 x                j  �       �                          d    ��        ���       d  ��           "                                                �                          � � ���	 �� *��  T������    	     
        
  G    � �� j��A       � j� �$ `j� �� @k� �d l  �� t  �� q@ � u� �$  v  �d v@ �� v` �� s@ �� 0s` �D  s� �� t  �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀���� ����� ����� ����� ����� � 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����   ����  ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    $�j � ��$  �
� �  �  
�  t    ��     ���           ��     � �       t    ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �%      �� �  ��        �t �  ���        �        ��        �        ��        �    ��     j�� j��        ��                         �w� $ �� �                                    �                 ����             t�� ���%��    ��                 32 Don Sweeney son     5:42                                                                        5  5      � �
"� �SC. kC6 �#kjO1kr?/ �E. �D �c�& � 	c�5 �
c�5c�5 � c�( �c�I � c�I � c�Y �c�Y � c�Q � c�N � V9 �	cW9 �c]A � ca1 �C � � C" � �k~0 � k�8 �c� � � c� � jK � � K � MJ� � m  J� �F!"�LF ""�^6#�H6$
�W m%"� � m &"� ]'"� � ](*�F)"�LF *"�^6+�H6 
�W6-�H6 
�WF/"�LF 0"�^61�H6 
�W6 
�W
 
�}5"�q 6"��7�m 
�|9�l 
�{ ~  *Gr �  *NW � =*@ �  *NX �  *NY                                                                                                                                                                                                                         �� R   �     �    @ 
       �     ] P E ^  ��                    	 �������������������������������������� ���������	�
��������                                                                                          ��    �GG�� ��������������������������������������������������������   �4, h� * � ���A������9� ���� ��                                                                                                                                                                                                                                                                                                                                '"(�@��                                                                                                                                                                                                                                     	         '    � �  D�J    	  ^�  	                           ������������������������������������������������������                                                                       
                                                                    u           �        �       �  �          	  
 	 
 	 	 ����������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� �������������������            �           
     V  
  %      �  	f�J �    L�                             ������������������������������������������������������                                                                    	                                                            	       �       ��        �          � �              	   	 	 �������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ����             x                                                                                                                                                                                                                                                           
                                                 �             


          �   }�    �    ��������������������������������  +����������������  '�  'q������������  +	����������������������������                                     '�                                           �ww�ww333wwwwwwww�ww�ww�ww�ww333wwww 0 I =               	                  � q�� �j�                                                                                                                                                                                                                                                                                   )n)n1n  
�              a      `      l      k                  m                                                                                                                                                                                                                                                                                                                                                                                                        � � �  � ��  � ��  � @��  � (��  � ��  �����|�����������������i�����Q�����������T�����8                 z � : v��        	 	 �   & AG� �  �   
              �                                                                                                                                                                                                                                                                                                                                      p B L    �      ��               !��                                                                                                                                                                                                                            Y��   �� � ���      �� @ 	 �� 
����������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� ��������������������������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ����             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    3      2      d                       B     �  �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$     `d     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@     \ 
pn ��  \ 
pn �$ ^$   L j� � �� j� � �$ /  ��/       �   d   5���� e�����  g��� 	 �     f ^�   `     ��v       5      ���
���2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                                                �����   �   �   �   ����                                     
�  

  
 � 
 
 
   
   
   
   
  ��                  ��   
   
   
   
   
   
 
 
 � 

  
�                 �   
    �   
    �   
    �   
   
   �  
   �  
   �  
   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "  "!  "" "  """           """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """""" "!   " ""  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  "!  "" "  """           """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��      �    �  �   �����������    ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                 � �� ��  ��                                                                                                                                                                                                �UCD�UTE
EUT �T8 �D�  ��  �  �   �   �      �  �  �� �� ��EO  TO  C�� ��� ��� ������̻�̻�̻�w˙�b��v&���}��ۻ����ȯ����                       �ϻ��̋��̨���z������ ��  ��  ��  ��  �                           ��  "   "/  ./� "�� �   �   ��     �                    �   ��  �  �   ��  �  �  �� �� ��  �� �,� �"/�""�"/� "/  �         "  "  ""  "+� �� � ��   �  "   "�  +�  
�� ��� D�D 4ETO3    �   �   �   D   E�  U�  UO                         "  "  "                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��               �   �   �  �  �  �  �   �   �                                       �  ���   �                          �   �   ��� ������ �   �      �       �                        �   ��  ���  � �    �               � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                       �  ��  ��  ww  ��  vv  w"   "   "  �� ��                   ����������                          �  �� ��  �    � ���                                                                                                                                                                                                           �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �        �  ��  ��  ww  ��  vv  w"   "   "  �� ��                   ����������                          �  �� ��  �    � ���                                       �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                                 �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                                 1    1   "    �   �   �� �����  �    �   �   ,   "   "                   ���ۼ����� 9��C��UTDD�D33��0��  "��
/� � �, �"  �"   �   ˻ڛ��Ȱ��  ��  ��  TJ  EJ  DT  4E  �P  ��  �   /   ��  ��� �                                     � 	�� �� �˙	���
������                Ͱ  ˻  ˻  ۻ  ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                  �   �   �   �   �      �                    ��� ���� ��    ��   �  ��  �  �  �         � �������������  �                                                                                                                                                              	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                   "   "   "       �         �        �   �     �       �   �   �   �   �      �                    ��� ���� ��             �  �˰ ��� �wp ���                                                                                                                                                                   �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw  ��  �   ��  �                                   � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                          w 
�� ɚ� ���
�˻Ɋ�����������-� �"+ ". "$ "$ �U  Z�  Z�  J�  J�  �D  ��  ��  ɘ ˰ "  �"/�"" "  �  �            g���z��ȩ�����ة�� ���  ̰  ̰  ˰  ��  �  N�� T4�CD  CD0 C40 C30 3;� ܰ �� �� �  �  "  �""�"" �"/���  � �  �      �     �   �   ��  �"" �""  ""   "                 �   ��   �                            � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                                                                                                                                                                "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��             �  �˰ ��� �wp ���      � �������������  �                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��   +� �".  ���  � ��  �       ��������  �� �""����� � �  � � �     �   �                     �   �                     �     �                                      � ����ݼ� ����     �   �   �   �   �   �                                                                                                                                                �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwwDwwAwwA""""wwwwwwqADDGG""""wwwwwwqAqwAwG""""wwwwDDtwwwww""""wwwwwqGDADGqGGqw""""wwwwwwDqGqG""""wwwwwwwwwwwwqwwqww""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUEUUEUUUUUUTDUUUU3333DDDDAEQQDUDEUTUUUU3333DDDDUETQEUADQDEUDUUUU3333DDDDUQUUDUDEUTUUUU3333DDDDEQUEQUEUEUQEUUDUUUU3333DDDDQEEDEEEDUTEUUUU3333DDDDQUUQUUQUUQUUUDUUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
"� �SC. kC6 �#kjO1kr?/ �E. �D �c�% � 	c�5 �
c�5c�5 � c�( �c�I � c�I � c�Y �c�Y � c�Q � c�N � V9 �	cW9 �c]A � ca1 �C � � C" � �k~0 � k�8 �c� � � c� � jK � � K � MJ� � m  J� �F!"�LF ""�^6#�H6$
�W m%"� � m &"� ]'"� � ](*�F)"�LF *"�^6+�H6 
�W6-�H6 
�WF/"�LF 0"�^61�H6 
�W6 
�W
 
�}5"�q 6"��7�m 
�|9�l 
�{ ~  *Gr �  *NW � =*@ �  *NX �  *NY3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������+�J�G�S���G�Z�K�Y� � � � � � � � � � �,��<�����������������������������������������$��4�U�K��4�[�T�K�G�[� � � � � � � � � � �,��<�������������������������������������������.�U�T��<�]�K�K�T�K�_� � � � � � � � � �,��<�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,��<� �� �������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                