GST@�                                                            \     �                                               d  �   ��                   ���2�����	 J���������������z���        �h     #    z���                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    
 �j
  ����
��
�"     "�j��   * ��
                                                                                 ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             �E  "          == �����������������������������������������������������������������������������                                ��  �   �   �   @  #   �   �                                                                                '       )n)n1n  �"E    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�9O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE & �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    I@/���@����,� |( P3��@@ E���@�3� T0 k� �4
�8
Y"t'!"t1'   ��'   �  I@/���@����,� |( P/��@@ E���@�3� T0 k� �4
�8
Y"t'!"t1'   ��'   �  I03���@����,� |( P/��@@ E���@�3� T0 k� �4
�8
Y"t'!"t1'   ��'   � ��I03���@����, |( P+��D@ E���@�3� T0 k� �4
�8
Y"t'!"t1'   ��'   � ��I03���@����-$|( P'��D@ E���@�3� T0 k� �8	�<	Y"t'!"t1'   ��'   � ��I07���@����-$|( P#��D@ E���P��3� T0 k� �8	�<	Y"t'!"t1'   ��'   � ��I@7���@����-$|( P��D@ J��P��3� T0 k� �8�<Y"t'!"t1'   ��'   � ��I@7�� @�� n�-o(|( ���D@ J��P��3� T0 k� �8�<Y"t'!"t1'   ��'   � ��I@7��@�� n�-o(|( ���D@ J��P��3� T0 k� �8�<Y"t'!"t1'   ��'   � ��I@7��@�� n�-o(|( ���D@ J��P��3� T0 k� �8�<Y"t'!"t1'   ��'   � ��I@7��@�� n�.o(|( ���D@ J��P��3� T0 k� �8�<Y"t'!"t1'   ��'   � ��I07� @�� n�.o(|( ���D@ J��P��3� T0 k� �8�<Y"t'!"t1'   ��'   � ��I07� @�� ��._(|( P��D@ J�#�
п�3� T0 k� �8�<Y"t'!"t1'   ��'   � ��I07� @�� ��._(|( P��D@ J�'�
п�3� T0 k� �8�<Y"t'!"t1'   ��'   � ��I07� @�� ��._(|( _���H@ J�/�
���3� T0 k� �8�<Y"t'!"t1'   ��'   � ��I07� @�� ��._(|( _���H@ J�3�
���3� T0 k� �<�@Y"t'!"t1'   ��'   � ��I@7� @�� ��._(|( _���H@ J�;�
���3� T0 k� �<�@Y"t'!"t1'   ��'   � ��I@7� @���.?(|( _���H@ J�C�
���3� T0 k� �<�@Y"t'!"t1'   ��'   � ��I@7� @���.?$|( _���H@ J�G�
���3� T0 k� �<�@Y"t'!"t1'   ��'   � ��I@7� @���.?$|( _���H@ J�O�
���3� T0 k� �<�@Y"t'!"t1'   ��'   � ��I@7� @���.?$|( O���H@ J�W�
���3� T0 k� �<�@Y"t'!"t1'   ��'   � ��@`7� @���/?$|( O���H@ J�_�
���3� T0 k� �<�@Y"t'!"t1'   ��'   � ��@`7�@���/o$|( O���H@ J�c�
���3� T0 k� �<�@Y"t'!"t1'   ��'   � ��@`7�@���/o$|( O���H@ E�k�
���3� T0 k� �<�@Y"t'!"t1'   ��'   � ��@`7�@���/o$|( O���H@ E�s�@��3� T0 k� �<�@Y"t'!"t1'   ��'   � ��@`7�@���/o$|( ����H@ E�w�@��3� T0 k� �<�@Y"t'!"t1'   ��'   � ��@7�@���0o$|( ����H@ E��@��3� T0 k� �<�@Y"t'!"t1'   ��'   � ��@7� `@��~�0
$|( ����H@ Eу�@��3� T0 k� �<�@Y"t'!"t1'   ��'   � ��@7� `@��~�0
$|( ����H@ E��@��3� T0 k� �<�@Y"t'!"t1'   ��'   � ��@7� `@��~�1
$|( ����L@ E��@��3� T0 k� �<�@Y"t'!"t1'   ��'   � ��@7� `@��~�1
 |( ����L@ E��@��3� T0 k� �@�DY"t'!"t1'   ��'   � ��@7� `@��~�2
 |( ����L@ E��A�3� T0 k� �@�DY"t'!"t1'   �'    � ��@7� @����2� |( ���L@ E��A�3� T0 k� �@�DY"t'!"t1'   �'    � ��@7� @����3�|( ���L@ A���A�3� T0 k� �@�DY"t'!"t1'   ��'    � ��@7� @����3�|( ���L@ A����3� T0 k� �@�DY"t'!"t1'   ��'    � ��@7� @����4�|( ���L@ A����3� T0 k� �@�DY"t'!"t1'   ��'    � ��B@7� @����4�|( ���L@ A����3� T0 k� �@�DY"t'!"t1'   ��'    � ��B@7� `@��~�4 o|( ��L@ A����3� T0 k� �@�DY"t'!"t1'   ��'    � ��B@7� `@��~�5 o|( w��L@ A����3� T0 k� �@�DY"t'!"t1'   ��'    � ��B@7� `@��~�5 o|( s��L@ A����3� T0 k� �@�DY"t'!"t1'   ��'    � ��B@7� `@��~�6 o|( o��L@ A����3� T0 k� �@�DY"t'!"t1'   ��'    � ��B@7� `@��~�6 o|( g��L@ A����3� T0 k� �@�DY"t'!"t1'   ��'    � ��A�7� �@��~�6 o|( c��L@ A����3� T0 k� �@�DY"t'!"t1'   ��'    � ��A�7� �@��~�7� |( _��L@ A����3� T0 k� �@�DY"t'!"t1'   ��'    � ��A�7� �@��~�7� |( W��L@ A���#�3� T0 k� �@�DY"t'!"t1'   ��'    � ��A�7� �@��~�8�  |( S��L@ A���#�3� T0 k� �@�DY"t'!"t1'   ��'    � ��A�7� �@��~�8�$ |( O��L@ A���'�3� T0 k� �@�DY"t'!"t1'   ��'    � ��D�7�@@��~�8�$!|( K��P@ A���+�3� T0 k� �@�DY"t'!"t1'   ��'    � ��D�7�@@����9�$!|( G��P@ A���+�3� T0 k� �@�DY"t'!"t1'   ��'    � ��D�7�@@����9�("|( C��P@ A���/�3� T0 k� �D �H Y"t'!"t1'   ��'    � ��D�7�@@����9�("|( ;��P@ A���/�3� T0 k� �D �H Y"t'!"t1'   ��'    � ��D�7�@@����:�,#|( 7��P@ A���3�3� T0 k� �D �H Y"t'!"t1'   ��'    � ��D�7�@@����:�,$|( 3��P@ A���3�3� T0 k� �D �H Y"t'!"t1'   ��'    � ��D�7�@@����:�0$|( /��P@ A���7�3� T0 k� �D �H Y"t'!"t1'   ��'    � ��D�7�@@����;�0%|( +��P@ A���7�3� T0 k� �D �H Y"t'!"t1'   ��'    � ��D�7�P@����;4&|( '��P@ A���;�3� T0 k� �D �H Y"t'!"t1'   ��'    � ��D�7�P	@����;8&|( #��P@ A���;�3� T0 k� �D �H Y"t'!"t1'   ��'    � ��D�7�P	@��� ;8'|( ��P@ A���?�3� T0 k� �D �H Y"t'!"t1'   ��'   � ��D�7�P	@��� <<(|( ��P@ A��?�3� T0 k� �G��K�Y"t'!"t1'   ��'    � ��D�7�P	@��� <@)|( ��P@ A��?�3� T0 k� �G��K�Y"t'!"t1'   ��'    � ��D�7�P	@��� <D*|( ��T@ A��C�3� T0 k� �G��K�Y"t'!"t1'   ��'    � ��D�7�P
@��� =H+|( ��T@ A��C�3� T0 k� �K��O�Y"t'!"t1'   ��'    � ��D�7�P@��� =L,|( ��T@ A��G�3� T0 k� �K��O�Y"t'!"t1'   ��'    � ��D�7�P@��� =L-|( ��T@ A��G�3� T0 k� �K��O�Y"t'!"t1'   ��'    � ��D�7�P@��� =P.|( ��T@ A��K�3� T0 k� �K��O�Y"t'!"t1'   ��'    � ��D�7�P@��� >T/|( ���T@ A��K�3� T0 k� �K��O�Y"t'!"t1'   ��'    � ��D�7�`@���>X0|( ���X@ A��K�3� T0 k� �K��O�Y"t'!"t1'   ��'    � ��D�7�`@���>\1|( ���X@ A��O�3� T0 k� �O��S�Y"t'!"t1'   ��'    � ��D�7�`@���?`2|( ���X@ A��O�3� T0 k� �O��S�Y"t'!"t1'   ��'    � ��D�7�`@���?d3|( ��X@ A�#�S�3� T0 k� �O��S�Y"t'!"t1'   ��'    � ��D�7�`@���?h4|( ��X@ A�#�S�3� T0 k� �O��S�Y"t'!"t1'   ��'    � ��D�7�`@���?�p6|( ��X@ A�'�S�3� T0 k� �O��S�Y"t'!"t1'   ��'    � ��D�7�`@���@�t7|( ��\@ A�+�W�3� T0 k� �O��S�Y"t'!"t1'   ��'    � ��D�7�`K����@�x8|( ��\@ A�+�W�3� T0 k� �S��W�Y"t'!"t1'   ��'    � ��D�7�`K����@�|9|( ��\@ A�/�[�3� T0 k� �S��W�Y"t'!"t1'   ��'    � ��D�7�`K����@��;|( ߱�\@ A�3�[�3� T0 k� �S��W�Y"t'!"t1'   ��'   � ��D�7��K����@��<|( ۰�\@ A�3�[�3� T0 k� �S��W�Y"t'!"t1'   ��'    � ��D�7��K����A��=|( ۰�\@ A�7�_�3� T0 k� �S��W�Y"t'!"t1'   ��'    � ��D�7�� K����A��?|( װ�\@ A�7�_�3� T0 k� �S��W�Y"t'!"t1'   ��'    � ��D�7��"K����A��@|( Ӱ�`@ A�;�_�3� T0 k� �S��W�Y"t'!"t1'   ��'    � ��D�7��#K����A��A|( ϰ�`@ A�;�c�3� T0 k� �W��[�Y"t'!"t1'   ��'    � ��D�7��$K����B��C|( ϯ�`@ A�?�c�3� T0 k� �W��[�Y"t'!"t1'   ��'   � ��D�7��&K����B��D|( ˯�`@ A�C�c�3� T0 k� �W��[�Y"t'!"t1'   ��'    � ��D�7��'K����BߨE|( ǯ�`@ A�C�g�3� T0 k� �W��[�Y"t'!"t1'   ��'    � ��D�7��)K����B߬F|( ǯ�`@ A�G�g�3� T0 k� �W��[�Y"t'!"t1'   ��'    � ��D�7��*K����B߰H|( ï�`@ A�G�g�3� T0 k� �W��[�Y"t'!"t1'   ��'    � ��D�7��+K����CߴI|( ���`@ A�K�g�3� T0 k� �W��[�Y"t'!"t1'   ��'    � ��D�7��,K����C߸J|( ���d@ A�K�k�3� T0 k� �W��[�Y"t'!"t1'   ��'    � ��LP7��.K����C߼K|( ���d@ A�O�k�3� T0 k� �[��_�Y"t'!"t1'   ��'    � ��LP7��/K���C��L|( ���d@ A�O�k�3� T0 k� �[��_�Y"t'!"t1'   ��'    � ��LP7��0K���C��M|( ���d@ A�S�o�3� T0 k� �[��_�Y"t'!"t1'   ��'    � ��LP7��1K���C��N|( ���d@ A�S�o�3� T0 k� �[��_�Y"t'!"t1'   ��'    � ��LP7��2K���D��P|( ���d@ A�W�o�3� T0 k� �[��_�Y"t'!"t1'   ��'   � ��LP7��4K���D��Q|( ���d@ A�W�o�3� T0 k� �[��_�Y"t'!"t1'   ��'    � ��LP7��5K���D��R|( ���d@ A�W�s�3� T0 k� �[��_�Y"t'!"t1'   ��'    � ��LP7��6K���OD��S|( ���d@ A�[�s�3� T0 k� �[��_�Y"t'!"t1'   ��'    � ��LP7��7K���OD��T|( ���h@ A�[�s�3� T0 k� �[��_�Y"t'!"t1'   ��'    � ��LP7��8K���OD��U|( ���h@ A�_�s�3� T0 k� �_��c�Y"t'!"t1'   ��'    � ��LP7��9K���OD��V|( ���h@ A�_�w�3� T0 k� �_��c�Y"t'!"t1'   ��'    � ��LP7��:K���OD��W|( ���h@ A�c�w�3� T0 k� �_��c�Y"t'!"t1'   ��'    � ��LP7��;K��� D��X|( ���h@ A�c�w�3� T0 k� �_��c�Y"t'!"t1'   ��'    � ��LP7��<K��� D��Y|( ���h@ A�c�w�3� T0 k� �_��c�Y"t'!"t1'   ��'    � ��L`7��=K��� D��Z|( ���h@ A�g�{�3� T0 k� �_��c�Y"t'!"t1'   ��'    � ��L`7��>K��� D��Z|( ���h@ A�g�{�3� T0 k� �_��c�Y"t'!"t1'   ��'    � ��L`7��?K��� D��[|( ���h@ A�k�{�3� T0 k� �_��c�Y"t'!"t1'   ��'    � ��L`7��@K����D��\|( ���h@ A�k�{�3� T0 k� �_��c�Y"t'!"t1'   ��'    � ��L`7��AK����D��]|( ���l@ A�k��3� T0 k� �_��c�Y"t'!"t1'   ��'    � ��L`7��BK���� D��^|( ���l@ A�o��3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`7��CK���� E� _|( ���l@ A�o��3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`7��DK����$E� `|( ���l@ A�o��3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`7��EK����(E�`|( ���l@ A�s��3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`7��EK����,E�a|( ���l@ A�s���3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`7��FK����0F�b|( ���l@ A�s���3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`7��GK����0F�c|( ���l@ A�w���3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`7�� HK����4F�d|( ���l@ A�w���3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`4� IK����8G�d|( ���l@ A�w���3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`4� JK����<G�e|( ���l@ A�{���3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`4� JK����@H�f|( ���l@ A�{���3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`4� KK����DH�g|( ���p@ A�{���3� T0 k� �c��g�Y"t'!"t1'   ��'    � ��L`4� LK����HI�g|( ��p@ A����3� T0 k� �g��k�Y"t'!"t1'   ��'    � ��L`4� MK����LJ�h|( ��p@ A����3� T0 k� �g��k�Y"t'!"t1'   ��'    � ��L`4� MK����PJ� i|( {��p@ A����3� T0 k� �g��k�Y"t'!"t1'   ��'    � ��L`4� NK����TK�$i|( {��p@ A�����3� T0 k� �g��k�Y"t'!"t1'   ��'    � ��L`0� OK���XL�$j|( {��t@ A�����3� T0 k� �g��k�Y"t'!"t1'   ��'    � ��L`0	� PK���`L�(k|( w��t@ A�����3� T0 k� �g��k�Y"t'!"t1'   ��'    � ��L`0
� PK���dM�(k|( w��t@ A�����3� T0 k� �k��o�Y"t'!"t1'   ��'    � ��L`0� QK���hN�,l|( w��t@ A�����3� T0 k� �k��o�Y"t'!"t1'   ��'    � ��L`0� RK���lO�,m|( s��t@ A�����3� T0 k� �k��o�Y"t'!"t1'   ��'    � ��L`0� RK���pP�0m|( s��x@ A�����3� T0 k� �k��o�Y"t'!"t1'   ��'    � ��L`0� SK���	?xP�4n|( s��x@ A�����3� T0 k� �o��s�Y"t'!"t1'   ��'    � ��L`,� TK���	?|Q�4n|( o��x@ A�����3� T0 k� �o��s�Y"t'!"t1'   ��'    � ��L`,� TK���	?�R�8o|( o��x@ A�����3� T0 k� �o��s�Y"t'!"t1'   ��'    � ��L`,� UK���	?�S�8p|( o��x@ A�����3� T0 k� �o��s�Y"t'!"t1'   ��'    � ��L`,� UK���	?�S�<p|( k��|@ A�����3� T0 k� �o��s�Y"t'!"t1'   ��'    � ��L`,� V@��	?�T�<q|( k��|@ A�����3� T0 k� �o��s�Y"t'!"t1'   ��'    � ��L`,� W@��	O�T�<q|( k��|@ A�����3� T0 k� �s��w�Y"t'!"t1'   ��'    � ��L`,� W@��	O�U�@r|( k��|@ A�����3� T0 k� �s��w�Y"t'!"t1'   ��'    � ��L`,@ X@��	O�U�@r|( g��|@ A�����3� T0 k� �s��w�Y"t'!"t1'   ��'    � ��L`,O�Y@��	O�U�Ds|( g��|@ A�����3� T0 k� �s��w�Y"t'!"t1'   ��'    � ��L`(O�Y@��	O�V�Ds|( g���@ A�����3� T0 k� �s��w�Y"t'!"t1'   ��'    � ��L`(O�Z@��	?�V�Ht|( c���@ A�����3� T0 k� �w��{�Y"t'!"t1'   ��'    � ��L`(O�[K���	?�V�Ht|( c���@ A�����3� T0 k� �w��{�Y"t'!"t1'   ��'    � ��L`(��\K���	?�W�Lu|( c���@ A�����3� T0 k� �w��{�Y"t'!"t1'   ��'    � ��LP(��]K���	?�W�Lu|( c���@ A�����3� T0 k� �w��{�Y"t'!"t1'   ��'    � ��LP(��^K���	?�W�Lv|( _���@ A�����3� T0 k� �w��{�Y"t'!"t1'   ��'    � ��LP(��_K���	O�W�Pv|( _���@ A�����3� T0 k� �w��{�Y"t'!"t1'   ��'    � ��LP(��`K���	O�W�Pw|( _���@ A�����3� T0 k� �{���Y"t'!"t1'   ��'    � ��LP(��aK���	O�W�Pw|( _���@ A�����3� T0 k� �{���Y"t'!"t1'   ��'    � ��LP$��bK���	O�W�Pw|( [���@ A�����3� T0 k� �{���Y"t'!"t1'   ��'    � ��D�$ ��cK���	O�W�Pw|( [���@ A�����3� T0 k� �{���Y"t'!"t1'   ��'    � ��D�$!��dK���	?�W�Pw|( [���@ A�����3� T0 k� �{���Y"t'!"t1'   ��'    � ��D�$"��fK���	?�W�Tw|( [���@ A�����3� T0 k� �{���Y"t'!"t1'   ��'    � ��D�$#��gK���	?�W�Tx|( [���@ A�����3� T0 k� �{���Y"t'!"t1'   ��'    � ��D�$$��hK���	?�W �Tx|( W���@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��Ep$%��iK���	?�W �Tx|( W���@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��Ep$&��kK���	O�W �Tx|( W���@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��Ep$'��lK���	O�W �Tx|( W���@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��Ep$(��mK���	O�W �Tx|( W���@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��Ep$*��nK���	O�W Tx|( S���@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��Ep$+��oK���	O�W Tx|( S���@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��E` ,��pK��� o�W Tx|( S���@ A�����3� T0 k� �����Y"t'!"t1'   ��'   � ��E` .��rK��� o�W Tx|( S���@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��E` /��sK��� o�W Tx|( S���@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��E` 1��tK��� o�WPTx|( O���@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��E`2��uK��� o�WPTx|( O���@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D04��vK��� �WPTx|( O���@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D05��wK��� �WPTx|( O���@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D07��xK��� �WPTy|( O���@ A�����3� T0 k� ������Y"t'!"t1'   ��'   � ��D08��yK��� �W�Ty|( K��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D0:��zK��� �W�Ty|( K��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D0;��zK��� �W�Ty|( K��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D0=�{K��� �W�Px|( K��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D0?�|K��� �W�Px|( K��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D0@�|K��� �W0Px|( K��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D0B�}K��� �W0Px|( K��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D@D�~K��� �W0Px|( G��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��D@E�~K��� �W0Px|( G��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��DO�I��K���O�W0Lx|( G��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��DO�J��K���O�W0Lx|( G��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�L��K���O�W0Lx|( G��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�N��K���O�W0Lw|( G��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�O��K���O�W0Lw|( C��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�Q��K����W0Lw|( C��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�R�|K����W0Hw|( C��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�T�xK����W0Hw|( C��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�T�tK����W0Hw|( C��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�UpK����W@Hw|( C��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�Wl~K����W@Hw|( C��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�Xh~K����W@Hw|( ?��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�Yd~K����W@Hw|( ?��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�Zd}K����W@Hv|( ?��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��L?�[�`}K����W@Dv|( ?��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�\�\}K�����W@Dv|( ?��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�]�\|K�����W@Dv|( ?��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�_�X|K�����W@Dv|( ?��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�`�T{K�����W@Dv|( ?��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�aTzK�����W@Dv|( ?��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�bPzK�����X@Dv|( ;��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�cPyK�����X@Dv|( ;��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�dLyK�����X@Dv|( ;��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�eLxK�����X@Dv|( ;��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�fHx@����X@@v|( ;��@ A�����3� T0 k� ������Y"t'!"t1'   ��'    � ��LO�gHx@����X@@v|( ;��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�hDw@����X@@v|( ;��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�iDw@����X@@u|( ;��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�j@v@����X@@u|( ;��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�j@vK�����X@@u!�( ;��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�k<uK�����X@@u!�( 7��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�l<uK�����X@@u!�( 7��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�m�8tK�����X@@u!�( 7��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�n�8tK�����X@@u!�( 7��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�o�8tK�����X@<u!�( 7��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�p�4sK�����X@<u!�( 7��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�p�4sK�����X@<u!�( 7��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�q�0rK�����X@<u!�( 7��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�r�0rK�����X@<u!�( 7��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�s�,rK�����X@<u!�( 7��@ A�����"�� T0 k� �����Y"t'!"t1'   ��'    � ��LO�t�,qK�����X@<u|( 7��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�t�,qK�����X@<u|( 7��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�u�(qK�����X@<u|( 7��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�v�(pK�����X@<u|( 3��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�v�(pK�����X@<t|( 3��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�w�$pK�����X@<t|( 3��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�x�$oK�����X@<t|( 3��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�y� oK�����X@<t|( 3��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�y� oK�����X@8t|( 3��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�z� nK�����X@8t|( 3��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�{�nK�����X08t|( 3��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��LO�{�nK�����X08t!�( 3��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'    � ��LO�|�mK�����Y08t!�( 3��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'    � ��LO�|�mK�����Y08t!�( 3��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'    � ��LO�}�mK�����Y08t!�( 3��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'    � ��LO�~�lK�����Y08t!�( 3��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'    � ��L?�~�lK���|Y08t!�( 3��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'    � ��L?��lK���|Y08t!�( 3��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'    � ��L?��lK���|Y08t!�( 3��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'   � ��L?Ԁ�kK���|Y04s!�( /��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'    � ��L?Ԁ�kK���|Y04s!�( /��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'    � ��L?Ԁ�kK���|Y04s!�( /��@ A�����"s� T0 k� �����Y"t'!"t1'   ��'    � ��L?��kK���|Y00s|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��L?��jK���xY00r|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��L?��jK���xY00r|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'   � ��L?��jK���xY0,q|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��L?��jK���OxY0,q|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��L?��iK���OxY0(p|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��L?��iK���OxY@(p|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A���iK���OxY@$o|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A���iK���OxY@ o|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A���hK���OxY@ n|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A���hK���OxY@m|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A��hK���OxY@m|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A��hK���OxY@l|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A�� hK���OxY@k|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A�� gK���OxY@j|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A_� gK��� xY@j|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A_� gK��� |Y@i|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A_�� gK��� |YPh|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A_�� fK��� |YPg|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A_���fK��� |YP f|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A_���fK����|Y_�e|( /��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A���eK�����Y_�d|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A��eK�����Y_�c|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A� dK�����Y_�b|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A� dK�����Y_�a|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A� cK�����Y_�a|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��@�� cK�����Y_�`|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��@��� b@����Y_�_|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��@���b@����Yo�^|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��@��~�a@����Yo�^|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��@��~�a@����Yo�]|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�~�`@����Yo�]|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�~�_@����Yo�\|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�}�_@�� �Yo�\|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�}�^@�� �Yo�\|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�|�^@�� �Yo�[|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�{�]@�� �Yo�[|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��{�]@�� �Yo�[|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��z�\@���Yo�[|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��z� \@���Yo�Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��y�$\@���Yo�Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��x�([@���Yo�Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��x�,[@���Yo�Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��w�0Z@���Yo�Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��w�4Z@���Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��v�<Y@���Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��v�@Y@���Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��u�DY@���Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��u�HX@���Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��t	HX@���Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��t	HX@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��s	LX@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��s	LX@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��r	LW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��r	/LW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��q	/PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��q	/PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��p	/PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��p	/PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��o�PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��o�PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��o�PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��n�PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��n�PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��m�PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��m�PW@����Y��Z|( +��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��m�PW@����Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��l�PW@����Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��l�PW@����Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�PW@����Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�PW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�PW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�PW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�PW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�PW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�PW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TW@����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK�����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK�����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK����YO�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK����Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK����Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK����Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�k�TWK����Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�k�TWK���O�Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�k�TWK���O�Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�k�TWK���O�Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�k�TWK���O�Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�k�TWK���O�Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��CO�k�TWK���O�Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y�Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TWK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TVK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TVK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TVK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��K��k�TVK���O�Y��Z|( '��@ A�����3� T0 k� �����Y"t'!"t1'   ��'    � ��A���ǒ@�_�(:�C<H	���T@ D�,8��Z3� T0 k� ���#�P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�D<H	���T@ D�,8��Z3� T0 k� ���#�P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�D<H	���T@ D�,9��Z3� T0 k� ���#�P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�D<H	���T@ D�,:��Z3� T0 k� ���#�P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�E<H	\��T@ D�,;��Z3� T0 k� ���#�P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�E<H	\��T@ Em,<��Z3� T0 k� ���#�P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�F<H	\�,�U@ Em(=��Z3� T0 k� ���#�P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�F<H	\�,�U@ Em(>��Z3� T0 k� ���#�P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�F<H	\�,�U@ Em(?��Z3� T0 k� ���#�P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�G<H	\�,�V@ Em$@��Z3� T0 k� ���$P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�G<H	\�,�V@ Em$A��Z3� T0 k� ���$P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�H<H	\�,�W@ Em$BL�Z3� T0 k� ���$P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�H<H	\�,�W@ Em$BL�Z3� T0 k� ���$P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�H<H	\�,�W@ D=$DL�Z3� T0 k� ���$P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�I<H	l�,�X@ D= EL�Z3� T0 k� ���#;P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�I<H	l�,�X@ D= FL�Z3� T0 k� ���#;P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�J<H	l�,�X@ D= G|�Z3� T0 k� ���#;P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�J<H	l�,�Y@ D=H|�Z3� T0 k� ���#;P Y"t'!"t1'  ��   � )�8A���ǒ@�_�(:�J<H	l�,�Y@ I�I|�Z3� T0 k� ���#;P Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	l�,�Y@ I�J|�Z3� T0 k� ���#[P Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	l�,�Z@ I�K|�Z3� T0 k� ���#[P Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	l�,�Z@ I�K|�Z3� T0 k� ���#[P Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	l�,�Z@ I�L|�[3� T0 k� ���#[P Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	\�,�[@ I�M|�[3� T0 k� ���#[P Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	\�,�[@ I�N|�[3� T0 k� ���#kP Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	\�,�[@ I�N|�[3� T0 k� ���#kP Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	\�,�[@ I�N��[3� T0 k� ���#kP Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	\�,�\@ I�N��\3� T0 k� ���#kP Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	\�,�\@ EmO��\3� T0 k� ���#kP Y"t'!"t1'  ��   � )�8A���ǒ@�c�(:�K<H	\�,�]@ EmO��\3� T0 k� ���#{P Y"t'!"t1'  ��   � )�8A�����2@� O8# o;�| P< �(2@ A�+���#3� T0 k� �  � Y"t'!"t1'   ��/   �   2A�����2@� O8# o;�!� P< �(2@ A�+���#"s� T0 k� �  � Y"t'!"t1'   /�/   �   3A�����2@� O8# o;�!� P< �(2@ A�+���#"s� T0 k� ��Y"t'!"t1'  ��/   �   4A�����2@� O8# o;�!� P< �(2@ A�+���#"s� T0 k� ��Y"t'!"t1'  ��/   �   5A�����2@� O8# o;�!� P< �(2@ B@+�P�#"s� T0 k� ��Y"t'!"t1'  ��/   �   6A�����2@� O8# o;�!� P< �(2@ B@+�P�#"s� T0 k� ��Y"t'!"t1'  ��/   �   7A�����1@� O8# o;�!�  P< �(2@ B@/�P�#"s� T0 k� �	�	Y"t'!"t1'  ��/   �   8A�����1@� O8# o;�!�  P< �(2@ B@/�P�#"s� T0 k� �
�
Y"t'!"t1'  ��/   �   9@����1@�  8#O;�!�$ P< �(1@ B@/�P�#"s� T0 k� �� Y"t'!"t1'  ��/   �   :@����1@�  8#O;�|$ P< �(1@ D�/���#3� T0 k� �� Y"t'!"t1'  ��/   �   ;@����1@�  8#O;�|$ P< �(1@ D�/���#3� T0 k� � �$Y"t'!"t1'  ��/   �   <@����0@�  8#O;�|$ P< �(0@ D�3���#3� T0 k� � �$Y"t'!"t1'  ��/   �   =@����0@�  8#O;�|( P< �(0@ D�3���#3� T0 k� �$�(Y"t'!"t1'  ��/   �   >@o����0@�  o8#O;�|( P< �(/@ D�3���#3� T0 k� �(�,Y"t'!"t1'  ��/   �  >@o����/@�  o8#O;�|( P< �(/@ D�7���#3� T0 k� �(�,Y"t'!"t1'  ��'   �  >@o���/@�  o8#O;�|( P< �(.@ D�7��#3� T0 k� �$�(Y"t'!"t1'  ��'   �  >@o���.@�  o8#�;�|( P< �(-@ F 7��#3� T0 k� � �$Y"t'!"t1'  ��'   �  >@o���.@�  o8#�;�|( P< �(-@ F ;��#3� T0 k� �� Y"t'!"t1'  ��'   �  >CO���.@� 
O8#�;�|( P< �,,@ F ?��#3� T0 k� �� Y"t'!"t1'  ��'   �  >CO���-@� 
O8#�;�|( P< �,,@ F ?��#3� T0 k� � �$Y"t'!"t1'  ��'   �  >CO���,@� 
O8#�;�!�( P< �,+@ F C��#"�� T0 k� � �$Y"t'!"t1'  ��'   �  >CO��o�,@� 
O8#�;�!�( �< �,+@ F C��""�� T0 k� � �$Y"t'!"t1'  ��'   �  >CO��o�+@� 
O8#�;�!�( �< �,*@ E�G��""�� T0 k� � �$Y"t'!"t1'  ��'   �  >CO��o�*@� 
4#�;�!�( �< �,*@ E�K��""�� T0 k� � �$Y"t'!"t1'  ��'   �  >CO��o�)@� 
4#�;�!�( �< �0)@ E�K��!"�� T0 k� � �$Y"t'!"t1'  ��'   �  >CO��o�(@� 
4#�7�!�( �< �0)@ E�O��!"�� T0 k� �$�(Y"t'!"t1'  ��'   �  =CO��o�'@� 
0#�7�!�( �< �0(@ E�S��!"�� T0 k� �$�(Y"t'!"t1'  ��'   �  <CO��o�&@� 
0#�7�!�( �< �0(@ B�W�� "�� T0 k� �$�(Y"t'!"t1'  ��'   �  ;E/��_�%@� 
,#�3�!�( �< �0'@ B�[� � "�� T0 k� �$�(Y"t'!"t1'  ��'   �  :E/��_�$@� 
,#�3�!�( �< �0'@ B�_� �"�� T0 k� �$�(Y"t'!"t1'  ��'   �  9E/��_�$@� 
(#�3�!�( �< �0&@ B�c� �"�� T0 k� �$�(Y"t'!"t1'  ��'   �  8E/��_�#@� 
(#�/�|( �< �4&@ B�g� �3� T0 k� �$�(Y"t'!"t1'  ��'   �  7E/��_�"@� 
/$#�/�|( �?��4%@ E�k� �3� T0 k� �(�,Y"t'!"t1'  ��'   �  6E/����!@� 
/ #�+�|( �?��4%@ E�o� �3� T0 k� �(�,Y"t'!"t1'  ��'   �  5E/���� @� 
/#o+�|( �?��4$@ E�s���3� T0 k� �(�,Y"t'!"t1'   ��'   �  4E/����@� 
/#o'�|( �?��4#@ E����3� T0 k� �(�,Y"t'!"t1'   .�'   �  3E/����@� 
/#o#�|( �?��4#@ E�����3� T0 k� �(�,Y"t'!"t1'   ��'   �  2B����@� 
/#o#�|( �?��8#@ DЇ���3� T0 k� �(�,Y"t'!"t1'   ��'   �  1B����@� 
/#o#�|( �?��8"@ DЋ���3� T0 k� �(�,Y"t'!"t1'   ��'   �  0B����@� �#o#�|( �?��8"@ DГ���3� T0 k� �,�0Y"t'!"t1'   ��'   �  .B����@� �#o#�|( �?��8!@ DЗ���3� T0 k� �,�0Y"t'!"t1'   ��'   �  ,B����@� � #o�|( �?��8!@ DЛ���3� T0 k� �,�0Y"t'!"t1'   ��'   �  *B����@� ��#�|( �?��8!@ F ����3� T0 k� �,�0Y"t'!"t1'   ��'   �  (B����@� ��$�|( �?��8 @ F ����3� T0 k� �,�0Y"t'!"t1'  ��'   �  &B����@� ��$ |( �?��8 @ F ����3� T0 k� �,�0Y"t'!"t1'  ��'   �  $B����@� ��$|( �?��8 @ F ����3� T0 k� �,�0Y"t'!"t1'  ��'   �  "B����@� ��$|( �?��<@ F ����3� T0 k� �,�0Y"t'!"t1'   ��'   �  !B���@����%|( �?��<@ F ����3� T0 k� �0�4Y"t'!"t1'   ��'   �  B���@����&|( �?��<@ F �� �3� T0 k� �0�4Y"t'!"t1'   ��'   �  C ��@����&	|( �?��<@ E�� �3� T0 k� �0�4Y"t'!"t1'   ��'   �  C ��@����'�
|( �?��<@ E�� �3� T0 k� �0�4Y"t'!"t1'   ��'   �  C ��@����'�|( �?��<@ E�� �3� T0 k� �0�4Y"t'!"t1'   ��'   �  C ���@����'�|( �?��<@ E��� �3� T0 k� �0�4Y"t'!"t1'   ��'   �  C ���@����(�|( �?��<@ E���0�3� T0 k� �0�4Y"t'!"t1'   ��'   �  I0���@���(�|( `?��@@ E���0�3� T0 k� �0�4Y"t'!"t1'   ��'   �  I0#���@���)|( `;��@@ E���0�3� T0 k� �4�8Y"t'!"t1'   ��'   �  I0#���
@���)|( `;��@@ E���0�3� T0 k� �4�8Y"t'!"t1'   ��'   �  I0'���	@���*|( `;��@@ E���0�
3� T0 k� �4�8Y"t'!"t1'   ��'   �  I@+���@���*|( `7��@@ E���@�	3� T0 k� �4�8Y"t'!"t1'   ��'   �  	I@+���@����+�|( `7��@@ E���@�3� T0 k� �4�8Y"t'!"t1'   ��'   �  I@/���@����+�|( `3��@@ E���@�3� T0 k� �4�8Y"t'!"t1'   ��'   �                                                                                                                                                                              � � �  �  �  c A�  �J����  �      6 \��� ]�6E6D 
x �� k��  � �	   ���     k�_��    ��            ? Z��           �    ���   0
            V�   � �
     ��Ճ7     V� ��}=    �� Z             M  Z��          ��     ���   8	
�          ����  � �
      ���    �������                       Z��          �P�    ���   (	"           Y�=   $ $     ��UB     Y�=��UB                     	 Z��          �      ���   H
w          Z�   � �
	   .����     Z�����    ��     
          o	 Z��          0�    ���   (
           ��  ��     B�
�!      ���
�!                             Z���\              4  ���    0

 2            ��}�          V���+    ��}����+                      �� :         �`     ��@   @
"
          w�     	   j +�]     w� +�+                      �8         ��     ��H  8
         �X�      ~  v"    �X�  v"               ��    
	 � !         �        ��F    

'		          �뿬   	     � ��    �뿬 �¦       %             ?         	 �@     ��@   8
          ����        � n    ���� n�                     A F         
 P     ��@   X
	           � �       � �,      � �,                             ����              4  ��@    0 0                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         ����  ��        � (�Y    ���� (�'        "               x                j  �       �                         ��    ��        � )      ��   )           "                                                �                         �����������
�� +   � n ��� ( )                	 

   �  ,V  ���J       �d 0[� �� 0\  �$ \� �D  \� ��  \� Ф g@ �D ]`���X � �  ]@ (� `e� )D  f� H� _����< ����J ����X � �d u� 
�\ V� 
�\ V� 
�\ W  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� � }`���� � 
�| V  
�\ W� 
�\ W� 
�\ W����� � �d 0k� �� l  ��  l@ � �c@ �  d@ ބ �^@ ބ �e� �� h@ � �h` �$ i� ?� �m@ @� 0n@ A n� A$ n� �� �`� �� a� ?� �o� @� 0p� A q  A$ q@ $ `r@ � s    s ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������� ��   ������  
�fD
��L���"����D" � j  "  B   J jF�"     
�j 
 ���
��
��"     "�j��   * �
� �  �  
�      ��     � +      ��    ��     ���           ��     � +          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �'"      �� � �  ���        � �T ���        �        ��        �        ��        �    ��	    ��������        ��                         5�$ 8   ���                                     �               D���              + ���%��   ����          �    �DET ei Fedorov      0:00                                                                        4  3     �:cV �Rc^ � �B�H �B�@ �B�X �CK � C"C �K � �	K � �
K � �C.K � C6S � C7C � C8C � C9N � C:I �J�e �J�] � J�d �J�] �J�Z � � � � � � �cj � cr � Uc� � mc� � �"� � � "� �� � �
�	 � "� � � !"� � �""� � �#*� � �$"� � � %"� �&� � � 
�	 �(� � � 
�	 �*"� � � +"� �,� � � 
�	 �.� � � 
� �0� � � 
�X  *GoX  *KO �4bp � � 5b� ~ �6br ~ �  b� � �  b� � �9br ~ � :b� � y;bt � � <b� � � =b� ~ �>bv ~ �  b� ~                                                                                                                                                                                                                         �� P         �     @ 
        �     c P E e  ���� W               �������������������������������������� ���������	�
��������                                                                                          ��    �� �� ��������������������������������������������������������   �4, .� < Ԃ@��A��.������������������(���                                                                                                                                                                                                                                                                                                             @�����                                                                                                                                                                                                                                         5  
  +    ��  .�J      �  	                           ������������������������������������������������������                                                                                                                                        �  �                �        �    �            	     ���������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ����                                .     �  4�J                                     ������������������������������������������������������                                                                                                                                     �  ma              m      >  ��               	 
     � ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� ������������������            x                                                                                                                                                                                                                                                 
                                        	                    �             


             �  }�                                                 V                                        ��������  R�  + ����������������������������  O������������  Rt��������  + ����������������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" A C 6                                 � Ї� �\                                                                                                                                                                                                                                                                                       )n)n1n  �"E        c            m            k      k            k                                                                                                                                                                                                                                                                                                                                                                                                        > �  
>�  J�  '#�  :#�  Bm �̞��������̞�h�̞������ �V ���� ������          <        ����           �   & AG� �  �   
           ���                                                                                                                                                                                                                                                                                                                                      K N   �   
    !             !��                                                                                                                                                                                                                            Y   �� �� Ѱ��      �� <      ���������������������������������������������� ��� �������������� ������� ������������  ����� ��������� � �������������� ������ ������ �� �� ��������������������������������� �� ������ ���  ������� ����� ������������������������� ����� ���������������������� ��� ������� ������� ������� �������� �� ��� � ���������� ��� ������ �������������   ����������������� ����������������������������� ��� ��� �� ������ ����� ������ ����� � ��������� ��������� ������������������   �� X     $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    ;      >   � ��                       B     �   �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��     �� p���� ���� p���� �$��   `d  �@���6 ��  �@���6 �$ ^$ �s@  �@  �s@      p 
�� ��   p  �`  -���� ��  -���� �$ ^$   �    E 
j� ��  E 
j�    ���`  � ��� ��  � ��� �$ f �  ��f   �      �  ��   (�������2����  g���          f ^�          ��        (      ���~���2�������J��*���      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                                             �                       �e iV�U�i                    ��������eeY�                 fU��Ul���ř�Yf�    V  UY e�V ��P �Uf Ŗf f�U                �  �  �\  �� 
]�    �U�eVl�Vl�f�f��f�iUl�f��VfU��f�V�����Ɯfli��e�fl\�Vf\ilVlUV����eU������elfl��fl�Y��eUV��f�e��fU�UVf�feYfU�l�fUVf�f�feUfY�l�ffP \UU �eP fe� �V  i`  V   `    \l �l� ��� ��l ��V �lV \e 
V��ll��V�fVllUVYlefll��VlfleVeV�eU��e����f�l���flf��V��f�ff��\l\UleU��f�fVlU�l�f�fY�feleU`iU` U`  �leZfeV eU` ej  V                                �                �l   e                       Uf��leUUV�eUeY�� Y�            eeV�Ul�Plƕ �e` �`              P                                                                                             wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           " "! "   "      ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ "!  "" "  """ "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      " "! "   "      ""            """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                      � ��� ��� ܷz �rywgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �     �  �   �   ��  �  �   �   ��  �           �   �   �                                                  �               �  �  ��  �   �   �           �     �                              �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .      �����                     ���                                       �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        ��̙��� ��� �� ��  ��  ��  ��  �I �D 
T3 
TD 
UD 
UD TD  T�  ˸  �  
�  ,� "� �"" �"  ��̊��˰�̻ �̰ �˰ ̻  ��  ��  �D� DD� 3EJ 4EJ 4ED ET DT �@ �� ��  �� ̰ �+/ �"/�"/����      ""  ",  "�  �   �   �             �   ��  ˚����ɪ��̙�    �   ��  �� �� ��Ш���������"  "  �"  �"  ˰  �   �   �       �   ��   ��   �                  �   �   �   �   �   �   �   �                .                  �   �               �  ��� ݼ� w{� �װ vw��"" �"" ��" ��  ��� ��� ��  ��                                                                                                                                      �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �          
 "� ""� ""� "                       �                             ���                         �  ��                    �����                                       ���                              �   ���                            �   �                                                                                                         �  �  �  �� ݚ� }�Ȫ��˙������˼� ��  ��  ��  ��  ��  I� H� �E X�T X�S T�D �[ ˻  ˸  ��  
� �,"��"" "  �" �  ""� �� ˻ �˻ ��ݪ��کɨ��ˀ�̽ ��� ��  ̽  ̻  ̻  ˉ  ��  �D  DC  C3  #;  ;�� �� ��  �� "�  "  �"/ / ����� ��  �      �   �          �  �  "     "  "  "   "�  �  �   �   
                            �          �   �          �                    ��  ���� ��    �����                         �     �                                                                                                                                                                                                            �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                                  �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �        �  ��  ��  ww  ��  vv  w       "   "   "                                     �   �  �  �� �  �  �      �   �                  �  �˰ ��� �wp ���                                                                                                                                                                �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���                        �   �   �   "   "   "  !�    ��               �  �           �   �   �                     �  �� �� ��     �����                                        � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                         ��w �������̻��̊��̹��˼��˼�ۻ̻�"   ""  ""  "                   ̰ ˽ �� �w �& vv                   � � �  �    �  �  �   �   �  �  �  �   S�  T�"��""��"!�"" "" "!                �  ̻� ��� ��p }r`          �  �  �   �   �  �                         �   �                �  ̻� ��� ��p�}r` "�"�����   �� �          ����   �       �                                   �    ���  ��                    ��  ��  ���                   ���              �   ��  ���  � �    �                                                                                                                                       �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��                       �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������             ��  �   ��  �                    �     �                                       �   ���                            �   �                                                                                                                 �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �                               ��                     �   �                      �������  ���    �    �����                                  �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                                                                �   �  � �� � � ��  �� �� ɘ�������� ��� ��  �� �� ��  ��   ��  ��  �۰ �ۀ���(����D344U3U4USTC�̻�˻�̼ͻ�̻ت˻ڪ˻ڪ���������������������       ��   �      �   �   �   �   �        ��  ؍  ۲  ز  ;�  D�� D?� D?  �?  ��  ��  ��� ��� ��� ��� �Ȁ ��� ��� ��� ����������� �� �� ��� ��  �          ��  �  �    �   �   ��   �        ��                  ��          � � ����� ��                       �   �   �   �   �   �                                                                                                                                                �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""����������D��M��M""""����������""""�����ADMA����""""����DD�M�""""��������AD�DM�""""�����������A�A�""""������AD�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��M��M�������D����3333DDDD�DD�M�D�������3333DDDDD�������M�DM�D����3333DDDD��A�M�M���M�����3333DDDDMM������D��D����3333DDDDA�A�A�D��M�D�����3333DDDD�������������D������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ADA�LL��L�D����3333DDDD x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(XxLL����������D����3333DDDD w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww""""����������A������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(""""�������I�I������ �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((�""""�������I��D���I������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`�D�M�D���M������3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(MD�M�A�����MD�����3333DDDD � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(�""""�����AMAD������ � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(�""""������������������ � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5fFfFDfFFfFffdFffff3333DDDD u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�xDDFFDfFFfdFffff3333DDDD  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww""""wwwwwwwGGD'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+""""wwwwwwqwAqwAwA34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�""""wwwwqwqAwAqAqAq9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(�A�A�A�A��LD�����3333DDDD U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(��A�LDL�L�D�L�����3333DDDD =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=""""wwwwwwDGAD    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( """"wwwwqqDAAq x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx""""wwwwwwwGGwGGwGwGw w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9wwUQUUQUUQUUQUUUDUUUUU3333DDDD  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(DEQQUUDUTEUUUU3333DDDD �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((�""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq:cV �Rc^ � �B�H �B�@ �B�X �CK � C"C �K � �	K � �
K � �C.K � C6S � C7C � C8C � C9N � C:I �J�e �J�] � J�d �J�] �J�Z � � � � � � �cj � cr � Uc� � mc� � �"� � � "� �� � �
�	 � "� � � !"� � �""� � �#*� � �$"� � � %"� �&� � � 
�	 �(� � � 
�	 �*"� � � +"� �,� � � 
�	 �.� � � 
� �0� � � 
�X  *GoX  *KO �4bp � � 5b� ~ �6br ~ �  b� � �  b� � �9br ~ � :b� � y;bt � � <b� � � =b� ~ �>bv ~ �  b� ~3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������"�"��9�G�[�R��-�U�L�L�K�_� � � � � � � � � �.�/�=�����������������������������������������$��<�Z�K�\�K��B�`�K�X�S�G�T� � � � � � � �.�/�=����������������������������������������$���<�K�X�M�K�O��0�K�J�U�X�U�\� � � � � � �.�/�=�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������-�2�3� ���������������������������������������.�/�=�	�
�������������������� � � � � � �����������������������������������������%��������������������.�/�=� ��!������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            