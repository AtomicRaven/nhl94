GST@�                                                            \     �                                               J���      �  �             ���2���$�	 ʱ����������h�������        �g      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"     "�j��   * ��
  �                                                                              ����������������������������������      ��    a bbQ  111  c c  	     
                g  	                  hn ")1         ==:�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             ��  )          == �����������������������������������������������������������������������������                                D   4           @  &   �   �                                                                                 '     "h)n1  �)�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g> ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E 4 �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ���K�|S��b�XEY|, ��W ��@TATH0 ��t - T0 k� �@#T� cA��1p (uBR0`1 ��    �  ����K��S��b�\EY|, ��X ��@TATH0 ��t - T0 k� �@#T� cA��1p (uBR0`1 ��    �  ����K��S��b�`DY|, ��X ��@TATH0 ��t - T0 k� �@#T� cA��1p (uBR0`1 ��    �  ����K��R��b�dDY|, ��X ��@TATH0 ��t - T0 k� �@#T� cA��1p (uBR0`1 ��    �  ����K��R��b�hDY|, ��Y ��@TATH0 ��t - T0 k� �@#T� cA��1p (uBR0`1 ��    �  ����K��R��b�lDY|, ��Y ��@TATH0 ��t - T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����K��R��b�lCY|, ��Z ��@TATH0 ��t - T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����K��R��b�pCY|, ��Z ��@TATH0 ��t - T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����K��R��b�tCY|, ��[ ��@TATH0 ��t - T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����K��R��b�xCa�, ��\ ��@TATH0 ��t - T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����K��R��b�|Ba�, ��\ ��@TATL0 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��R��b�|Ba�, ��] ��@TATL0 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��R��bÀBa�, ��^ ��@XATL0 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��R��bÄBa�, ��_ ��@XATL0 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��R��bÈAa�, ��_ ��@XATL0 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��R �bÈAa�, ��` ��@XATL0 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��R �bÌAa�, ��a ��@XATL0 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��R �bÐAa�, ��b ��@XATL1 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��R �bÐ@a�, ��b ��@XATL1 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��R �bÔ@a�, ��c ��@XATL1 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��RC�bØ@Y|, ��d ��@XATL1 ��t - T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K��RC�bØ@Y|, ��d ��@XATL1 ��!� - T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��K��QC�bÜ?Y|, ��e ��@XATL1 ��!� - T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��K��QC�bà?Y|, ��f ��@XATL1 ��!� - T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��K��QC�bà?Y|, �f ��@XATL1 ��!� - T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B��QC�bä?Y|, �g ��@XATL1 ��!� - T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B��QC�bä?Y|, �h ��@XATL1 ��!� - T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B��QC�bè>Y|, �h ��@XATL1 ��!� . T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B��Q�bì>Y|, �i ��@XATL1 ��!� . T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B��Q�bì>Y|, �i ��@XATL1 ��!� . T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B��Q�bð>Y|, �j ��@XATL1 ��!� . T0 k� �@#԰ cA��1p (uBR0`1 ��    �  � ��B��Q�bð>Y|, �k ��@XATL1 ��!� . T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����B��Q�bô=Y|, �k ��@XATL1 ��t . T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����E�Q�bô=Y|, �l ��@XATL1 ��t . T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����E�Q�bø=Y|, #�l ��@XATL1 ��t . T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����E�Q�bü=Y|, #�m ��@XATL1 ��t . T0 k� �@#� cA��1p (uBR0`1 ��    �  ����E�Q�bü=Y|, #�m ��@XATL1 ��t . T0 k� �@#� cA��1p (uBR0`1 ��    �  ����E�Q�b��=Y|, #�n ��@XATL1 ��t . T0 k� �@#� cA��1p (uBR0`1 ��    �  ����E�Q�b��<Y|, #�n ��@XATL1 ��t . T0 k� �@#� cA��1p (uBR0`1 ��    �  ����E��Q�b��<Y|, #�o ��@XATL1 ��t . T0 k� �@#� cA��1p (uBR0`1 ��    �  ����E��QS�b��<Y|, #�p ��@XATL1 ��t . T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����E��QS�b��<Y|, #�p ��@XATL1 ��t . T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����E��QS�b��<Y|, #�q ��@XATL1 ��t . T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����E��QS�b��<Y|, #�q ��@XATL1 ��!� . T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����E��RS�b��<Y|, #�q ��@\ATL1 ��!� . T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����E��RS�b��;Y|, #�r ��@\ATL1 ��!� . T0 k� �@$� cA��1p (uBR0`1 ��    �  ����E��RS�b��;Y|, #�r ��@\ATL1 ��!� . T0 k� �@$� cA��1p (uBR0`1 ��    �  ����E� SS�b��;Y|, #�s ��@\ATL1 ��!� . T0 k� �@$� cA��1p (uBR0`1 ��    �  ����E�SS�b��;Y|, #�s ��@\ATL1 ��!� . T0 k� �@$� cA��1p (uBR0`1 ��    �  ����EtSS�b��;Y|, #�t ��@\ATL1 ��!� . T0 k� �@$� cA��1p (uBR0`1 ��    �  ����EtTc�b��;Y|, #�t ��@\ATL1 ��!� . T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����EtTc�b��;Y|, #�u ��@\ATL1 ��!� . T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����EtUc�b��;Y|, #�u ��@\ATL1 ��!� . T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����Et Vc�b��;Y|, #�u ��@\ATL1 ��!� . T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����Et$Vc�b��<Y|, #�v ��@\ATL1 ��t. T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����Et,Wc�b��<Y|, #�v ��@\ATL1 ��t. T0 k� �@#T� cA��1p (uBR0`1 ��    �  ����Et0Xc�b��<Y|, #�w ��@\ATL1 ��t- T0 k� �@#T� cA��1p (uBR0`1 ��    �  ����Et4Yc�b��<Y|, #�w ��@\ATL1 ��t- T0 k� �@#T� cA��1p (uBR0`1 ��    �  ����Et8Zc�b��<Y|, #�w ��@\ATL1 ��t- T0 k� �@#T� cA��1p (uBR0`1 ��    �  ����Et<[S�b��<Y|, #�x ��@\ATL1 ��t- T0 k� �@#T� cA��1p (uBR0`1 ��    �  ����EdD\S�b��=Y|, #�x ��@\ATL1 ��t- T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����EdH]S�b��=Y|, #�y ��@\ATL1 ��t- T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����EdL^S�b��=Y|, #�y ��@\ATL1 ��t- T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����EdL_S�b��=Y|, #�y ��@\ATL1 ��t- T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����EdP`S�b��>Y|, #�z ��@\ATL1 ��t- T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����EdTaS�b��>Y|, #�z ��@\ATL1 ��t- T0 k� �@#t� cA��1p (uBR0`1 ��    �  ����EdXcS�b��?Y|, #�z ��@\ATL1 ��t, T0 k� �@#t� cA��1p (uBR0`1 ��    �  ����EdXdS�b��?Y|, #�{ ��@\ATL1 ��t, T0 k� �@#t� cA��1p (uBR0`1 ��    �  ����Ed\e�b��@Y|, #�{ ��@\ATL1 ��t, T0 k� �@#t� cA��1p (uBR0`1 ��    �  ����Ed`f�b��@Y|, #�{ ��@\ATL1 ��t, T0 k� �@#t� cA��1p (uBR0`1 ��    �  ����ET`g�b��AY|, #�| ��@\ATL1 ��t, T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ETdi�b��BY|, #�| ��@\ATL1 ��t,  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ET`i�b��BY|, #�| ��@\ATL1 ��t,  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ET\i�b��CY|, #�} ��@\ATL1 ��t,  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ETXj�b��DY|, #�} ��@\ATL1 ��t,  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ETXj�b��DY|, �} ��@\ATL1 ��t,  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ETTk�b� EY|, �} ��@\ATL1 ��t,  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ETPk�b� FY|, �~ ��@\ATL1 ��t+  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����EDLk�b� GY|, �~ ��@\ATL1 ��t+  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����EDHl�b� GY|, �~ ��@\ATL1 ��t+  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����EDDl�b� HY|, � ��@\ATL1 ��t+  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ED@l�b� IY|, S�~ ��@\ATL1 ��t+  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ED<l�b� JY|, S�~ ��@\ATL1 ��t+  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����C�8l�b� KY|, S�~ ��@\ATL1 ��t+  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����C�4l�b��LY|, S�~ ��@\ATL1 ��t+  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����C�0l�b��LY|, S�} ��@\ATL1 ��t+  T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����C�(l�b��MY|, ��} ��@\ATL1 ��t+  T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����C�$l�b��NY|, ��} ��@\ATL1 ��t+  T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����C� l�b��OY|, ��} ��@\ATL1 ��t+  T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����C�l�b��PY|, ��| ��@\ATL1 ��t+  T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����C�k�b��QY|, ��| ��@\ATL1 ��t*  T0 k� �@#� cA��1p (uBR0`1 ��    �  ����C�k�b��RY|, ��{ ��@\ATL1 ��t*  T0 k� �@#� cA��1p (uBR0`1 ��    �  ����C�k�b��SY|, �{ ��@`ATL1 ��t*  T0 k� �@#� cA��1p (uBR0`1 ��    �  � ��Itk�b��TY|, �z ��@`ATL1 ��t*  T0 k� �@#� cA��1p (uBR0`1 ��    �  � ��It j�b��UY|, �y ��@`ATL1 ��t*  T0 k� �@#� cA��1p (uBR0`1 ��    �  � ��Is�j�b��WY|, �y ��@`ATL1 ��t*  T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Is�j�b��XY|, ��x ��@`ATL1 ��t*  T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Is�j�b��YY|, ��w ��@`ATL1 ��t*  T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Is�j�b��ZY|, ��v ��@`ATL1 ��t*  T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��I��j�b��ZY|, ��v ��@`ATL1 ��t*  T0 k� �@#�� cA��1p (uBR0`1 ��    �  �3��C���Bs�я�Y|, �O2G�D�AT�����>T0 k� ����cA��1p (uBR0`1  ��    �  �3��C���Bk�ы�Y|, ��R2C�D�AT�����AT0 k� ����cA��1p (uBR0`1  ��    �  �3��C���Bc���Y|, ��SBC�DۥAT�����CT0 k� ����cA��1p (uBR0`1  ��    �  �3��C���B_���Y|, ��UB?�DӥAT�����DT0 k� ����cA��1p (uBR0`1  ��    �  �3��C���B[���Y|, ��VB;�D˥AT�����FT0 k� ����cA��1p (uBR0`1  ��    �  �3��C���BS��{�Y|, ��XB7�D��AT���	��IT0 k� ����cA��1p (uBR0`1  ��    �  �3��D��2O��{�Y|, ��ZB3�D��AT���	��JT0 k� ����cA��1p (uBR0`1  ��    �  �3��D��2G��w�Y|, ��[B3�D��AT���	��LT0 k� ����cA��1p (uBR0`1  ��    �  �3��D��2C��s�Y|, ��\B/�D��AT���	�MT0 k� ����cA��1p (uBR0`1  ��    �  �3��D��2;��k�Y|, ��_B'�D��AT�� �
�PT0 k� ����cA��1p (uBR0`1  ��    �  �3��D��27��g�Y|, ��`B'�D��ATC�!�
�RT0 k� ����cA��1p (uBR0`1  ��    �  �3��D��23��c�Y|, �aR#�C��ATC�"�
�ST0 k� ����cA��1p (uBR0`1  ��    �  �3��D��2/��_�Y|, �bR�C�w�ATC�#�
�TT0 k� ����cA��1p (uBR0`1  ��    �  �3��D��2+��[�Y|, �cR�C�k�ATC�$�
�VT0 k� ����cA��1p (uBR0`1  ��    �  �3��D{�2#��PY|, �fR�C�[�ATC�'�
�XT0 k� ����cA��1p (uBR0`1  ��    �  � ���Ds�"��LY|, �gR�C�O�ATC�(�
�ZT0 k� ����cA��1p (uBR0`1  ��    �  � ���Dg�"��DY|, �hR�C�G�AT��)��[T0 k� ����cA��1p (uBR0`1  ��    �  � ���D_�"��@Y|, �iR�C�?�AT��+��\T0 k� ����cA��1p (uBR0`1  ��    �  � ���DO�"��8Y|, |kQ��C�+�AT��-��_T0 k� ����cA��1p (uBR0`1  ��    �  �3��DG����0Y|, tlQ��C�#�AT��/�x`T0 k� ����cA��1p (uBR0`1  ��    �  �3��D?����,Y|, pma��C��AT��0�taT0 k� ����cA��1p (uBR0`1  ��    �  �3��D7���$Y|, hna��C��AT��2�lbT0 k� ����cA��1p (uBR0`1  ��    �  �3��D+��� Y|, `oa��C��AT��3�hdT0 k� ����cA��1p (uBR0`1  ��    �  �3��D���Y|, Pqa��C��AT��6�\fT0 k� ����cA��1p (uBR0`1  ��    �  �3��C����	Y|, Hra��C��AT��8��XgT0 k� ����cA��1p (uBR0`1  ��    �  �3� C����	Y|, @sa��E�ߥAT��:��PhT0 k� ����cA��1p (uBR0`1  ��    �  �3� C����
Y|, <ta��E�ץAT��;��HiT0 k� ����cA��1p (uBR0`1  ��    �  �3� C����� �Y|, ,va��E�åAT��?��<lT0 k� ����cA��1p (uBR0`1  ��    �  �3�C������ �Y|, $wa��E⻥AT��@��8mT0 k� ����cA��1p (uBR0`1  ��    �  �3�C����� �Y|, x1��E⳦AT��B��0nT0 k� ����cA��1p (uBR0`1  ��    �  �3�C������Y|, y1��E⧦AT��D��,oT0 k� ����cA��1p (uBR0`1  ��    �  �3�C�����Y|, z1��E⟦AT��E��$pT0 k� ����cA��1p (uBR0`1  ��    �  �3�C����Y|, � {1��D2��AT��I��rT0 k� ����cA��1p (uBR0`1  ��    �  �3�C����Y|, ��|1��D2��AT��K��sT0 k� ����cA��1p (uBR0`1  ��    �  �3�C��"��Y|, ��}1��D2{�AT��L��tT0 k� ����cA��1p (uBR0`1  ��    �  �3�C��"��Y|, ��~1��D2s�AT��N��uT0 k� ����cA��1p (uBR0`1  ��    �  �3�C��"��Y|, ��1��D2g�AT��P�� uT0 k� ����cA��1p (uBR0`1  ��    �  �3�C��"��Y|, �Ѐ1�D2W�AT��S���wT0 k� ����cA��1p (uBR0`1  ��    �  �3�I���"��Y|, �Ȁ	�w�D2O�AT��U���xT0 k� ����cA��1p (uBR0`1  ��    �  �3�I�{�"���Y|, ���	�s�D2C�AT��W���xT0 k� ����cA��1p (uBR0`1  ��    �  � ��I�s�"���Y|, �	�k�D2;�AT��X���yT0 k� ����cA��1p (uBR0`1  ��    �  � ��I�k�"���Y|, �	�g�D23�AT��Z���yT0 k� ����cA��1p (uBR0`1  ��    �  � ��I�c�"��xY|, �	�c�D2'�AT��[�1�zT0 k� ����cA��1p (uBR0`1  ��    �  � ��I�[���pY|, �	�_�DB�AT��]�1�zT0 k� ����cA��1p (uBR0`1  ��    �  �3�I�O���`Y|, �~	�S�DB�AT��`�1�{T0 k� ����cA��1p (uBR0`1  ��    �  �3�I�G���XY|, ��~	�O�DB�AT��a�1�|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I�C�#��PY|, ��~	�K�DA��AT��c��|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I�;�'��LY|, �x~	�G�DA�AT��d��|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I�7�+��DY|, �p}	�G�DA�AT��f��|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I�/�/��<Y|, �h}	�C�DA�AT��g��|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I�+�3��0Y|, �`}	�?�DAױAT��h��|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I�#�;��$Y|, �P|	�7�DAǲAT�j��}T0 k� ����cA��1p (uBR0`1  ��    �  �3�I���C��Y|,  H|	�7�DQ��AT�k��|}T0 k� ����cA��1p (uBR0`1  ��    �  �3�I���G��Y|,  @|	�3�DQ��AT�l��t}T0 k� ����cA��1p (uBR0`1  ��    �  �3�I���K��Y|,  8|	�/�DQ��AT�m��l}T0 k� ����cA��1p (uBR0`1  ��    �  �3�I���S��Y|,  0|	�/�DQ��AT�n��d|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I���W���Y|,  ({	�+�DQ��AT�o��`|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I���_��Y|,  {	�+�EᓷAT�p��X|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I���c��Y|,  {	�'�EዷAT�q��P|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I���k��Y|,  {	�'�EჸAT�q��L|T0 k� ����cA��1p (uBR0`1  ��    �  �3�I����o��Y|,  {	�'�E�w�AT�r��D{T0 k� ����cA��1p (uBR0`1  $�    �  �3�I����w��Y|, �z	�'�E�o�AT�s��<{T0 k� 3���cA��1p (uBR0`1  ��    �  �3�I������o�Y|, �z	�#�E�_�AT��t��0zT0 k� 3���cA��1p (uBR0`1  ��    �  �3�I������o�Y|, �z	�#�E�W�AT��t��,yT0 k� 3���cA��1p (uBR0`1  ��    �  �3�I������o�Y|, �z	�#�E�O�AT��t��$yT0 k� 3���cA��1p (uBR0`1  ��    �  �3�I������o� Y|, �z	�#�E�G�AT��u�� xT0 k� ����cA��1p (uBR0`1  ��    �  �3�I������o� Y|, �z	��E�?�AT��u��wT0 k� ����cA��1p (uBR0`1  ��    �  �3�I������o�!Y|, o�z	��E�7�AT�|u ���wT0 k� ����cA��1p (uBR0`1  ��    �  �3�I�������"Y|, o�z	��E�/�AT�xu ���vT0 k� ����cA��1p (uBR0`1  ��    �  � ��I����� �"Y|, o�z	��E�'�AT�tu ���uT0 k� ����cA��1p (uBR0`1  ��    �  � ��I������#Y|, o�{	��E��AT�tu ��� tT0 k� ����cA��1p (uBR0`1  ��     �  � ��I������$Y|, o�{	��E��AT�pu ����sT0 k� ����cA��1p (uBR0`1  ��     �  � ��E������%Y|, �{��E��AT�lu ����rT0 k� ����cA��1p (uBR0`1  ��     �  � ��E������&Y|, �{��F�AT�hu ����qT0 k� ����cA��1p (uBR0`1  ��     �  � ��E������'Y|, �|��F�AT�du �� �pT0 k� ����cA��1p (uBR0`1  $�     �  � ��E������'a�, �|��F ��AT�du �� �oT0 k� 3���cA��1p (uBR0`1  ��    �  � ��E�����|(a�, �|��F ��AT�`t �� �nT0 k� 3���cA��1p (uBR0`1  ��    �  � ��E�� ��x)a�, �|A�F ��AT�\t �� �mT0 k� 3���cA��1p (uBR0`1  ��    �  � c�E�� �	�t*a�, ��|A�F ��AT�\t �� �lT0 k� 3���cA��1p (uBR0`1  ��    �  � c�E�� �
�p+a�, ��|A�F ��AT�Xs ����kT0 k� 3���cA��1p (uBR0`1  ��    �  � c�E����h-a�, ��|A�F ��AT�Ts ����jT0 k� ����cA��1p (uBR0`1  ��    �  � c�E��� �d.a�, ��{A�F ��AT�Pr ����hT0 k� ����cA��1p (uBR0`1  ��    �  � c�E���(�`/a�, �|{�#�F ��AT�Pr ����gT0 k� ����cA��1p (uBR0`1  ��    �  � �F ��<�T1a�, t{�#�F ��AT�Hq ����eT0 k� ����cA��1p (uBR0`1  $�    �  � �F ��D�P2a�, pz�#�F ��AT�Hp ����cT0 k� ����cA��1p (uBR0`1  ��    �  � �F ��L�L3Y|, lz�#�F ��AT�Do ����bT0 k� ����cA��1p (uBR0`1  ��    �  � �F ��X�D4Y|, hz�#�E���AT�Do ���aT0 k� ����cA��1p (uBR0`1  ��    �  � �F ��`�@5Y|, `z�#�E���AT�@n ���`T0 k� ����cA��1p (uBR0`1  ��    �  ��F ��h�<7Y|, \z #�E���AT�<m ���^T0 k� ����cA��1p (uBR0`1  ��    �  ��F �	p48Y|, �Xz #�E���AT�<l ���]T0 k� ����cA��1p (uBR0`1  ��"    �  ��E��	x09Y|, �Tz #�E���AT�8k ���[T0 k� ����cA��1p (uBR0`1  ��"    �  ��E��		�,:Y|, �Pz #�E���AT�8j �� �ZT0 k� ����cA��1p (uBR0`1  ��"    �  ��E��
	�$;Y|, �Hz #�E���AT�4j �� �YT0 k� ����cA��1p (uBR0`1  ��"    �  ��E��	� <Y|, �Dz #�B���AT�0i �� �WT0 k� ����cA��1p (uBR0`1  $�"    �  �#�E���=Y|, @z #�B���AT�0h �� �VT0 k� 3���cA��1p (uBR0`1  ��/    �  �#�E���?Y|, 8z #�B���AT�,f �� �TT0 k� 3���cA��1p (uBR0`1  ��/    �  �#�E���
Aa�, 0z #�B���AT�(d �� �QT0 k� 3���cA��1p (uBR0`1  ��/    �  �#�E���
 Ba�, (z a#�B���AT�(c �� �PT0 k� 3���cA��1p (uBR0`1  ��/    �  �#�E���
�Ca�, �$z a#�B���AT�$b ����NT0 k� ����cA��1p (uBR0`1  ��/    �  �#�E���
�Da�, � z a#�B���AT�$a ����MT0 k� ����cA��1p (uBR0`1  ��/    �  �#�E���
�Ea�, �z a#�B���AT� _ ����KT0 k� ����cA��1p (uBR0`1  ��/    �  �#�E��#���Ea�, �y a#�B���AT� ^ ����JT0 k� ��� cA��1p (uBR0`1  ��/    �  ��E��#���Fa�, �y a#�B���AT] ����HT0 k� ��� cA��1p (uBR0`1  $�/    �  ��E��#���Ga�, �y a#�B���AT\ ����GT0 k� 3�� cA��1p (uBR0`1  ��/    �  ��E��#���Ha�, �y a#�B���ATZ ����ET0 k� 4 �cA��1p (uBR0`1  ��/    �  �� E��#���Ia�, �x a#�B���ATY ����DT0 k� 4 �cA��1p (uBR0`1  ��/    �  �� E��#���IY|, x a#�B���AT W ����CT0 k� 4�cA��1p (uBR0`1  ��    �  � c� E��#���JY|,  x a#�B���AT V ����AT0 k� 4�cA��1p (uBR0`1  ��    �  � c� @`�3���JY|,  w a#�B�� AT U ����@T0 k� � �cA��1p (uBR0`1  ��     �  � c��@`�3���KY|, ~�w a#�B��AT S ����?T0 k� ��� cA��1p (uBR0`1  ��     �  � c��@`�3�޼KY|, ~�v a#�B��AT R ����>T0 k� ����cA��1p (uBR0`1  ��     �  � c��@`�3�޸LY|, �u a#�B��AT!P ����=T0 k� ����cA��1p (uBR0`1  ��     �  � ��@`�3�޴LY|, �u #�B��AT!O ����;T0 k� � 
�
cA��1p (uBR0`1  $�     �  � ��B��3�ްMY|, �t #�B��AT!�N ����:T0 k� 4	�	cA��1p (uBR0`1  ��    �  � ��B��3�ްMY|, �s #�B��AT!�L ���9T0 k� 4	�	cA��1p (uBR0`1  ��    �  � ��B��3� ެMY|, �s #�B��AT!�K ���8T0 k� 4�cA��1p (uBR0`1  ��    �  � ��B� 3� ިNY|, �r '�B��AT!�I ���7T0 k� 4�cA��1p (uBR0`1  ��    �  ���B�3� ޤNY|, �q�'�B��	AT"�H ���6T0 k� 4�cA��1p (uBR0`1  ��    �  ���B�3�!ޤNY|, ��p�'�B��
AT"�F ���5T0 k� ��cA��1p (uBR0`1  ��    �  ���B�3�!ޠNY|, ��p�+�B��
AT"�E ���4T0 k� ��cA��1p (uBR0`1  ��    �  ���B�3�"ޠNY|, ��o�+�B��AT"�C ���3T0 k� ��cA��1p (uBR0`1  ��    �  ���B�3�"�OY|, ��n�+�B��AT "�B ���3T0 k� ��cA��1p (uBR0`1  ��    �  �#��C 3�"�OY|, ��m�/�B��AT "�@ ���2T0 k� ��cA��1p (uBR0`1  ��    �  �#��C$3�#�OY|, �l�3�B��AT #�> ���1T0 k� ��cA��1p (uBR0`1  ��    �  �#��C,3�#�OY|, �k�3�B��AT #�= ����0T0 k� ��cA��1p (uBR0`1  ��    �  �#��C03�$�OY|, �j�7�B��AT #�; ����/T0 k� �@#4� cA��1p (uBR0`1  �    �  �#��E@3�$�OY|, �h�;�B� AT #� 8 ��� -T0 k� �@#4� cA��1p (uBR0`1 �    �  �#��ED3�%��OY|, ��g�?�B�AT #�$7 � �,T0 k� �@#4� cA��1p (uBR0`1��    �  ���EL3�%��NY|, ��f�C�B�AT $�$5 �  ,T0 k� �@#4� cA��1p (uBR0`1��    �  ���ET3�%��NY|, ��e C�B�AT $�$4 �  +T0 k� �@#D� cA��1p (uBR0`1��    �  ���E\3�&��NY|, ��d G�B�AT$$�(2 �  *T0 k� �@#D� cA��1p (uBR0`1��    �  ���E`3�&��NY|, ��c K�@AT$$�(1 �  )T0 k� �@#D� cA��1p (uBR0`1��    �  ���B�h3�&��NY|, ��b O�@ AT$$�(0 (T0 k� �@#D� cA��1p (uBR0`1��    �  � ��B�p3�'��NY|, ��a O�@$AT$$�,. (T0 k� �@#D� cA��1p (uBR0`1��    �  � ��B�x3�'��NY|, ��` S�@(AT$$ ,-  'T0 k� �@#T� cA��1p (uBR0`1��    �  � ��B��3�'��NY|, ��` S�@,AT$% 0, $&T0 k� �@#T� cA��1p (uBR0`1��    �  � ��B��3�(��NY|, ��_ W�@0AT$% 0* (%T0 k� �@#T� cA��1p (uBR0`1��    �  � ��B��3�(��NY|, � ^ [�@4AT$% 0) ,%T0 k� �@#T� cA��1p (uBR0`1��    �  � ��E�3�(��NY|, �] [�@8AT$% 4( 0$T0 k� �@#T� cA��1p (uBR0`1��    �  � ��E�3�)��NY|, �\ _�@<AT$% 4& 0$T0 k� �@#d� cA��1p (uBR0`1��    �  � ��E�3�)��NY|, �[ _�@@AT$% 4% 4$T0 k� �@#d� cA��1p (uBR0`1��    �  � ��E�3�)��NY|, �[ c�@DAT$% 8$ 8$T0 k� �@#d� cA��1p (uBR0`1��    �  � ��E�3�)��NY|, �Z g�@LAT(% 8#� <$T0 k� �@#d� cA��1p (uBR0`1��    �  � ��E�3�*��NY|, �Y g�@PAT(& 8"� @$T0 k� �@#d� cA��1p (uBR0`1��    �  � ��E�3�*��NY|, �X k�@TAT(& <!� D$T0 k� �@#t� cA��1p (uBR0`1��    �  � ��E��3�*��NY|, �W k�@XAT(& <� D$T0 k� �@#t� cA��1p (uBR0`1��    �  � ��E��3�*��NY|, �$W o�@\AT(& <� H#T0 k� �@#t� cA��1p (uBR0`1��    �  � ��E��3�+��NY|, �(V o�@`AT(& @� L#T0 k� �@#t� cA��1p (uBR0`1��    �  � ��E��3�+��NY|, �,U s�@dAT(& @� P#T0 k� �@#t� cA��1p (uBR0`1��    �  � ��E��3�+��MY|, �0U s�@hAT(& @� T#T0 k� �@#�� cA��1p (uBR0`1��    �  � ��D� 3�+��MY|, �4T w�@hAT(& D� T#T0 k� �@#�� cA��1p (uBR0`1��    �  � ��D�3�,��MY|, �<S w�@lAT(& D� X#T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��D�3�,��MY|, �@S {�@pAT(' D� \#T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��D�3�,��MY|, �HR {�@tAT(' D� `#T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��D�$3�,��MY|, �LQ �@xAT(' H� `#T0 k� �@#�� cA��1p (uBR0`1 /�    �  � ��D�,3�-��MY|, �TQ �@|AT(' H� d"T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��D�43�-��MY|, �XP ��@�AT,' H� h"T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��D�<3�-��MY|, �`O ��@�AT,' H� l"T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��D�D 3�-��MY|, �dO ��@�AT,' L� l"T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��LrL 3�.��MY|, �lN ��@�AT,' L� p"T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��LrX!3�.��MY|, �pM ��@�AT,' L� t"T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Lr`!3�.��MY|, �xM ��@�AT,' L� t"T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Lrh!3�.��MY|, πL ��@�AT,( P� x"T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Lrp"3�.��MY|, ߈L ��@�AT,( P� x"T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Lrt"3�/��MY|, ߌK ��@�AT,( P� |"T0 k� �@#İ cA��1p (uBR0`1 ��    �  � ��Lr|#3�/��MY|, ߔK ��@�AT,( P� �"T0 k� �@#İ cA��1p (uBR0`1 ��    �  � ��Lr�#3�/��MY|, ߜJ ��@�AT,( T� �!T0 k� �@#İ cA��1p (uBR0`1 ��    �  � ��Lr�#3�/��MY|, ߤJ ��@�AT,( T� �!T0 k� �@#İ cA��1p (uBR0`1 ��    �  � ��Lr�$3�/��MY|, ߬I ��@�AT,( T
� �!T0 k� �@#İ cA��1p (uBR0`1 ��    �  � ��Lr�$3�0� MY|, ߴI ��@�AT,( T	,$ �!T0 k� �@#� cA��1p (uBR0`1 ��    �  � ��Lr�%3�0�MY|, ߼H ��@�AT,( X,$ �!T0 k� �@#� cA��1p (uBR0`1 ��    �  � ��Lr�%3�0�MY|, ��H ��@�AT,( X,$ �!T0 k� �@#� cA��1p (uBR0`1 ��    �  � ��Lr�%3�0�MY|, ��G ��@�AT,( X,$ �!T0 k� �@#� cA��1p (uBR0`1 ��    �  � ��L��&3�0�MY|, ��G ��@�AT,( X,$ �!T0 k� �@#� cA��1p (uBR0`1 ��    �  � ��L��&3�0�MY|, ��F ��@�AT0( X,$ �!T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L��&3�1� MY|, ��F ��@�AT0) \,4 �!T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L��'3�1�$MY|, ��E ��@�AT0) \,4 �!T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L��'3�1�,MY|, ��E ��@�AT0) \,4 �!T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L��(3�1�4MY|, ��D ��@�AT0) \,4 �!T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L��(3�1�8MY|, �D ��@�AT0) \,4 � T0 k� �@$� cA��1p (uBR0`1 ��    �  � ��L��(3�1�@MY|, �C ��@�AT0) \,4 � T0 k� �@$� cA��1p (uBR0`1 ��    �  � ��L��)3�2�DMY|, �C ��@�AT0) `,D � T0 k� �@$� cA��1p (uBR0`1 ��    �  � ��L��)3�2�LMY|, �C ��@�AT0) ` ,D � T0 k� �@$� cA��1p (uBR0`1 ��    �  � ��L��)3�2�TMY|, �$B ��@�AT0) c�,D � T0 k� �@$� cA��1p (uBR0`1 ��    �  � ��L��)3�2�XLY|, �,B ��@�AT0) c�,D � T0 k� �@#4� cA��1p (uBR0`1 ��    �  � ��L� *3�2�`LY|, �4A ��@�AT0) c�,D � T0 k� �@#4� cA��1p (uBR0`1 ��    �  � ��L�*3�2�hLY|, �<A ��@�AT0) g�,D � T0 k� �@#4� cA��1p (uBR0`1 ��   �  � ��L�*3�3�lLY|, �DA ��@�AT0) g�,D � T0 k� �@#4� cA��1p (uBR0`1 ��    �  � ��L�+3�3�tLY|, �L@ ��@�AT0) g�,D � T0 k� �@#4� cA��1p (uBR0`1 ��    �  � ��L�+3�3�|LY|, �T@ ��@�AT0* g�,D � T0 k� �@#T� cA��1p (uBR0`1 ��    �  � ��L�+3�3��LY|, �\? ��@�AT0* g�,D � T0 k� �@#T� cA��1p (uBR0`1 ��    �  � ��L� +3�3��LY|, �d? ��@�AT0* g�,D � T0 k� �@#T� cA��1p (uBR0`1 ��    �  � ��L�$,3�3��LY|, �p? ��@�AT0* k�,T � T0 k� �@#T� cA��1p (uBR0`1 ��    �  � ��L�(,3�3��LY|, �x> ��@�AT0* k�,T � T0 k� �@#T� cA��1p (uBR0`1 ��    �  � ��L�,,3�3��LY|, ��> ��@�AT0* k�,T � T0 k� �@#d� cA��1p (uBR0`1 ��    �  � ��L�0-3�4��LY|, ��> ��@�AT4* k�,T � T0 k� �@#d� cA��1p (uBR0`1 ��    �  � ��L�8-3�4��LY|, ��= ��@�AT4* k�,T �T0 k� �@#d� cA��1p (uBR0`1 ��    �  � ��L�<-3�4��LY|, ��= ��@�AT4* k�,T �T0 k� �@#d� cA��1p (uBR0`1 ��    �  � ��L�@-3�4��LY|, ��= ��@�AT4* k�t �T0 k� �@#d� cA��1p (uBR0`1 ��    �  � ��L�D.3�4��LY|, ��< ��@�AT4* o�t �T0 k� �@#t� cA��1p (uBR0`1 ��    �  � ��L�H.3�4��LY|, ��< ��@�AT4* o�t �T0 k� �@#t� cA��1p (uBR0`1 ��    �  � ��L�L.3�4��LY|, ��< ��@�AT4* o�t �T0 k� �@#t� cA��1p (uBR0`1 ��    �  � ��L�P.3�4��LY|, ��; ��@�AT4* o�t �T0 k� �@#t� cA��1p (uBR0`1 ��    �  � ��L�T/3�5��LY|, ��; ��@�AT4+ o�t �T0 k� �@#t� cA��1p (uBR0`1 ��    �  � ��L�X/3�5��LY|, ��; ��@�AT4+ o�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L�\/4 5��LY|, ��; ��@�AT4+ o�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L�`/4 5��LY|, ��: î@�AT4+ o�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L�h04 5�LY|, ��: î@�AT4+ s�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L�l0D 5�LY|, ��9 î@�AT4+ s�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L�p0D 5� LY|, � 9 î@�AT4+ s�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L�t0D 5�(LY|, �9 Ǯ@�AT4+ s�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L�x0D 5�0LY|, �9 Ǯ@ AT4+ s�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��L�|1D 6�8LY|, �8 Ǯ@ AT4+ s�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Ls�1D 6�@LY|, � 8 Ǯ@ AT4+ s�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Ls�1D 6�HLY|, �(8 Ǯ@AT4+ w�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Ls�1D6�PLY|, �08 ˮ@AT8+ w�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Ls�1D6�XLY|, �47 ˮ@AT8+ w�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Ls�26�`LY|, �<7 ˮ@AT8, w�t �T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��Ls�26�hLY|, �D7 ˮ@AT8, w�t �T0 k� �@#İ cA��1p (uBR0`1 ��    �  � ��DӔ26�pLY|, �H7 ˮ@AT8, w�t �T0 k� �@#İ cA��1p (uBR0`1 ��   �  � ��DӘ26�xLY|, �P7 ˮ@AT8, w�t �T0 k� �@#İ cA��1p (uBR0`1 ��    �  � ��DӜ36ЀLY|, �X6 Ϯ@AT8, w�t �T0 k� �@#İ cA��1p (uBR0`1 ��    �  � ��DӠ37ЈLY|, �\6 Ϯ@AT8, w�t �T0 k� �@#İ cA��1p (uBR0`1 ��    �  � ��DӤ37��LY|, �d6 Ϯ@AT8, w�t  �T0 k� �@#԰ cA��1p (uBR0`1 ��    �  � ��E��47��LY|, �h6 Ϯ@AT8, {�t  �T0 k� �@#԰ cA��1p (uBR0`1 ��    �  � ��E��47��LY|, �p5 Ϯ@AT8, {�t  �T0 k� �@#԰ cA��1p (uBR0`1 ��    �  � ��E��5 d7��LY|, �t5 Ϯ@AT8, {�t  �T0 k� �@#԰ cA��1p (uBR0`1 ��    �  � ��E��5 d7��LY|, �|5 Ӯ@AT8, {�t! �T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����E��6 d7��LY|, ��5 Ӯ@AT8, {�t! �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����Es�7 d7��LY|, ��5 Ӯ@AT8, {�t! �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����Es�7 d7��LY|, ��4 Ӯ@AT8, {�t! �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����Es�8 �7��LY|, ��4 Ӯ@AT<, {�t! �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����Es�8 �7��LY|, ��4 Ӯ@AT<, {�t" �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����Es�9 �7��LY|, ��4 Ӯ@AT<, {�t" �T0 k� �@$� cA��1p (uBR0`1 ��   �  ����Es�9 �8��LY|, ��4 ׮@AT<, {�t" �T0 k� �@$� cA��1p (uBR0`1 ��    �  ����Es�: �8��LY|, ��4 ׮@AT<, �t" �T0 k� �@$� cA��1p (uBR0`1 ��    �  ����Es�;D8��LY|, ��3 ׮@AT<, �t" �T0 k� �@$� cA��1p (uBR0`1 ��    �  ����Es�<D9��LY|, ��3 ׮@AT<, �t# �T0 k� �@$� cA��1p (uBR0`1 ��    �  ����Es�=D9��LY|, ��3 ׮@ AT<, �t# �T0 k� �@#4� cA��1p (uBR0`1 ��    �  ����Es�?D:� LY|, ��3 ׮@ AT<, �t# �T0 k� �@#4� cA��1p (uBR0`1 ��    �  ����Es�@D:�LY|, ��3 ׮@ AT<, �t# �T0 k� �@#4� cA��1p (uBR0`1 ��    �  ����Es�A�;�LY|, ��3 ۮ@ AT<, �t# �T0 k� �@#4� cA��1p (uBR0`1 ��    �  ����Ec�B�<�LY|, ��2 ۮ@ AT<, �t# �T0 k� �@#4� cA��1p (uBR0`1 ��    �  ����Ec�C�<�LY|, ��2 ۮ@$AT<- �t$ �T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����Ec�E�=� LY|, ��2 ۮ@$AT<- �t$ �T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����Ec�F�>�$LY|, ��2 ۮ@$AT<- �t$ �T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����Ec�G�?�,LY|, ��2 ۮ@$AT<- �t$ �T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����Ec�I�@�0LY|, ��2 ۮ@(AT<- �t$ �T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����Ec�J�@�8LY|, ��1 ۮ@(AT<- ��t$ �T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����Ec�L�A�<LY|, ��1 ۮ@(AT<- ��t$ �T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����Ec�M�B�@LY|, ��1 ߮@(AT@- ��t% �T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����Ec�N�C�DLY|, ��1 ߮@(AT@- ��t% �T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����Ec�P�D�LLY|, ��1 ߮@,AT@- ��t% �T0 k� �@#d� cA��1p (uBR0`1 ��    �  ����Ec�Q�E�PLY|, ��1 ߮@,AT@- ��t% �T0 k� �@#t� cA��1p (uBR0`1 ��    �  ����Ec�S�G�TLY|, ��1 ߮@,AT@- ��t% �T0 k� �@#t� cA��1p (uBR0`1 ��    �  ����Ec�T�H�XLY|, � 1 ߮@,AT@- ��t% �T0 k� �@#t� cA��1p (uBR0`1 ��    �  ����ES�V�I�`LY|, �0 ߮@,AT@- ��t% �T0 k� �@#t� cA��1p (uBR0`1 ��    �  ����ES�W�J�dLY|, �0 ߮@0AT@- ��t& �T0 k� �@#t� cA��1p (uBR0`1 ��    �  ����ES�Y�K�hLY|, �0 ߮@0AT@- ��t& �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ES�Z�L�lLY|, �0 �@0AT@- ��t& �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ES�\�N�pLY|, �0 �@0AT@- ��t& �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ES�]�O�tLY|, �0 �@0AT@- ��t& �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ES�_�P�xLY|, �0 �@0AT@. ��t& �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ES�`�Q��LY|, � 0 �@4AT@. ��t& �T0 k� �@#�� cA��1p (uBR0`1 ��   �  ����ES�a�S��LY|, � / �@4AT@. ��t& �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ES�c�T��LY|, �$/ �@4AT@. ��t' �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����ES�d�V��LY|, �(/ �@4AT@. ��t' �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����EC�e�W��LY|, �,/ �@4AT@. ��t' �T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����EC�f� X��LY|, �0/ �@4AT@. ��t' �T0 k� �@#�� cA��1p (uBR0`1 ��   �  ����EC�g��Z��LY|, �0/ �@4AT@. ��t' �T0 k� �@#�� cA��1p (uBR0`1 ��   �  ����EC�h��[��LY|, �4/ �@8AT@. ��t'  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����EC�i��]��LY|, �8/ �@8AT@. ��t'  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����EC�j��^��LY|, �</ �@8AT@. ��t'  T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����EC�k��`��LY|, �@/ �@8AT@. ��t'  T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����EC�l��a��LY|, �D/ �@8AT@. ��t(  T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����EC�m��c��LY|, �H. �@8ATD. ��t(  T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����EC�m��d��LY|, �L. �@8ATD. ��t(  T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����EC�n��e��LY|, �P. �@<ATD. ��t(  T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����EC�o��g��LY|, �T. �@<ATD. ��t(  T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����EC�o��h��LY|, �X. �@<ATD. ��t( T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����E3�p��i��LY|, �`/ �@<ATD. ��t( T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����E3�p��j��LY|, �d/ �@<ATD. ��t( T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����E3�p��l��LY|, �h/ �@<ATD. ��t( T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����E3|qӼm��LY|, �l/ �@<ATD. ��t( T0 k� �@#� cA��1p (uBR0`1 ��    �  ����E3xq�n��LY|, �p/ �@@ATD. ��t) T0 k� �@#� cA��1p (uBR0`1 ��    �  ����E3tq�n��LY|, �x0 �@@ATD. ��t) T0 k� �@#� cA��1p (uBR0`1 ��   �  ����E3lq�o��LY|, �|0 �@@ATD/ ��t) T0 k� �@#� cA��1p (uBR0`1 ��    �  ����E3hq�p��LY|, �1 �@@ATD/ ��t) T0 k� �@#� cA��1p (uBR0`1 ��    �  ����E3dq�q��LY|, �1 �@@ATD/ ��t) T0 k� �@$� cA��1p (uBR0`1 ��    �  � ��E3\q�q��LY|, �1 �@@ATD/ ��t) T0 k� �@$� cA��1p (uBR0`1 ��    �  � ��E#Xq�r��LY|, �2 �@@ATD/ ��t ) T0 k� �@$� cA��1p (uBR0`1 ��    �  � ��E#Tp�s��LY|, �2 �@@ATD/ ��t ) T0 k� �@$� cA��1p (uBR0`1 ��    �  � ��E#Pp�s��LY|, �3 �@@ATD/ ��t ) T0 k� �@$� cA��1p (uBR0`1 ��    �  � ��E#Lp�t��LY|, �4 �@DATD/ ��t ) T0 k� �@#4� cA��1p (uBR0`1 ��    �  � ��E#Hp�t��LY|, �4 �@DATD/ ��t ) T0 k� �@#4� cA��1p (uBR0`1 ��    �  � ��E#Do�t��LY|, �5 �@DATD/ ��t ) T0 k� �@#4� cA��1p (uBR0`1 ��    �  � ��E#@o�u��LY|, �6 �@DATD/ ��t * T0 k� �@#4� cA��1p (uBR0`1 ��    �  � ��E#<n�xu� LY|, �6 �@DATD/ ��t * T0 k� �@#4� cA��1p (uBR0`1 ��    �  � ��E#<n�xu�LY|, �7 �@DATD/ ��t * T0 k� �@#D� cA��1p (uBR0`1 ��    �  � ��E#8m�tu�LY|, �8 �@DATD/ ��t * T0 k� �@#D� cA��1p (uBR0`1 ��    �  � ��E#4m�pu�LY|, �9 �@DATD/ ��t * T0 k� �@#D� cA��1p (uBR0`1 ��    �  � ��E4l�pu�LY|, �9 �@DATD/ ��t * T0 k� �@#D� cA��1p (uBR0`1 ��    �  � ��E0k�lu�LY|, �: �@DATD/ ��t * T0 k� �@#D� cA��1p (uBR0`1 ��    �  � ��E,k�hu� LY|, �; �@HATD/ ��t * T0 k� �@#T� cA��1p (uBR0`1 ��    �  � ��E,j�du�(LY|, �< �@HATD/ ��t * T0 k� �@#T� cA��1p (uBR0`1 ��    �  � ��E(j�`u�,LY|, �= �@HATD/ ��t * T0 k� �@#T� cA��1p (uBR0`1 ��   �  � ��B�(i\t�0LY|, �> �@HATD/ ��t * T0 k� �@#T� cA��1p (uBR0`1 ��    �  � ��B�(h\t�8LY|, �? �@HATD/ ��t * T0 k� �@#T� cA��1p (uBR0`1 ��    �  � ��B�(hXt�<LY|, @ �@HATD/ ��t * T0 k� �@#t� cA��1p (uBR0`1 ��    �  � ��B�$gTs�DLY|, A �@HATH/ ��t * T0 k� �@#t� cA��1p (uBR0`1 ��    �  � ��B�$gPs�HLY|, B �@HATH/ ��t * T0 k� �@#t� cA��1p (uBR0`1 ��    �  � ��B�$fPr�PLY|, C �@HATH/ ��t + T0 k� �@#t� cA��1p (uBR0`1 ��    �  � ��B�$fPr�XLY|, D �@HATH/ ��t + T0 k� �@#t� cA��1p (uBR0`1 ��    �  � ��B�$ePq�\LY|, $F �@HATH/ ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B�$d�Lq�dLY|, #,G �@HATH/ ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B�$d�Lq�hLY|, #4H �@LATH/ ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B�(c�Lq�pLY|, #8I �@LATH/ ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B�(b�Lp�xLY|, #@J �@LATH/ ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  � ��B�(a�LpҀLY|, #HK �@LATH/ ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����B�(a�Lo҄LY|, 	3LL �@LATH/ ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����B�,`�LoҌLY|, 	3TM �@LATH0 ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����B�,_�LnҔLY|, 	3\N �@LATH0 ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����B�,_LmҜLY|, 	3`O �@LATH0 ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�0^LmҠLY|, 	3dP �@LATH0 ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�0]LlҨLY|, 	ClQ �@LATH0 ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�4]LlҰLY|, 	CpQ �@LATH0 ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�4\LkҸLY|, 	CtR �@LATH0 ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�4[�Lk��LY|, 	CxS �@LATH0 ��t + T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�8[�Pj��LY|, 	C|S �@LATH0 ��t + T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����K�8Z�Pi��LY|, 	3�T �@LATH0 ��t , T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����K�8Y�Th��LY|, 	3�T �@PATH0 ��t , T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����K�<Y�Th��LY|, 	3�U �@PATH0 ��t , T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����K�<X�Xg��LY|, 	3�U �@PATH0 ��t , T0 k� �@#İ cA��1p (uBR0`1 ��    �  ����K�<W�\f��LY|, 	3�V �@PATH0 ��t , T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����K�<W�`f��LY|, 	C�V �@PATH0 ��t , T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����K�@V�`e��LY|, 	C�V �@PATH0 ��t , T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����K�@U�de�LY|, 	C�V �@PATH0 ��t , T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����K�@U�hd�LY|, 	C�W �@PATH0 ��t , T0 k� �@#԰ cA��1p (uBR0`1 ��    �  ����K�DU�lc�KY|, 	C�W �@PATH0 ��t , T0 k� �@#� cA��1p (uBR0`1 ��    �  ����K�HU�lc�KY|, 	3�W �@PATH0 ��t , T0 k� �@#� cA��1p (uBR0`1 ��    �  ����K�LU�lc�KY|, 	3�W �@PATH0 ��t , T0 k� �@#� cA��1p (uBR0`1 ��    �  ����K�PT�pc�JY|, 	3�W �@PATH0 ��t , T0 k� �@#� cA��1p (uBR0`1 ��    �  ����K�TT�tb� JY|, 	3�W �@PATH0 ��t , T0 k� �@#� cA��1p (uBR0`1 ��    �  ����K�XT�tb� JY|, 	3�W �@PATH0 ��t , T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�XT�tb�$IY|, 	C�W �@PATH0 ��t , T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�\S�xb�(Ia�, 	C�W �@PATH0 ��t , T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�`S�xb�,Ia�, 	C�W �@PATH0 ��t , T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�dS�|b�4Ha�, 	C�W �@TATH0 ��t , T0 k� �@#�� cA��1p (uBR0`1 ��    �  ����K�hS�|b�8Ha�, 	C�V �@TATH0 ��t , T0 k� �@#4� cA��1p (uBR0`1 ��    �  ����K�hS�|b�<Ha�, 	3�V ��@TATH0 ��t , T0 k� �@#4� cA��1p (uBR0`1 ��    �  ����K�lS�|b�@Ha�, 	3�V ��@TATH0 ��t , T0 k� �@#4� cA��1p (uBR0`1 ��    �  ����K�pS�|b�DGa�, 	3�V ��@TATH0 ��t , T0 k� �@#4� cA��1p (uBR0`1 ��    �  ����K�pS��b�DGa�, 	3�V ��@TATH0 ��t - T0 k� �@#4� cA��1p (uBR0`1 ��    �  ����K�tS��b�HGa�, 	3�V ��@TATH0 ��t - T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����K�tS��b�HFa�, ��W ��@TATH0 ��t - T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����K�tS��b�LFa�, ��W ��@TATH0 ��t - T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����K�xS��b�PFY|, ��W ��@TATH0 ��t - T0 k� �@#D� cA��1p (uBR0`1 ��    �  ����K�xS��b�TEY|, ��W ��@TATH0 ��t - T0 k� �@#D� cA��1p (uBR0`1 ��    �  �                                                                                                                                                                            � � �  �  �  c,�  �J����   �      � \��%� ]��� � �����        � �    ��� �           
            Z  Z �           �      ���   0	
	
           jJ�  � �	    � ��      jQ� ��U    	��              	 Z �         ��    ���@(	
           b�<           �\q     b�< �\q                        >	 Z �         p     ���   8�
          Z��   \ \	     ��X     ZW� �$x    	o�*   
            ' Z �          	��     ���  P



           � ��     .���      ����                               ���                d  ���    8	 1	             v�   H H	     B ��U     v�{ �q^    ����                & Z ��        ��     ���  (
	         ����          V ~ǽ    ���� ~�$       	                 	  K��           �P     ��@   8	(	          �         j �B     � �       1                 ����           �      ��@    
'           19?        ~+<     19?+<                        
     �          �`     ��J   8
	          ���l          � ���    ���l ���                          � �         	  �     ��@   X          *u� ��	     ��     *����    �+ �                 ��       
       �  ��@    0 0             �          � �]2     � �Z�       $                    J��           ��     ��@   @

               ��      �                                                                           �                               ��        ���          ��                                                                 �                          �  ��        �*     �*         "                   x                j  �   �    �                               ??       �,   �~    ,   ��    z�                                      . 4        �                          � � � �� � ~ � � ���,  
  	             
   �   / u  g��J       -� �h@ .� i@ .�  i` G$ d` �D _� G$ d` �D }� �� i` :d i� 
�< V� 
� V� 
�| W  $  ]  
�| W� 
� V� 
�| W  �d �t� �d u� 
�\ W� 
�� W� 
�\ W� �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ���� ����� � 
�| V ���� ����� � 
�| W ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���� �  ���  ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"     "�j��   * �
� �  �  
� ��    ��     � �  �   ��    ��     � �       1��  ��     �          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �      ��T ���        � � � ���        �        ��        �        ��        �      ��    ���	����        ��                         �$ (  ������                                     �                  ����             
  �
���%� �    ���               10 Hawerchukulet ny    0:01                                                                       1   0      �@cV �6c�&kj � �c� � �CI � CA �CB\ � CJT �	CKl �
B� � �C< �CD � C"L � C#T � 
�N �J�T �J�L � J�D �c� � c�
 �c�" � � � �	� � �	� � �� � �� �k~ � k� �� � �� � �"� � �  "� � �!"� � �"*� � �#"� � $"�# �%� �&
�  w'" �  (*H� � )*Kp � *)�� �  *O� �  *O� � -)�� �  *R� �  *O� � 0*x � 1*Qx �  *O� � 3*Qx �  *O� � 5*Qx �  *O� �  *O� �  *O� �  *O� �  *R� � ;*G� � <*Hp �  *R� � >*Kp �  *O�                                                                                                                                                                                                                         � P                     %� 
-     G P E V  ��                     �������������������������������������� ���������	�
��������                                                                                          ��   �� � ��������������������������������������������������������  �B�, &� ���                                                                                                                                                                                                                                                                                                                                                                    A@� @� A�                                                                                                                                                                                                                                              ��  L�J      ��                             �������������������������������������������������������                                                                                                                                        �    �4           �  x        �b     �             	 	 � ������������������� ����� �� ������������   ��������� ���������������� ����������������� ��� �������� �������������������������� ����� �����������������������������������������������������  ������������� ����� �����  ������                                     j            ��  4�J      :  	                           ������������������������������������������������������                                                                                                                                             �  �   +  b   �    V          ��               	 
     ������ �� ����������������� ����������������������������������������� �������� �� ���������� ���������������� �� ���� ������ ��������������������� ��� � ���� ����� ������ ������������������ �������������������������������� ������� ���                 �                                                                                                                                                                                                                                                                                                          
        �             


             �   }�   �    �#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" E B 5                                 � �� �\                                                                                                                                                                                                                                                                                  �      "h)n1  �)�             �3       d                  l      a      m                                                                                                                                                                                                                                                                                                                                                                                                                  ;#   >#  Iq� +# B#  Cm�  �̎���˖���������� ! � ��f�� ��  ������                       ���           �   &  AG� �   �                                                                                                                                                                                                                                                                                                                                                          [ X   �    N  ~�     "         !��                                                                                                                                                                                                                        Y��   �� �� �      �� 4  �� 
� ������������������� ����� �� ������������   ��������� ���������������� ����������������� ��� �������� �������������������������� ����� �����������������������������������������������������  ������������� ����� �����  ������������ �� ����������������� ����������������������������������������� �������� �� ���������� ���������������� �� ���� ������ ��������������������� ��� � ���� ����� ������ ������������������ �������������������������������� ������� ���             $������̼����˼̻���˻�̼������̼��̼��̻���Ƽ�ff��ff��ff��ff�fff�����fffffffffffffffffffffff�fff����f���ffl�ffflffffffffffffffff����˼̼�̻�̼��k˻�f˻�ff���f����˻�̼���̼̻���˻��˼���˼��˻���̼��˻��̼�˻���̼˼�̼�������fff�ffƶfff�fff�fff��f��fh��f��ffffffffffffffffffff���f���f����ffffffffffffffffffffffffffff̼��ffl�ffl�ffl�flk�ffl�ffl�ffl�ffl���˻̻����˻̻������̼����̼���˼��˼�̻���˻���������̼���̼����f���f���l���i���h���i���ʛ˶��˘�����������x����˪�ff��fk���j������������wy���w�fʇfl��jk��iʚ�ffk�ffk�flj��fl�vj��v���z��ˊ�{�˼��̻���������̼�����̻��������̻�˻�˻��˻�����̻������̼�˻˼̺������̺�������Ǚ�̪���ˉ������j���ȉw�������������������ˉ���lk���ˈw����y��������̙��ʘ�����y��ˈ�������x�˫��˻x˻��˻�����˻˻̻���˺�����˺��˼���˻����̻�̻���������̻���˼�˻��̼Ƨwww�˨��̷���ʈ��˙��̩�ˬ�����ww�����������fll���ƙ��l���ƙ���������������Ƽ����������������������������������������˪w�fȇ�fiw�f��̻˻�����˻�˻�k��ʌ���w����wxwuw����xwlff�������������ffff�fff����x�������fʇ�ll����j|f�k{fffy�������˘��̈�����������������������ʩ��f�������������������������f��|ly��j���h��f�ǖl\�fj��f�Ȧ�x���w�x����Xy�wx���x�wwffl��������                                         4     �     ���J���J    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       p���� ��   p���� �$ ^h  ��   p   	b��      
           �� �   6   
���(    �     �z � �N ^$a�       ��m        �c    �   ��������J � ��� �� �  � �N  � �  ��J  �      �     � �������2����   g���  �     f ^�  0     �� �      �       ��&H���2�������J������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  "  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��  DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰ wwwywww�www�www�www�www�www�www����������!��������������������a��������݈����������a������������(-�a������!�-���www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�www�������������������������������������!�����!�-����������!-�����������!������www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�www������m����������݈����������������a݈�����m����!�����������a�-������www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�wwwy-��������!�����������������������������������!��������                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         Dw D  4Dp 4Dw 4Dw 4DwpsGDDstDCsDD433G  DG   7                                    G   G   w   wp  wp  wp  wp  wwp p   ww                     	   2        �� 	�� 	�� ��� � � # 2 0 0                      y   2   s   ��wy�ypy�yp���p�w�t#w2#7 s7p pL��t���}���|���|���|���}�ww陙G   �p  �p  �p  �p  �p  �p  �p  J��t���{���z���z���z���{�ww陙G   �p  �p  �p  �p  �p  �p  �p  L��t���}���}����}��}��ww���G   �p  �p  �p  �p  �p  �p  w   J��t���{���{����{��{��ww���G   �p  �p  �p  �p  �p  �p  w    ��  ��  	�  ��  ��  �2  2#  0 �w�y� �	� � � � � � � � � " �wy��wy���	�	� �  	�  	�  	��w�y��y��w��w��w��w� " �  	�                           ""                             ff`                            330330330330330330330    ��p��p}}�p}}�pw��pwwp��p��pwp ww wwpwww  ww                                                                    ��p}�p}}�p}��pw�}pwww������     eW fWpffgw�p��p�p�w eVpvVpvvWpvgepwfvpwww�������w�y��y��w��w��w��w�"w���p��p y�p y�p��7��p�7 2#peVpfVpvvWpvvWpwgepwwp��p��p     w  wDpDDGG�G���p vdp         eg Uf ffpO�p��pwN�p         �� �� ��pO�p��pwN�p  y�  r'  p                    wy��wy���y�y�r'x�py�  y�  y� �p  �w �w �p Gp 7p wwpwwwwwpwp  wp  wp  p  p  w  w  w wp wpwwp wp wp wpwwwwwwwwC3GtDDDtDDDtDDDtDDDtwwtt334DDG      w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                                                �����   �   �   �   ����                                     
�  

  
 � 
 
 
   
   
   
   
  ��                  ��   
   
   
   
   
   
 
 
 � 

  
�                 �   
    �   
    �   
    �   
   
   �  
   �  
   �  
   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "  "!    " ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "  "!    " ""            """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       "! "   "      ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �   ��  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� �   �".  .                            �   �    �   �       �   �   �                .          ܰ  ˻  ��  �w  �&  vv        +  "  "     �  �               �  � �                       � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                                        0             �  �  � 
�� ��r ˚w
���	������ ��� ��� ",  "�  ". 34 DC3 DD3 �DC ��  ��  
"   "  "  ""  "!    �                    �   �   �   w   b�  g�� z�� ����̹���˙�̼̰������������蜚��L��>\���" ""  ""  �+ "	��"�������.�"��"! "  ��           �   ��  �   �    �  ��   �"" �"  �                        .   .   �                                 ��"� �"� ����            ���.�                         ��   �  ��  �  �  �         � ".��".��/����  �                                                                                                                                       �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���                         �  ��� ݼ� w��                                      "   "   "                                            �  "� "     �  �   �   �            "   "   "�  �                            �   ���                            �   "                                                                                                                           ̙ �ɪ���˭�̻� �� �   ""  ""  .         �� ̻ �� ��w �rb �wg���z�����ٙ�����ˍ�ݙ8����DD��3D��33L�3� �3+ ��" �" ""  ".  �  �   �                        �T  �U  �D  +�� ��� 
�  �"" �"" ��"/��� ��� �  ��               �   �   �   �   �   �   �@      �    �  �   �""��""����                "   "   "       �         �        �   �     �       �       "       .      �                    �"  �""� "�                                                                                                                                                                                                                 �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �                                                                                                                                                                                                                                                                                                    ̰ �� ̻ {��'��vz� w��  ��  ��  ̘  	�  
� "��,̻�"�� "#3  34  D  
�  �  " "" """ ! ��  ��                               ˹� �ɩ ��� �͋ ��� ��� ��̀��Ȑ���лܹнȝ0ݙ�@43�PCD�@@E�@ E�@ U�� H�  K�  �   ��    �� "�" ���                             "   "   .  ��                �   �   �   "   "   "  !�    ��                                 �   �                      �".��".  ���    �                    ".  ".  ���                                                                                                                                                                                                   �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �             "� /���  �       �   �   �                       "/ "�  �                                         �   �                      �".��".  ���    �                    ".  ".  ���                                                                                                                                                                                                   �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �"  "�  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �                    ".  ".  ���                                                                                                                                                                                                  	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��                        �          �   � � /  �"" �"  �                       �   �                      �".��".  ���    �        � ��                    ���� �                                                                                                                                                                                         �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �    �   �  .�  ."  �               �                         ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �                    ".  ".  ��� ���                                                                                                                                                                                                   �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �   �                                        �   �"           �    �� ��  �� �� ��� �           �   � �                   �         �  "� "  �  ��                                                                                                                                        �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �               �   �   P   T   U   T   S   C   3   30  30  ;�  ��  ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �                                                                                                                                                                                                                                           2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ D�D D@  �D�JJN�J��J��J��J��JJD�N�                    �   �       
    �  ��	���������                                                                                                                                                                                                                                                                                                                                                                                                                                                                               "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=""""��������AA�A    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ADA�LL��L�D����3333DDDD + , -   . / 0 1  	 2         3       4 (((((((2	10/(.(-(,(+LL����������D����3333DDDD 5 6   7   8 9 1 :   $ % ) ! " #   ; ) ! " # $ % ) (#("(!()(%($ :198(((7(6(5""""����������A������    <     = 8 0 1 > ? @ A B C D E F G H BC D I J KFE(DC(B(A(@?>108(=((( (<""""�������I�I������ L  . M + , N    O P Q R S S S T S S S T S ST S S ST S S ST S S SRQPO(( (N(,(+(M(.L""""�������I��D���I�������  7  N 5 U V W X Y S Z [ \ ] ^ _ ^ ^ ^ _ ^ ^_ ^ ^ ^_ ^ ^ ^_ ^]\[Z SY(X(W(V(U(5(N((7�D�M�D���M������3333DDDD  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`D�M�A�����MD�����3333DDDD 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
""""�����AMAD������ w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw""""������������������ w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xwwfFfFDfFFfFffdFffff3333DDDD + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+DDFFDfFFfdFffff3333DDDD � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(�""""wwwwwwwGGD � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(�""""wwwwwwqwAqwAwA �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(�""""wwwwqwqAwAqAqAq = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=A�A�A�A��LD�����3333DDDD    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( �A�LDL�L�D�L�����3333DDDD x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx""""wwwwwwDGAD w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww""""wwwwqqDAAq  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(""""wwwwwwwGGwGGwGwGw �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((�UQUUQUUQUUQUUUDUUUUU3333DDDD ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`DEQQUUDUTEUUUU3333DDDD M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M""""������������������������ � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(�""""�������DAADAI � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(��A�AM�M�DM��M334CDDDD 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5DD����M��DM�����3333DDDD x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x""""wwwwwwDGqGq w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwwGwwDGwwwwwwww + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+ADAH�DJ�H�H�����3333DDDD � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(��H��J�AD�DH�D����3333DDDD � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(�""""�������DD����� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq@cV �6c�&kj � �c� � �CI � CA �CB\ � CJT �	CKl �
B� � �C< �CD � C"L � C#T � 
�N �J�T �J�L � J�D �c� � c�
 �c�" � � � �	� � �	� � �� � �� �k~ � k� �� � �� � �"� � �  "� � �!"� � �"*� � �#"� � $"�# �%� �&
�  w'" �  (*H� � )*Kp � *)�� �  *O� �  *O� � -)�� �  *R� �  *O� � 0*x � 1*Qx �  *O� � 3*Qx �  *O� � 5*Qx �  *O� �  *O� �  *O� �  *O� �  *R� � ;*G� � <*Hp �  *R� � >*Kp �  *O�3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������������������������������� � � �m�n�|�}�c�d�v�w��� � � � � ������������������������������������������������� � � ������������������ � � � � ����������������������������������������������������2�G�]�K�X�I�N�[�Q��a��b� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%� �������������������-�2�3� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������,�>�0� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            