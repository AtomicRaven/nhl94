GST@�                                                            \     �                                                ��g      �  d   P         ����e J���J�������̸����������        6i     #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     "�j  " ���
��
�"    B�jl �   B ��
  ��                                                                              ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������=  0b  4  11                                         �  �  �  �                    
*          = �����������������������������������������������������������������������������                                �5  5       5�   @  #   �   �                                                                                '   $    )n)n1n  
*    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    �tm�O�D���IX�S�|,�G�I�M�L
�_����`qT0 k� ������(%2't �d1Q1   ��*    �  ��|l�W�D���IX�[�|,�K�I�M�T
�_����hpT0 k� ������(%2't �d1Q1   ��*    �  �	�l�g�D���I/\�k�|,�W�I#�M�`�_����xpT0 k� ������(%2't �d1Q1   ��*    �  �	�l�k�D��I/`�s�|,�[�I#�M�dғ�_���ЀoT0 k� ������(%2't �d1Q1   ��*    �  �	�l�s�D��I/`p{�|,�c�I#�M�lғ�_���ЈoT0 k� ������(%2't �d1Q1   ��*    �  �	�l�{�D��I/dp��|,�g�I#�M�pҗ�_���АnT0 k� ������(%2't �d1Q1   ��*    �  �	#�l���D�+�Idp��|,�o�I�M�|қ�_���РnT0 k� ������(%2't �d1Q1   ��*    �  �	#�lC��D�3�Ihp��|,�s�I�M��қ�_���ШmT0 k� ������(%2't �d1Q1   ��*    �  �	#�lC��D�?�Ihp��|,�w�I�M��қ�_����mT0 k� ������(%2't �d1Q1   ��*    �  �	#�lC��D�O�Ilp��|,�{�I�M��ҟ�_�����lT0 k� ������(%2't �d1Q1   ��*    �  �	�lC��D�W�B�lp��|,��I#�MØҟ�_�����kT0 k� ������(%2't �d1Q1   ��*    �  �	�l���D�c�B�pp��|,рI#�MÜ��_�����kT0 k� ������(%2't �d1Q1   ��*    �  �	�l���D�s�B�pp��|,фI#�Mä��_�����jT0 k� �� �� (%2't �d1Q1   ��*    �  �	�l���D�{�B�tp��|,фI#�Mè��_�����iT0 k� ����(%2't �d1Q1   ��*    �  �	#�l�ǯDă�B�x`��|,шI�Mì��_�����iT0 k� ����(%2't �d1Q1   ��*    �  �	#�l�˰Dă�B�x`��|,ш
I�Mðқ�_�����hT0 k� ����(%2't �d1Q1   ��*    �  �	#�l�׳D��B�|`��|,шI�Mø җ�_����gT0 k� �|��(%2't �d1Q1   ��*    �  �	#�l�ߵD�{�B��`��|,шI�Mü!җ�_����fT0 k� �t�x(%2't �d1Q1   ��*    �  ���l��D�{�E�`��|,ш@c�Mü#ғ�_����fT0 k� �l�p(%2't �d1Q1   ��*    �  �� k��D�w�E�a�|,�@c�M��&ҏ�_����$dT0 k� �h�l(%2't �d1Q1   ��*    �  ��k��BDs�E�a�|,�@c�M��'ҋ�_����,dT0 k� �d�h(%2't �d1Q1   ��*    �  ��k���BDs�E�a�|,�@c�M��)ҋ�_����4cT0 k� �` �d (%2't �d1Q1   ��*    �  ��j���BDo�E�a�|,�@��M��,҃�_����@bT0 k� �X�\(%2't �d1Q1   ��*    �  ��j��BDk�E�a�|,�@��M��-��_���HaT0 k� �T�X(%2't �d1Q1   ��*    �  ��i��BDk�E�a�|,�@��M��/�{�_���PaT0 k� �T�X(%2't �d1Q1   ��*    �  �� i��BDk�E�Q�|,�@��M��0�w�_���X`T0 k� �L�P(%2't �d1Q1   �*    �  �t,h��BDg�E�� Q'�|,�|@��M��3�o�_�{��h_T0 k� �8�<(%2't �d1Q1   ��/    �  �t0g��BDc�E�� Q+�|,�| A�M��4�k�[�w��p_T0 k� �,�0(%2't �d1Q1   ��/    �  �t4g��BDc�E���Q+�|,1x!A�M��6�g�[�o��x^T0 k� �$�((%2't �d1Q1   ��/    �  �t<f��BD_�E���Q/�|,1x"A�M��72c�[�k���]T0 k� �� (%2't �d1Q1  ��/    �  �t@e��BD_�E���Q3�|,1t#A�M��82_�[�g���]T0 k� ��(%2't �d1Q1  ��/    �  �tDd��BD_�E���Q3�|,1t$A�M��:2[�[�c���\T0 k� ��(%2't �d1Q1  ��/    �  �tHd�#�BD[�E���Q3�|,1p$AS�M��;2W�[�_���\T0 k� � �(%2't �d1Q1  ��/    �  �tTb�'�BDW�E���Q7�|,1l&AS�M��=2K�[�W���[T0 k� ��!��!(%2't �d1Q1  ��/    �  �tXa�'�BDW�E���A;�|,1h&AS�M��=2G�[�S���ZT0 k� ��$��$(%2't �d1Q1  ��/    �  �t\`�'�BDW�E���A;�|,1d'AS�N��>2C�[�O���ZT0 k� ��'��'(%2't �d1Q1  ��/    �  t`_�'�BDS�F��A;�|,1`'C�N��>2;�[�K�	�YT0 k� ��)��)(%2't �d1Q1  ��/    �  {dd^�'�BDS�F��A;�|,1\(C�O��>27�[�G�	�YT0 k� ��,��,(%2't �d1Q1   ��/    �  wdh]�+�BDS�F� A;�|,1\(C�O��?23�[�@ 	�YT0 k� ��/��/(%2't �d1Q1   ��/    �  sdl\�+�BDO�F� �;�|,�X(C�P��?2+�[�< 	�XT0 k� ��2��2(%2't �d1Q1   ��/    �  odp[�+�BDO�F  �;�|,�T(C�P��?B'�[�8 	�XT0 k� ��4��4(%2't �d1Q1   ��/    �  kdtY�'�BDO�F  �;�|,�P)C�Q�?B#�[�4��XT0 k� ��7��7(%2't �d1Q1   ��/    �  gdxW�'�BDK�F �;�|,�H)C�Q�@B�[�,��XT0 k� ��<��<(%2't �d1Q1   /�/    �  cd|V�'�BDK�F �;�|,�D)C�R��@B�[�(��WT0 k� ��?��?(%2't �d1Q1   ��/    �  _d|U�'�BDG�F $�;�|,�<)C�R��?R�[�$��WT0 k� �xB�|B(%2't �d1Q1   ��/    �  \d�S4#�BDG�D�,�;�|,�8)C�S��?R�[�$� WT0 k� �pD�tD(%2't �d1Q1   ��/    �  Yd�R4#�BDG�D�0�7�|,�4)C�S��?Q��[� �WT0 k� �hG�lG(%2't �d1Q1   ��/    �  Vd�Q4�BDC�D�8�7�|,�0)C�S��?Q��[��WT0 k� �\J�`J(%2't �d1Q1   ��/    �  ST�O4�BDC�D�@�7�|,�,(C�T��?Q��[��WT0 k� �TL�XL(%2't �d1Q1   ��/    �  PT�N4�BDC�D�D�3�|,�((C�T��>Q��[��WT0 k� �LO�PO(%2't �d1Q1   ��/    �   MT�M4�BD?�D�L�3�|,�$(C�T��>Q��[�� XT0 k� �@Q�DQ(%2't �d1Q1   ��/    � ! JT�L4�BD?�D�T�/�|,� 'C�|U��=Q��[��(XT0 k� �8T�<T(%2't �d1Q1   $�/    � " KT�J4�BD?�D�\�+�|,�'C�tU��=Q��[��0XT0 k� 28T�<T(%2't �d1Q1   ��/    � # L�I4�BD;�D�`�+�|,�&C�pU��<���[��4XT0 k� 2<T�@T(%2't �d1Q1   ��/    � $ M�H4�BD;�E�h	�'�|,�&C�lV��<���[��<XT0 k� 2<S�@S(%2't �d1Q1   ��/    � % N�GD�BD;�E�p	�#�|,�%DdV��;��[��@YT0 k� 2<S�@S(%2't �d1Q1   ��/    � & O�FD�BD;�E�x
�#�|,�$D`V��:��[� �HYT0 k� 2<S�@S(%2't �d1Q1   ��/    � ' P�ED�BD7�E�|��|,�$DXW��9��_���PZT0 k� �@S�DS(%2't �d1Q1   ��/    � ( Q�BD�BD7�E����|, "DLW��8��_���\[T0 k� �@R�DR(%2't �d1Q1   ��/    � ) R�AC��BD7�E����|, �!DDX��7��_���`[T0 k� �@R�DR(%2't �d1Q1   ��/    � * S�@C��BD3�E����|, � D@X��6��_���h\T0 k� �DR�HR(%2't �d1Q1   ��/    � * T�?C��BD3�E����|, �D8X��5��^r��l\T0 k� �DR�HR(%2't �d1Q1   ��/    � * U�>C��BD3�E����|, �D0Y��4�{�^r��p]T0 k� �DQ�HQ(%2't �d1Q1   ��/    � * V�=C��BD3�E����|, �D(Y��3�s�^r��x^T0 k� �DQ�HQ(%2't �d1Q1   ��/    � * W�<C��BD/�Ep����|, �D$Y��1�k�^r�	�|^T0 k� �HQ�LQ(%2't �d1Q1   ��/    � * X�|;S��BD/�Ep����|, �DZ��0�c�^r�	_T0 k� �HQ�LQ(%2't �d1Q1   ��/    � * Y�|:S��BD/�Ep����|,��DZ��/�[�^r�	`T0 k� �HQ�LQ(%2't �d1Q1   ��/    � * Z�x9S��BD/�Ep� �|,��DZ��.�S�^r�
aT0 k� �LP�PP(%2't �d1Q1   ��/    � * [�t7S��BD+�Ep� �|,� D�[��+�C�^��
bT0 k� �LP�PP(%2't �d1Q1   ��/    � * \�p6S��BD+�Ep� �|,�EB�[��*�;�^��cT0 k� �LP�PP(%2't �d1Q1   ��/    � * ]�l5S��BD+�Ep� ߳|,�EB�[��(�3�^� dT0 k� �PO�TO(%2't �d1Q1   ��/    � * ^�h5S��BD+�E`� ׳|,�EB�[��'�+�^� eT0 k� �PO�TO(%2't �d1Q1   ��/    � * _Td4S��BD'�E`� Ӳ|,�EB�[��%�'�^� fT0 k� �PO�TO(%2't �d1Q1   ��/    � * _T`3S��BD'�E`� ˲|,�EB�[��$��^�ҤgT0 k� �PO�TO(%2't �d1Q1   ��/    � * _T\2S��BD'�E`� Ǳ|,�EB�[��"��^�ҨhT0 k� �TO�XO(%2't �d1Q1   ��/    � * `TX1S��BD'�E`� ��|,�EB�[��!��^�ҨiT0 k� �TN�XN(%2't �d1Q1   ��/    � * `TT0S��BD'�EP� ��|,�EB�Z����^�ҨjT0 k� �TN�XN(%2't �d1Q1   ��/    � * `TP/S��BD#�EP���|,�E��Z����^�ҨkT0 k� �TN�XN(%2't �d1Q1   ��/    � * `TD.S��BD#�EP���|,� E°Y�����^�$ҬnT0 k� �XN�\N(%2't �d1Q1   ��/    � * aT@-��BD#�EP���|,�$E¬X�����^�,ҬoT0 k� �XM�\M(%2't �d1Q1   ��/    � * aT<,��BD#�EP���|,�$E¤W�����^�0ҬpT0 k� �XM�\M(%2't �d1Q1   ��/    � * aD8+��BD#�C����|,�(EW�����^�8ҬqT0 k� �\M�`M(%2't �d1Q1   �/    � * aD0+��BD�C�P��|, (EV����^�@ҬrT0 k� �dK�hK(%2't �d1Q1   �'    � * aD,*��BD�C�P��|, ,EU����^�DҬsT0 k� �dI�hI(%2't �d1Q1   ��'    � * aD )Sw�BD�C�Pw�|, 0EҀT����^�DҬuT0 k� �XJ�\J(%2't �d1Q1   ��'    � * aD)So�BD�L0�Ps�|, 0E�xS����^�DҬvT0 k� �PL�TL(%2't �d1Q1   ��'    � * aD(Sg�Lt�L0�@k�|, 4E�pR�
��^�HҬwT0 k� �HM�LM(%2't �d1Q1   ��'    � * aD(S_�Lt�L0�@c�|, 4E�hQ���^�HҬxT0 k� �@M�DM(%2't �d1Q1   ��'    � * aD'S[�Lt�L0�@[�|, 8E�`Q���^�LR�yT0 k� �8M�<M(%2't �d1Q1   ��'    � * aD'SS�Lt�L0�@S�|, 8AbXP���^�L
R�zT0 k� �$M�(M(%2't �d1Q1   ��'    � * a��'SK�Lt�L0�@O�|, 8AbPO���^�P	R�{T0 k� �L�L(%2't �d1Q1   ��'    � * a��'SC�Lt�L0�@G�|, <AbHO���^�TR�|T0 k� �K�K(%2't �d1Q1   ��'    � * a��&C;�Lt�L0�@?�|, <AbDN����Y�TR�}T0 k� ��K��K(%2't �d1Q1   ��'    � * a��&C3�Lt�L0�07�|, @Ab<M����Y�XR�~T0 k� ��J��J(%2't �d1Q1   ��'    � * a��&C+�Lt�L0�0/�|, @EB4M����Y�\R�T0 k� ��E��E(%2't �d1Q1   ��'    � * a��&C#�Lt�L0�0+�|, @EB,L�����Y�\R��T0 k� ��B��B(%2't �d1Q1   ��'    � * a��&C�Lt�L0�0#�|, DEB$K�����Y�`R��T0 k� ��?��?(%2't �d1Q1   ��'    � * a��&C�Lt�L0� 0�|, DEBK�����Y�`R�T0 k� ��<��<(%2't �d1Q1   ��'    � * a��%C�Lt�L0� 0�|, DEBJ����Y�dR�T0 k� ��:��:(%2't �d1Q1   ��'    � * a��%C�Lt�L@�!0�|, HEBI���{�Y�hR�T0 k� ��9��9(%2't �d1Q1   ��'    � * aӼ%B��L��L@�!0�|, HEBH���w�Y�hR�T0 k� ��7��7(%2't �d1Q1   ��'    � * aӴ%B��L��L@�"0�|, LEA�H���s�Y�lR�~T0 k� ��6��6(%2't �d1Q1   ��'    � * aӬ%B�L��L@�"?��|, LEA�G���o�Y�l R�~T0 k� ��5��5(%2't �d1Q1   ��'    � * a�%2�L��L@�"?�|, LEA�F���k�Y�p R�~T0 k� ��4��4(%2't �d1Q1   ��'    � * a�%2ߵL��L@�#/�|, PA�E���g�Y�s�R�~T0 k� ��3��3(%2't �d1Q1   ��'    � * a�$2׵L��L@�#/�|, PA�D���_�Y�w�R�~T0 k� ��2��2(%2't �d1Q1   ��'   � * a�$2ϵL��L@�#/�|, PA�D���[�Y�w�R�}T0 k� ��1��1(%2't �d1Q1   ��'    � * a�$2ǵL��L@�$/߱|, PA�C���W�Y�{�R�}T0 k� ��0��0(%2't �d1Q1   ��'    � * aC�$2��L��L@�$/۲|, TA�B���S�Y�{�R�}T0 k� ��/��/(%2't �d1Q1   ��'    � * aCx$2��L��L@�%/ӳ|, TA�A���O�Y��R�}T0 k� ��/��/(%2't �d1Q1   ��'    � * aCp$2��L��L@�%/ϳ|, TA�@���K�Y��R�}T0 k� �|.��.(%2't �d1Q1   ��'    � * aCh%B��L��L@�%�˴|, XA�?���G�Y���R�|T0 k� �x-�|-(%2't �d1Q1   ��'    � * aC`%B��L��L@�&�ǵ|, XA�>���C�Y���R�|T0 k� �p,�t,(%2't �d1Q1   ��'    � * aCX%B��L��L@�&�ö|, XA�=���C�Y���R�|T0 k� �h+�l+(%2't �d1Q1   ��'    � * aCP%B��L��L@�&���|, \Eј=���?�Y���R�|T0 k� �d/�h/(%2't �d1Q1   ��'   � * a�H&B��L��L@�'���|, \Eѐ<���;�Y���R�|T0 k� �`2�d2(%2't �d1Q1   ��'    � * a�@&B��L��L@�'���|, \Eь;���7�Y���R�{T0 k� �\4�`4(%2't �d1Q1   ��'    � * a�8&B��L��L@�'���|, \Eф:���3�Y���R�{T0 k� �X5�\5(%2't �d1Q1   ��'    � * a�0'B�L��L@�(���|, `E�|9���/�Y���R�{T0 k� �T6�X6(%2't �d1Q1   ��'    � * a�('Bw�L��L@�(���|, `E�t8���+�Y���R�{T0 k� �L6�P6(%2't �d1Q1   ��'    � * a� 'Bs�L��L@�(���|, `E�l8���'�Y���R�{T0 k� �D6�H6(%2't �d1Q1   ��'    � * a�(Bo�L��L@�(���|, `E�d7���'�Y���R�zT0 k� �<6�@6(%2't �d1Q1   ��'   � * a�(Bg�L��L@�)���|, dE�\6���#�Y���R�zT0 k� �45�85(%2't �d1Q1   ��'    � * a�)Rc�L��L@�)��|, dE�T5����Y���R�zT0 k� �05�45(%2't �d1Q1   ��'    � * a� *R[�L��L@�)��|, dE�L4����Y���R�zT0 k� �(4�,4(%2't �d1Q1   ��'    � * a��*RW�L��L@�*��|, dE�D4����Y���R�zT0 k� � 3�$3(%2't �d1Q1   ��'    � * a��+RS�L��L@�*��|, hE�<3����Y���R�zT0 k� �7�7(%2't �d1Q1   ��'    � * a��+RK�L��L@�*��|, hE�42����Y���R�zT0 k� �;�;(%2't �d1Q1   ��'    � * a��,RG�L��L@�*��|, hE�,2����Y���R�yT0 k� �=�=(%2't �d1Q1   ��'    � * a��-RC�L��L@�+��|, hE�$1�����Y���R�yT0 k� � >�>(%2't �d1Q1   ��'    � * a��.R;�L��L@�+��|, lE�0�����Y���R�yT0 k� ��@��@(%2't �d1Q1   ��'   � * a��.�7�L��L@�+��|, lEQ0�����Y���R�yT0 k� ��9��9(%2't �d1Q1   ��'    � * a��/�3�L��L@�+��|, lEQ/�����Y���R�yT0 k� ��4��4(%2't �d1Q1   ��'    � * a��0�/�L��L@�,��|, lEQ/�����Y���R�yT0 k� ��/��/(%2't �d1Q1   ��'    � * a��1�'�L��L@�,��|, lEP�.������Y���R�yT0 k� ��+��+(%2't �d1Q1   ��'    � * a��2�#�L��L@�,��|, pEP�.������Y���R�xT0 k� ��)��)(%2't �d1Q1   ��'    � * a��2��L��L@�,��|, pEP�-������Y���R�xT0 k� ��'��'(%2't �d1Q1   ��'    � * a��3��L��L@|-��|, pEP�-������Y���R�xT0 k� ��&��&(%2't �d1Q1   ��'    � * a��4��L��L@|-��|, pEP�,�����Y���R�xT0 k� ��$��$(%2't �d1Q1   ��'    � * a��5��L��L@|-��|, pEP�+�����Y���R�xT0 k� ��#��#(%2't �d1Q1   ��'   � * a�x6��L��L0|-��|, tEP�+�����Y���R�xT0 k� ��"��"(%2't �d1Q1   ��'    � * a�p7��Lt�L0|.��|, tEP�*�����Y���R�xT0 k� ��!��!(%2't �d1Q1   ��'    � * a�h8��Lt�L0x.��|, tEP�*�����Y���R�xT0 k� �� �� (%2't �d1Q1   ��'    � * a�`9��Lt�L0x.��|, tE@�*�����Y���R�wT0 k� ����(%2't �d1Q1   �'    � * a�X9���Lt�L0x.��|, tE@�*�����Y���R�wT0 k� ����(%2't �d1Q1   ��'    � * a�P:���Lt�L0t//��|, xE@�)�����Y���R�wT0 k� ����(%2't �d1Q1   ��'    � * a�H;���Lt�E�p//��|, xE@�(�����Y���R�wT0 k� ����(%2't �d1Q1   ��'    � * a�@<���BD�E�l0/��|, xE@�'����ߘY���R�wT0 k� ����(%2't �d1Q1   ��'    � * a�8=���BD�E�h0/��|, xA�&����ߗY���R�wT0 k� �|��(%2't �d1Q1   ��'    � * a�0>���BD�E�d1/��|, xA�%����ۗY���R�wT0 k� �p�t(%2't �d1Q1   ��'    � * a�(?���BD�E�`2/��|, xA�$����זY���R�wT0 k� �h�l(%2't �d1Q1   ��'    � * a� @���BD�E�\2/��|, |A�#����זY���R�wT0 k� �\�`(%2't �d1Q1   ��'    � * a�A���BD�E�X3/��|, |A�"����ӕY���R�vT0 k� �T�X(%2't �d1Q1   ��'    � * a�B���BD�E�X4/��|, |A�!����ӕY���R�vT0 k� �P�T(%2't �d1Q1   ��'    � * a	rC���BD�E�T4/��|, |A� ����ϔY���R�vT0 k� �H�L(%2't �d1Q1   ��'    � * a	rD���BD�E�P5/��|, |A|����ϔY���R�vT0 k� �D�H(%2't �d1Q1   ��'    � * a	q�E���BD�E�L6���|, |At�ӿ�ϓY���R�vT0 k� �<�@(%2't �d1Q1   ��'    � * a	q�F���BD�E�H7���|, �Ap�ӿ�˓Y���R�vT0 k� �4�8(%2't �d1Q1   ��'    � * a	q�F���BD�F D8���|, �Ah�Ӿ�˓Y���R�vT0 k� �0
�4
(%2't �d1Q1   ��'    � * a	��G���BD�F D9���|, �Ad�׽�ǒY���R�vT0 k� �(	�,	(%2't �d1Q1   ��'    � * a	��G���BD�F @:���|, �A \�׽�ǒY���R�vT0 k� �(�,(%2't �d1Q1   ��'    � * a	��H���BD�F <;���|, �A X�׼�ÑY���R�vT0 k� �$�((%2't �d1Q1   ��'    � * a	��H��BD�F <<���|, �A P�׼�ÑY���R�vT0 k� �� (%2't �d1Q1   ��'    � * a	��I��BD�F 8=���|, �A H�׻���Y���R�uT0 k� ��(%2't �d1Q1   ��'    � * a	q�I��BD�F 8>���|, �A D�׻���Y���R�uT0 k� ��(%2't �d1Q1   ��'    � * a	q�J��BD�F 8@���!�, �A <�׻���Y���R�uT0 k� ��(%2't �d1Q1   ��'    � * a	q�J��BD�F 4A���!�, �A 4�׺���Y���R�uT0 k� � � (%2't �d1Q1   ��'    � * a	q�J��BD�F 4B���!�, �A 0�׺���Y���R�uT0 k� �����(%2't �d1Q1   ��'    � * a	q�K��BD�E�4C��!�, �A (�׺���Y���R�uT0 k� ������(%2't �d1Q1   ��'    � * a	��K��BD�E�0D��!�, �A $�׹���Y���R�uT0 k� ������(%2't �d1Q1   ��'    � * a	��K��BD�E�0E�!�, �A �׹���Y���R�uT0 k� ������(%2't �d1Q1   ��'    � * a	��K��BD�E�0F�!�, �A0�׹���Y���R�uT0 k� ������(%2't �d1Q1   �'    � * a	��K��BD�E�0G�!�, �A0 �׹���Y���R�uT0 k� ������(%2't �d1Q1   ��'    � * a	��K��BD�E�0H�!�, �A0 �׸���Y���R�uT0 k� ������(%2't �d1Q1   ��'    � * a	q�K��BD�E�0J�!�, �A0 �׸���Y���R�uT0 k� ������(%2't �d1Q1   ��'    � * a	q�K��BD�E�0K�!�, �A0 �׸���Y���R�uT0 k� ������(%2't �d1Q1   ��'    � * a	q�K��BD�B�4L�|, �A0 �׷���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * a	q�K��BD�B�4M�|, �A0$�׷���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * a	q�K��BD�B�4N�|, �A0$�׷���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * aA�K��BD�B�8O�|, �A0$�׷���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * aA�L��BD�B�8P�	|, �A0$�׶���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * aA�L��BD�B�8P�
|, �A0$�׶���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * aA�L��BD�B�<Q�
|, �A@$�׶���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * aA�L��BD�B�@R�
|, �A@(�׶���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * a1�M��BD�B�@S��|, �A@(�׵���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * a1�M��BD�B�DT��|, �A@(�׵���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * a1�Mу�BD�B�HU��|, �A@(�׵���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * a1�N��BD�B�HV��!�, �G�(�׵���Y���R�tT0 k� ������(%2't �d1Q1   ��'    � * a1�N��BD�B�LW��!�, �G�(�״���Y���R�tT0 k� ����(%2't �d1Q1   ��'    � * aфN�{�BD�B�PW��!�, �G�(�״���Y���R�tT0 k� ����(%2't �d1Q1   ��'    � * aрN�{�BD�B�TX��!�, �G�(�״���Y���R�tT0 k� ����(%2't �d1Q1   ��'    � * aрO�w�BD�B�XY��!�, �G�(�״���Y���R�tT0 k� ����(%2't �d1Q1   ��'    � * a�|OAw�BD�B�\Z��!�, �G�(�׳���Y���R�tT0 k� ����(%2't �d1Q1   ��'    � * a�xOAs�BD�B�`[��!�, �G�(�׳���Y���R�tT0 k� ����(%2't �d1Q1   ��'    � * a�xPAs�BD�B�d[��!�, �G�(�׳���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�tPAo�BD�B�h\��!�, �G�,�׳���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�pPAo�BD�B�l]��!�, �G�,�׳���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�pPAo�BD�B�p^��!�, �G�,�ײ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�lQAk�BD�B�x^��|, �G�,�ײ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�lQAk�BD�B�|_��|, �G�,�ײ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�hQAg�BD�B��`��|, �G�,�ײ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�hQAg�BD�B��a��|, �G�,�ײ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�dRAc�BD�B��a��|, �G�,�ױ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�dRAc�BD�B��b��|, �G�,�ױ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�`RQc�BD�B��c��|, �G�,�ױ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�`RQ_�BD�B��c��|, �G�,�ױ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�\SQ_�BD�B��d��|, �G�,�ױ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�\SQ_�BD�B��d��|, �G�,�Ӱ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�XSQ[�BD�B��e��|, �G�,�Ӱ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�XS�[�BD�B��f��|, �G�0�Ӱ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�TT�[�BD�Bмf��|, �G�0�Ӱ���Y���R�sT0 k� ����(%2't �d1Q1   ��'    � * a�TT�W�BD�B��g��|, �G�0�Ӱ���Y���R�sT0 k� ��	��	(%2't �d1Q1   ��'    � * a�PT�W�BD�B��g��|, �G�0�Ӱ���Y���R�sT0 k� ��
��
(%2't �d1Q1   ��'    � * a�PT�S�BD�B��h��|, �G�0�Ӱ���Y���R�sT0 k� ��
��
(%2't �d1Q1   ��'    � * a�LT�P BD�B��i��|, �G�0�ӯ���Y���R�sT0 k� ��
��
(%2't �d1Q1   ��'    � * a�LU�PBD�E��i��|, �G�0�ӯ���Y���R�sT0 k� ��
��
(%2't �d1Q1  �'    � * a�HU�LBD�E��j��|, �G�0�ӯ���Y���R�sT0 k� ��
��
(%2't �d1Q1  ��/    � * a�HU�LBD�E��j��|, �G�0�ӯ���Y���R�sT0 k� ��
��
(%2't �d1Q1  ��/    � * a�DU�LBD�E��k��|, �G�0�ӯ���Y���R�sT0 k� ��
��
(%2't �d1Q1  ��/    � * a�DU�LLt�E��k��|, �G�0�ӯ���Y���R�sT0 k� ��
��
(%2't �d1Q1  ��/    � * a�DV�HLt�E�l��|, �G�0�Ӯ���Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�@V�HLt�E�l��|, �G�0�Ӯ���Y���R�rT0 k� �l
�p
(%2't �d1Q1  ��/    � * a�@V�HLt�E�m��|, �G�0�Ӯ��Y���R�rT0 k� �X
�\
(%2't �d1Q1  ��/    � * a�<V�DLt�E�m�� |, �G�0�Ӯ��Y���R�rT0 k� �D
�H
(%2't �d1Q1  ��/    � * a�<V�DLt�E�$n�� |, �G�0�Ӯ��Y���R�rT0 k� �0
�4
(%2't �d1Q1 	 ��/    � * a�<W�D	Lt�E�,n�� |, �G�4�Ӯ��Y���R�rT0 k� � 
�$
(%2't �d1Q1 	 ��/    � * a�8W�@
Lt�E�<o��!|, �G�4�Ӯ��Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�8W�@Lt�E�Do��"|, �G�4�ӭ��Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�4W�@Lt�E�Po��"|, �G�4�ӭ�{�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�4W�<Lt�E�Xp��"|, �G�4�ӭ�{�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�4X�<Lt�E�`p��#|, �G�4�ӭ�{�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�0X�<Lt�E�hp��#|, �G�4�ӭ�{�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�0X�<L��E�pp��#|, �G�4�ӭ�{�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�0X�8L��E�xp��$|, �G�4�ӭ�{�Y���R�rT0 k� �l
�p
(%2't �d1Q1  ��/    � * a�,X�8L��E��p��$|, �G�4�ӭ�{�Y���R�rT0 k� �X
�\
(%2't �d1Q1  ��/    � * a�,X�8L��E��p��$|, �G�4�ӭ�w�Y���R�rT0 k� �D
�H
(%2't �d1Q1  ��/    � * a�,Y�8L��E��p��%|, �G�4�Ӭ�w�Y���R�rT0 k� �0
�4
(%2't �d1Q1  ��/    � * a�(Y�8L��E��p��%|, �G�4�Ӭ�w�Y���R�rT0 k� � 
�$
(%2't �d1Q1  ��/    � * a�(Y�4L��E��p��%|, �G�4�Ӭ�w�Y���R�rT0 k� �
�
(%2't �d1Q1  ��/    � * a�(Y�4L��E��p��&|, �G�4�Ӭ�w�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�$Y�4L��E��p��&|, �G�4�Ӭ�w�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�$Y�4L��E��o��&|, �AP4�Ӭ�w�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�$Y�0L��E��o��'|, �AP4�Ӭ�w�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a�$Z�0L��E��n��'|, �AP4�Ӭ�s�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * a� Z�0L��E��n��'|, �AP4�Ӭ�s�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * aA Z�0L��E��m��(|, �AP4�Ӭ�s�Y���R�rT0 k� ��
��
(%2't �d1Q1  ��/    � * aA Z�0L��E��m��(|, �AP8�ӫ�s�Y���R�rT0 k� �l
�p
(%2't �d1Q1  ��/    � * aAZ�,L��K��l��)|, �AP8�ӫ�s�Y���R�rT0 k� �X
�\
(%2't �d1Q1  ��/    � * aA[�,L��K��l��)|, �AP8�ӫ�s�Y���R�rT0 k� �D
�H
(%2't �d1Q1  ��/   � * aA[�,L��K��k/�)|, �AP8�ӫ�s�Y���R�rT0 k� �0
�4
(%2't �d1Q1  ��/    � * a� 3�FWE�DE�D�\�A� �<���Z3����T0 k� @f�Df(%2't �d1Q1   ��" 
   � <�J� 3�F WE�@F�D�\�A� �<���Z3���T0 k� �He�Le(%2't �d1Q1   ��" 
   � <�L��3�F$XE�8G�H�\�
A� �;���Z3���T0 k� �Pe�Te(%2't �d1Q1   ��" 
   � <�O��3�F(XE�4H�H�\�BM �;���Z3���T0 k� �Tf�Xf(%2't �d1Q1   ��" 
   � <�R��7�E�0YE�(J�P�	�|BM �p:���Z3���~T0 k� �Xc�\c(%2't �d1Q1   ��" 
   � <�U��;�E�4YE�$K�T�	�tBM �h9���Z3���~T0 k� �X`�\`(%2't �d1Q1   ��" 
   � <�X��;�E�8ZE� M�\�	�pBM �`9���Z3���~T0 k� �\^�`^(%2't �d1Q1   ��" 
   � <�[��?�E�<ZE�N�\�	�l D� �X8���Z3���}T0 k� �\]�`](%2't �d1Q1   ��"    � <�^��?�E�DZE�O�`�	�g�D� �P8���Z3���x}T0 k� �`\�d\(%2't �d1Q1   ��"    � <�a��C�@-H[E�Q�d�	�c�D��H7��Z3���p}T0 k� �t\�x\(%2't �d1Q1   ��"    � <�e �G�@-T\E�S�p�	�[�D��<5��Z3���`|T0 k� ��\��\(%2't �d1Q1   ��"    � <�i�K�@-X\FU�t�	�S�D��44��Z3���X|T0 k� ��]��](%2't �d1Q1   ��"    � <�m�O�@-`\F V�x�	�O�D��,4��Z3���P|T0 k� ��]��](%2't �d1Q1   ��"    � <�q�S�E�d]F�X��
�	�K�F�$3��Z3���H|T0 k� ��\��\(%2't �d1Q1   ��"    � <�u�W�E�l]F�Y��	�	�G�F� 2��Z3���@|T0 k� ��\��\(%2't �d1Q1   ��"    � <�y�_�E�x^F�\���	�?�F�0��Z3���0{T0 k� ��\��\(%2't �d1Q1   ��"    � <�}�c�E��^F�^���	�?�F�.�#�Z3���({T0 k� ��]��](%2't �d1Q1   ��"    � <�� �g�E��^F�`���	�;�F-�'�Z3��� {T0 k� ��]��](%2't �d1Q1   ��"    � <��-$�k�E��_F�a���	�7�F ,�/�Z3���{T0 k� ��]��](%2't �d1Q1   ��"    � <��-(�o�E��_F�c���	�3�E��+�3�Z3���zT0 k� ��^��^(%2't �d1Q1   ��"    � <��-,�s�E��_F�d���	�/�E� �*�;�Z3���zT0 k� ��^��^(%2't �d1Q1   ��"    � <��-0�w�E��`F�f�� �	�/�E� �(�?�Z3��� zT0 k� ��^��^(%2't �d1Q1   ��"    � <��-<̓�E��`E��i����	�+�E�( �&�K�Z3����yT0 k� ��_��_(%2't �d1Q1   ��"    � <��@͇�E��aE��k����	�'�B�,!�$�S�Z3����yT0 k� ��[��[(%2't �d1Q1   ��"    � <��D͏�E��aE��m����	�'�B�0"�#�[�Z3����yT0 k� ��X��X(%2't �d1Q1   ��"    � <��L͓�E��aE��n����	�#�B�4#�"�_�Z3����xT0 k� ��W��W(%2't �d1Q1   ��"    � <��P	͛�E��aE��p����	�#�B�<$� �g�Z3����xT0 k� ��U��U(%2't �d1Q1   ��"    � <��X	͟�E��aE��q����	�#�B�@$���o�Z3��^�xT0 k� ��T� T(%2't �d1Q1   ��"    � <��\
ݧ�E��aE��s����	��B�D%���w�Z3��^�wT0 k� �S�S(%2't �d1Q1   ��"    � <��d
ݫ�E��aE��t������B�H&����Z3��^�wT0 k� �R�R(%2't �d1Q1   ��"    � <��hݳ�E��aE��u������B�P'��̇�Z3��^�wT0 k� �Q�Q(%2't �d1Q1   ��"    � <��pݷ�E� `E��v������B�T'��̏�Z3��^�vT0 k� � Q�$Q(%2't �d1Q1   ��"    � <��|�ǚ@~`E��v������B�l)��ܛ�Z3��^�vT0 k� �0O�4O(%2't �d1Q1   ��"    � <�����˚@~`E��v������B�x*��ܣ�Z3��^�uT0 k� �8L�<L(%2't �d1Q1   ��"    � <�����Ӛ@~$_E��w������B��*��ܯ�Z3��^�uT0 k� �DK�HK(%2't �d1Q1   ��"    � <�����ۚ@~,_E��w������B��+��ܷ�Z3��^�uT0 k� �LJ�PJ(%2't �d1Q1   ��"    � <������@~8_E��w������B��,��ܿ�Z3��^|tT0 k� �TH�XH(%2't �d1Q1   ��"    � <������@~@^B��w���� ��B��,���ǀZ3��^ttT0 k� �\G�`G(%2't �d1Q1   ��"    � <������@~H^B��w���� ��B��-���ρZ3��^ltT0 k� �hG�lG(%2't �d1Q1   ��"    � <�������@~P]B� v���� ��B��.���ׁZ3��^dsT0 k� �pF�tF(%2't �d1Q1   ��"    � <�������@~\]B�v��� ��B��.���߁Z3��N\sT0 k� �xF�|F(%2't �d1Q1   ��"    � <������@~l\B�v��� �B��0����Z3��NLsT0 k� ��E��E(%2't �d1Q1   ��"    � <������@~t[B�v��� �B��0��
���Z3��NDsT0 k� ��D��D(%2't �d1Q1   ��"    � <������@�|[E�u��� �B��1��	��Z3��N<sT0 k� ��E��E(%2't �d1Q1   ��"    � <�����'�@��ZE� u��| �B��2����Z3��N4rT0 k� ��D��D(%2't �d1Q1   ��"    � <�����/�@��ZE�$u��| �B� 2����Z3��N,rT0 k� ��D��D(%2't �d1Q1   ��"    � <�����7�@��YE�(t���| �B�3����Z3��N$rT0 k� ��C��C(%2't �d1Q1   ��"    � <�����?�@��YE�0t��| �B�3���#�Z3��NrT0 k� ��C��C(%2't �d1Q1   ��"    � <�����G�E�XE�4s��| �B� 4���+�Z3��NsT0 k� ��I��I(%2't �d1Q1   ��"    � <����[�E�WE�@r��| �B�05���;�Z3��N sT0 k� ��M��M(%2't �d1Q1   ��"    � <����c�E�WE�Dr��| �B�86���C�Z3��=�sT0 k� ��P��P(%2't �d1Q1   ��"    � <��� �k�E�VE�Lq��|$��B�D6�� �K�Z3��=�sT0 k� ��S��S(%2't �d1Q1   ��"    � <���(�s�E�VE�Pq��|$��B�L7�� �W�Z3��=�rT0 k� ��T��T(%2't �d1Q1   ��"    � <���0�{�E�UE�Xp��|$��B�T7����_�Z3��=�rT0 k� ��U��U(%2't �d1Q1   ��"    � <���8���E�UE�\o�#�|$��B�\8����g�Z3��=�rT0 k� ��U��U(%2't �d1Q1   ��"    � <���D���E�TE�`o�'�|$��B�d8����o�Z3��=�rT0 k� �V�V(%2't �d1Q1   ��"    � <���L���E�TE�hn�+�|$��B�l9����w�Z3��=�rT0 k� �V�V(%2't �d1Q1   ��"    � <���T���E SE�lm�/�|$��B�t9�����Z3��=�rT0 k� �V�V(%2't �d1Q1   ��"    � <���d���ERE�xk�7�|$��B��:������Z3��=�rT0 k� �$U�(U(%2't �d1Q1   ��"    � < �lγ�ERE�|j�;�|$��B��;������Z3��=�rT0 k� �,U�0U(%2't �d1Q1   ��"    � < �xλ�E$QE��i�C�|$��B��;N�����Z3��=�rT0 k� �4U�8U(%2't �d1Q1   ��"    � < ���ǚE,QCL�h�G�|$�#�B��<N�����Z3��-�rT0 k� �<U�@U(%2't �d1Q1   ��"    � < 	���ϚE4QCL�g�K�|$�'�B��<N�����Z3��-�rT0 k� �HT�LT(%2't �d1Q1   ��"    � < ���ךE�<PCL�f�O�|$�+�B��=N��ͻ�Z3��-�sT0 k� �PR�TR(%2't �d1Q1   ��"    � < ���ߚE�HPCL�d�S�|$�/�B��=N���ÇZ3��-�sT0 k� �XP�\P(%2't �d1Q1   ��"    � < ����E�POCL�c�[�|$�3�B��>.���ˇZ3��-�sT0 k� �`O�dO(%2't �d1Q1   ��"    � < ����E�XOE��b�_�|$�;�B��>/��ӇZ3��-�sT0 k� �hN�lN(%2't �d1Q1   ��"    � < �����E�`OE��a�c�|$�?�B�?/��ۇZ3��-�tT0 k� �tM�xM(%2't �d1Q1   ��"    � < �����E�hNE��_�g�|$�C�B�?/���Z3��-|tT0 k� �|M��M(%2't �d1Q1   ��"    � < ����E�tNE��^�k�|(�G�B�$?/���Z3��-xuT0 k� ��L��L(%2't �d1Q1   ��"    � < ����E�|ME��]�o�|(�O�B�0@���Z3��-puT0 k� ��H��H(%2't �d1Q1   ��"    � < �� ��E��ME��[�s�|(�S�B�<@����Z3��luT0 k� ��E��E(%2't �d1Q1   ��"    � < ��!��E��ME��Z�w�|(�W�B�HA���Z3��hvT0 k� ��B��B(%2't �d1Q1   ��"    � < !��!�+�E��LE��Y�{�|(�_�B�TA���Z3��dvT0 k� ��@��@(%2't �d1Q1   ��"    � < #��"�3�E��LE��X��|(�c�B�\A#���Z3��`wT0 k� ��>��>(%2't �d1Q1   ��"    � < &��#�;�@�KE��W���|(�k�B�hB�'���Z3��`wT0 k� ��;��;(%2't �d1Q1   ��"    � < ( $�C�@�KE��V���|,�s�B�tB�+��'�Z3���\wT0 k� ��8��8(%2't �d1Q1   ��"    � < *%�K�@�JE��T���|,�w�B��B�/��/�Z3���XxT0 k� ��6��6(%2't �d1Q1   ��"    � < ,%�S�@�IE��S���|,��B��B�7��7�Z3���XxT0 k� ��5��5(%2't �d1Q1   ��"    � < /&�[�@�IE��R���|,̇�O�B�;��?�Z3���TyT0 k� ��3��3(%2't �d1Q1   ��"    � < 2 '�c�@�HE��Q���|,
̋�O�B�?��G�Z3���PyT0 k� ��2��2(%2't �d1Q1   ��"    � < 5((�k�E�HE��P���|,
̓�O�B�G��S�Z3���PyT0 k� ��8��8(%2't �d1Q1   ��"    � < 80)�s�E�HE��O���|,
̛�O�B�K��[�Z3���PzT0 k� ��=� =(%2't �d1Q1   ��"    � < ;8*�{�E�GE��N���|,
̣�O�C�S��c�Z3���LzT0 k� �A�A(%2't �d1Q1   ��"    � < >@*���E�GE��M���|,
���O�C�W��k�Z3���LzT0 k� �C�C(%2't �d1Q1   ��"    � < @H+���EFE��L���|,
���O�C�_��s�Z3���L{T0 k� �E�E(%2't �d1Q1   ��"    � < BP,���E�FE��K���|,	���O�C�c��{�Z3���H{T0 k� �$@�(@(%2't �d1Q1   ��"    � < DX-���E�FE��J���|,	�ÛO�C�k����Z3���H{T0 k� �0=�4=(%2't �d1Q1   ��"    � < F`.���E� EE��I���|,	�˚O�C�s����Z3���H|T0 k� �8;�<;(%2't �d1Q1   ��"    � < Hh/���E�(EE��H���|,	�әO�C�w����Z3���H|T0 k� �@9�D9(%2't �d1Q1   ��"    � < Jp0���E�0DE� G���|,�ۘO�C�����Z3���H|T0 k� �H8�L8(%2't �d1Q1   ��"    � < Lx1���E�8DE� F���|,��O�C������Z3���H}T0 k� �T6�X6(%2't �d1Q1   ��"    � < N�2�ǚE�DCE�F���|,��O�D������Z3���H}T0 k� �\5�`5(%2't �d1Q1   ��"    � < P�3�ϚE�LCE�E���|,��O�D������Z3���H}T0 k� �d4�h4(%2't �d1Q1   ��"    � < R�4�ךE�TBE�D���|,���O D������Z3���L~T0 k� �l3�p3(%2't �d1Q1   ��"    � < T�5�ߚ@p\AE�C���|,��OD����ǋZ3� �L~T0 k� �x0�|0(%2't �d1Q1   ��"    � < V�6��@pdAE�B���|,��ODϫ��ϋZ3� �L~T0 k� ��-��-(%2't �d1Q1   ��"    � < X�7��@pl@E�A���|,��ODϳ��׋Z3� �LT0 k� ��,��,(%2't �d1Q1   ��"    � < Z/�8���@px@E�A���|,��ODϻ��ߋZ3� �PT0 k� ��*��*(%2't �d1Q1   ��"    � < \/�9��@p�?E�@���|,�'�O$D�����Z3� �PT0 k� ��(��((%2't �d1Q1   ��"    � < ^/�:��@p�>E�?���|,�/�O(D�����Z3��TT0 k� ��'��'(%2't �d1Q1   ��"    � < `/�;��@p�>E� >���|,�;�O0D������Z3��T�T0 k� ��&��&(%2't �d1Q1   ��"    � < b/�<��@p�=E�$=���|,�C�O4E�����Z3��XT0 k� ��%��%(%2't �d1Q1   ��"    � < d/�=�#�@p�<E�$=���|,�K�O<E�����Z3��XT0 k� ��$��$(%2't �d1Q1   ��"    � < f/�>�+�@p�;E�(<���|,�S�O@E�����Z3��\T0 k� ��$��$(%2't �d1Q1   ��"    � < h/�@�3�@p�;E�,;���|,�_�E�HE�����Z3��\T0 k� ��#��#(%2't �d1Q1   ��"    � < j/�A�;�@p�:E�,:���|,�g�E�PE����#�Z3��`~T0 k� ��"��"(%2't �d1Q1   ��"    � < l/�B�C�@��9E�0:���|,�o�E�TE���+�Z3��d~T0 k� ��"��"(%2't �d1Q1   ��"    � < n/�C�K�@��8E�09���|,�w�E�`E� �7�Z3��d~T0 k� ��"��"(%2't �d1Q1   ��"    � < p�D�S�@��7E�48���|,���E�pE� �?�Z3��h~T0 k� ��"��"(%2't �d1Q1   ��"    � < r�E�[�@��7E�88���|,���B�|E� �G�Z3��l~T0 k� ��!� !(%2't �d1Q1   ��"    � < t�F�g�@��6E�87���|,���B��E�$ �O�Z3��p}T0 k� � � (%2't �d1Q1   ��"    � < v�H�o�@��5E�<6���|,��B��E�, �W�Z3��t}T0 k� ��(%2't �d1Q1   ��"    � < x�$I�w�@��4E�<6���|,��B��F�4 �_�Z3��x}T0 k� ��(%2't �d1Q1   ��"    � < z�,J��@��3E�@5���|,��B��F�< �g�Z3��|}T0 k� �� (%2't �d1Q1   ��"    � < |�4KЇ�@�2E�D5���|,��B��F�D �o�Z3�݀|T0 k� �$�((%2't �d1Q1   ��"    � < ~�<LЋ�@�1E�D4���|,ÖB��F�L �w�Z3�݄|T0 k� �0�4(%2't �d1Q1   ��"    � < ��@M	�@�0E�H3���|,ϗB��F�T σ�Z3���|T0 k� �8�<(%2't �d1Q1   ��"    � < ��HO	�@� /E�H3��|,חB��F�\ ϋ�Z3���|T0 k� �@�D(%2't �d1Q1   ��"    � < ��PP	�@�(/E�L2��|,ߘB��F�d ߓ�Z3���|T0 k� �H�L(%2't �d1Q1   ��"    � < ��XQ	�@�0.E�L2��|,�B��F�l ߛ�Z3���{T0 k� �P�T(%2't �d1Q1   ��"    � < � `R	�@�8-E�P1��|,�B��F�t ߣ�Z3���{T0 k� �X�\(%2't �d1Q1   ��"    � < � hS
 ��@�@,E�P1��|,��B�F�| ߫�Z3���{T0 k� �`�d(%2't �d1Q1   ��"    � < � pU
 ��@�H+E�T0��|,�B�F��߳�Z3���{T0 k� �h�l(%2't �d1Q1   ��"    � < � tV
 ��@�P*E�T/��|,�B�F��߻�Z3���{T0 k� �p�t(%2't �d1Q1   ��"    � < � |W
 ×@�X)E�X/��|,�B�$F���ÎZ3���{T0 k� �x�|(%2't �d1Q1   ��"    � < ��X
 Ǘ@�`(E�X.��|,#�B�,F���ˎZ3���zT0 k� ����(%2't �d1Q1   ��"    � < ��Z�ϗ@�h'E=\.��|,+�B�4G���׎Z3���zT0 k� ����(%2't �d1Q1   �"    � < ��[�ӗ@�p%E=\->�|,3�B�@G���ߎZ3���zT0 k� ����(%2't �d1Q1   ��"    � < ��\�ז@�x$E=`->�|,?�B�HG����Z3���zT0 k� ����(%2't �d1Q1   ��"    � < ��]�ߖ@��#E=`,>�|,G�B�PG����Z3���zT0 k� ����(%2't �d1Q1   ��"    � < ��^��@��"E=d+>�|,O�B�\G�����Z3���zT0 k� ����(%2't �d1Q1   ��"    � < ��_��@��!E-d*>�|,[�B�dG�����Z3���yT0 k� ����(%2't �d1Q1   ��"    � < ��`��@�� E-h*.�|,c�B�lG����Z3���yT0 k� ����(%2't �d1Q1   ��"    � < ��a��@��E-h).#�|,k�E�tG����Z3���yT0 k� ����(%2't �d1Q1   ��"    � < ��bp��@��E-l(.#�|,w�E�|G����Z3���yT0 k� ����(%2't �d1Q1   ��"    � < ���cp��@��E-p'.'�|,�E��G���#�Z3���yT0 k� ����(%2't �d1Q1   ��"    � < ���dq�@��B�t&.+�|,��E��G���+�Z3���yT0 k� ����(%2't �d1Q1   ��"    � < ���fq�@��B�x%�/�|,���E��G��;�Z3�� xT0 k� ����(%2't �d1Q1   ��"    � < ���g��@q�B�|$�3�|,���E��G��C�Z3��xT0 k� ����(%2't �d1Q1   ��"    � < ���h��@q�B��#�7�|,���E��G��K�Z3��xT0 k� ����(%2't �d1Q1   ��"    � < �� i��@q�B��#�;�|,���E��G�(�S�Z3��xT0 k� ����(%2't �d1Q1   ��"    � < ��j�'�@q�B��"�?�|,���E��G�0�[�Z3��xT0 k� ����(%2't �d1Q1   ��"    � < ��k�+�@q�B��!�C�|,�˨E��G�8�c�Z3��$xT0 k� ����(%2't �d1Q1   ��"    � < ��l3�@q�B�� �G�|,�өE��G�D�k�Z3��,xT0 k� ����(%2't �d1Q1   ��"    � ; �� m7�@q�B�� �K�|,�۩E��G�L�w�Z3��0wT0 k� ����(%2't �d1Q1   ��"    � : ��(n;�@rB���O�|,��@a�G�T��Z3��8wT0 k� �#��'�(%2't �d1Q1   ��"    � 9 ��<pG�@rB���[�|,���@a�G�h���Z3��HwT0 k� �3��7�(%2't �d1Q1   ��"    � 8 ��DpO�@rB���_�|,��@a�G�p���Z3� �PwT0 k� �;��?�(%2't �d1Q1   ��"    � 7 ��LqS�@r B���c�|,��@a�H�|���Z3� �XwT0 k� �C��G�(%2't �d1Q1   ��"    � 6 ��Tr�[�@�(
B���k�|,��@bHф���Z3� �`wT0 k� �K��O�(%2't �d1Q1   ��"    � 5 ��\s�c�@�0	B���o�|,��@bHь���Z3� �hwT0 k� �S��W�(%2't �d1Q1   ��"    � 4 �dt�g�@�8B���s�|,�'�@bHј���Z3� �pwT0 k� �[��_�(%2't �d1Q1   ��"    � 3 �lt�o�@�@B���{�|,�3�@bHѠ�ÏZ3� �xvT0 k� �c��g�(%2't �d1Q1   ��"    � 2 �tu�s�@�HB����|,�;�@b HѨ�ːZ3� ހvT0 k� �k��o�(%2't �d1Q1   ��"    � 1 ��w���EXB�����|,�O�@b0HѼ�ېZ3� ސvT0 k� �w��{�(%2't �d1Q1   ��"    � 0 ��x���E\B�����|,�W�@b4H����Z3��ޘvT0 k� �{���(%2't �d1Q1   ��"    � / ���x���Ed B�����|,�c�@b<H����Z3��ޠvT0 k� �����(%2't �d1Q1   ��"    � . ���y���Eo�B�����|,�k�@bDH����Z3��ިvT0 k� ������(%2't �d1Q1   ��"    � - ���z���Ew�B��Σ�|,�s�@bHH�����Z3����vT0 k� ������(%2't �d1Q1   ��"    � , ���z���E�B��Ϋ�|,��EPH ���Z3����vT0 k� ������(%2't �d1Q1   ��"    � + ���{���E��B�ί�|,χ�ETH ���Z3����uT0 k� ������(%2't �d1Q1   �"    � * ���{���FB��B�η�|,ϓ�E\H ���Z3����uT0 k� ������(%2't �d1Q1   ��/    � ) ���|���FB��B�ο�|,ϛ�EdH ��Z3����uT0 k� ������(%2't �d1Q1   ��/    � ( ���}�ǂFB��B����|,���ElH �'�Z3����uT0 k� ������(%2't �d1Q1   ��/    � ' ���}�ςFB��B�$���|,���EtH �/�Z3����uT0 k� ����(%2't �d1Q1   ��/    � & ���~�ׂFB��B�,���|,���ExH �7�Z3����uT0 k� ���#�(%2't �d1Q1   ��/    � % ���~�߂FB��B�4���|,���E�H $�?�Z3����uT0 k� �7��;�(%2't �d1Q1   ��/    � $ �����FR��B�<���|,�˶E�H ,�G�^����uT0 k� �O��S�(%2't �d1Q1   ��/    � # �����FR��B�D���|,�ӷE�H 4�O�^��� uT0 k� �g��k�(%2't �d1Q1   ��/    � " ������FR��B�L���|,�۷E�H <�W�^���uT0 k� �����(%2't �d1Q1   ��/   � ! ������FR��B�T���|,��E��H D�c�^���uT0 k� ������(%2't �d1Q1   ��/    �   ����FR��B�\���|,��E��H L�k�^���uT0 k� ������(%2't �d1Q1   ��/   �  ����Fb��B�d��|,���E��H T�s�^��� tT0 k� ������(%2't �d1Q1   �/    �  ��0~�Fb��B�t��|,��E��H `�^���0tT0 k� 3�����(%2't �d1Q1   ��/    �  ��8~'�Fb��B�|��|,��E��H h�^���8tT0 k� 3�����(%2't �d1Q1   ��/    �  ��@~/�Fb��Bބ�'�!�,��E��I p���^���@tT0 k� 3�����(%2't �d1Q1   ��/    �  ��H};�Fb��Bތ�/�!�,�'�F�I x���^���HtT0 k� 3�����(%2't �d1Q1   ��/    �  ��P}C�Fb��Bޔ�7�!�,�/�F�I�|���^���PtT0 k� 3�����(%2't �d1Q1   ��/    �  ��X|K�Fc�B���?�!�,�7�F�J�����^���XtT0 k� ������(%2't �d1Q1   ��/   �  ��d|S�Fc�B���K�!�,�C�F�J�����^���`tT0 k� ������(%2't �d1Q1   ��/    �  ��l{[�Fc�B���S�!�,�K�F�J�����^���htT0 k� ������(%2't �d1Q1   ��*    �  ��t{�c�Fc�B���[�!�, S�E� K���×^���ptT0 k� ������(%2't �d1Q1   ��*    �  �҄z�s�Fc#�B��
�k�!�, g�E�K2��Ә^��πtT0 k� ������(%2't �d1Q1   ��*    �  �Ҍy�{�Fc'�B��
�s�!�, o�E�L2��ۘ^��ψtT0 k� ������(%2't �d1Q1   ��*    �  ���x���Fc+�B��	�{�!�, w�E�$L2���^��ϐsT0 k� ������(%2't �d1Q1   ��*    �  ���x���Fc3�I�	���|,��I(L2���^��ϘsT0 k� ������(%2't �d1Q1   ��*    �  ���w���Fc7�I�	���|,���I0M2���^��ϠsT0 k� ������(%2't �d1Q1   ��*    �  ���w���Fc;�I����|,���I8MB����^��ϨsT0 k� ������(%2't �d1Q1   ��*    �  ���v���Fc?�I����|,���I@MB���^���sT0 k� ������(%2't �d1Q1   ��*    �  ���v���FcG�I����|,���IDMB���^���sT0 k� ������(%2't �d1Q1   ��*    �  ���u�FcK�I ��|,���ILMB���^���sT0 k� ������(%2't �d1Q1   ��*    �  ���t�ÌES�I/��|,���I#XMB���^���sT0 k� ������(%2't �d1Q1   ��*    �  ���t�ˍE[�I/��|,���I#\M2��'�^���sT0 k� ������(%2't �d1Q1   ��*    �  ���s�ӍE_�I/��|,���I#dM2��/�^���sT0 k� ������(%2't �d1Q1   ��*    �  ���s�ێEg�I/��|,���I#hM2��3�^���sT0 k� ������(%2't �d1Q1   ��*    �  ��r��Ek�I/ ��!�,���I#pM2��;�^���sT0 k� ������(%2't �d1Q1   ��*    �  �r��Es�I(��!�,���ItM3 �C�^���sT0 k� ������(%2't �d1Q1   ��*    �  �q��Ew�I,��!�,���IxM��G�^�� sT0 k� ������(%2't �d1Q1   ��*    �  � q��E��I4��!�,���I�M��S�_3���sT0 k� ������(%2't �d1Q1   ��*    �  �(p��E��I8�!�,��I�M��[�_3���rT0 k� ������(%2't �d1Q1   ��*    �  �0p��E��I/<��!�,��I#�M��_�_3��� rT0 k� ������(%2't �d1Q1   ��*    �  �<o��E���I/@��!�,��I#�M� �g�_3���(rT0 k� ������(%2't �d1Q1   ��*    �  �Do�#�E���I/D��!�,��I#�M�(�k�_3���0rT0 k� ������(%2't �d1Q1   ��*    �  ��Ln�+�E���I/H�'�!�,�#�I#�M�,�o�_s���8rT0 k� ������(%2't �d1Q1   ��*    �  ��\n�;�E���IL�;�!�,�3�I�M�8�{�_s���LqT0 k� ������(%2't �d1Q1   ��*    �  ��dm�?�E���IP�C�|,�;�I�M�@	��_s���PqT0 k� ������(%2't �d1Q1   ��*    �  ��lm�G�D���IT�K�|,�?�I�M�D	�_s���XqT0 k� ������(%2't �d1Q1   ��*    �  �                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��_R ]�&H&G � �� [��   4 4   � GyN     [6  G�b    ��,            ,
  Z a          Pb     ���  8	(          m   � �	   � K�&     �� K�:    a�,                	 Z a�        ���    ���   @
"          ���/  � $       ��    ��� �k    � �               Z a         j��    ���    		'
           k�G  � �   }�     l< {R    ���                S Z a          p�   
  ���  8		           )�&   R R
     .��|�     ){���A�    ,                 6
  Z a          ��b     ��� X
          dx  ��     B�<D     dx�<D                           �����         �`   �  ���    0 0	            �;           V g��     �; g�       �           	 ��           �0  �  ��@   8�	          ��   
	  j #�     �� �     � �                 ��          �P      ��H   (
           ����         ~ ��X    ��φ ��X    ��                      �          �  �  ��@   (           ��T�          ���O�    ��67��j    ��q               @��         	 �@     ��@   0

	 
         �ۑ��     � ��    �۠, ��R    � �                      �� `       
         ��@    8	 1 	            rP        � ��]     rT ��]    ��                    A ��        �0     ��@   P
B 	               ��      �                                                                           �                               ��        ���          ��                                                                 �                          
1)  ��        ��L� (� 
1)�Q�t �  ��r                x                j  �  �   �                          
    ��        ��M       
  �R                                                            �                          G K }��� g  ��� � ����L�M    
   	          
  �   x �� ]-�J       9$ �e� :$  f� :d g  �� d  �� 0d@ �  d� �D d� m� n@ m�  n` m� n���� ����  ����. ����< ����J ����X � J$ ]@ �d �t� �d  u� � v  �d x@ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �� �R� 
�\ U� 
� V  
� V ���� � 
�< W� 
� W����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���� a  *����  ������  
�fD
��L���"����D" � j  "  B   J jF�"     "�j  " ��
��
��"    B�j l �  B �
� �  �  
�      ��     �   �   ��    ��     �           ��     �           � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �/'      �� � � ��        � �T ���        �        ��        �        ��        �   �     F�� 
         ��                         �$ (  ������                                     �                  ����               ���%��   * a�� F �            28 Steve Larmer tu     0:01                                                                        1  1     � �
*� �@C. �PC6
8 C8.kj �N kr � �B�1 � B�A	B�+ 
B�3 �B� � �B� � � B� �B� � �B� � �K( � C> �K7 � K!? �K"2 �K%" � K'! �c�@ � c�HN"� �N "� �>� �>
� ��} ��} �  *&~ � )�v?!� �?"
� � � #*Kv � )�v �%*~ � &*Fv �'*8v �  *Gv � )*Gv �  *Av �  *Av � ,*Fv �-*8v �  *Gv �/*8v �  *Gv �  *AvF 
�D r  *Ou �4
� � {  *Ou ~ 6*Ru ~ *}0 )�tM )�tP )�tA  *Gt2<*8tB  *Gt>*<tD *:t � @"�4 �A�" � 
�1                                                                                                                                                                                                 |� R        �    @ 
        "     W P E ^  ���� 5               �������������������������������������� ���������	�
��������                                                                                          ��    �Y� '  ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, ,�  �@��A�2�                                                                                                                                                                                                                                                                                                                                                   �  ��A,����                                                                                                                                                                                                                                      b    *    ��  4�J      )�  	                           ������������������������������������������������������                                                                                                                                      ��             �          � �             	 
     ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ���                                 /         L�J     Ҁ                             ������������������������������������������������������                                                                                                                                       �    �              z          �
 y             	 	 ���������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������                                                                                                                                                                                                                                                     
                                                                        �             


            �   }�    �                                                            'v                        ������������   &  +
����������������������������   ����������������������������  'r��������������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" A C 6                                 � ,��� �\                                                                                                                                                                                                                                                                                       )n)n1n  
*        a      c      l      c      d      e      m      k                                                                                                                                                                                                                                                                                                                                                                                                           > �  >�  J�  @�  D#�  EZm �̞�� �N ���
����f������������8�����7������     
     <  ���F : k ~ 
         �   & AG� �                ��                                                                                                                                                                                                                                                                                                                                      N I   �                 "         !��                                                                                                                                                                                                                        Y   �� �~ ��      �� 9      ����������������� ������ ������������������������������ ����������� �������������� � �������������������������� � ����� ���������� �������������������� ��������� ������� ������������  �������� ���������������������������� ������������� ��������������� ��� ����������������������� �� ������������������ ����� ������������������  �������� �������������������� ������������������������������ �� ����������� � �� �  � �� � ���������� ���� ������ ������� ���������������     �     $ffllf���flll����llll����ll�l����l��������l�l���fl�Ƹ��ˈ�l���ƪ�˻��˪��˫�̼�ff�f�f��ff�lff���flll���˼ff�̼ffffff�ffffffffffff���̶�ff�fff����flflfl��ffll�fl�lʻ�̻��l̻��˻�l�ll����l�l�����ll����̼��������l�l�����lll�����l�l���ʬƬ�fl��flffff��ffl�f�f�f�f��fˉ�f���f��ffl�ffffffff�fffƬ��Ɖ����ffffffffffff�fffff�ffffffflf�fllfff�ffffffffffffffl�fffl��l�����l������ll��f���fll�����fll�f���ffllff�ffflff��klflj����ffff�ffffffl�fk��f���f�Ƽf�̖f��ff�fl�f��fʨ�����ʩ����̚��l����ll�Ɖ�������˙�����̺���ʙ�f����l��f�k���lj���̛lll�˪̪fˬ��̛�kllll���lll�f���f�l�f���lf��f���ll����l��l�����l��������l������l�f���f���j��ɫ��ɘ��i���i���ʈ�����������������������������������������������������ʋ̼Ɖ��l�����������j���j�������̩���ɩ�̺����f�ƺl�l�f��yl�̙f�ƨ��l�f�ƨ���flf�����ff�l����ffllf���flll����f�{�f�z��ʊ��jy��f����x��ƚ��̙�����������������ʪ��˚��̺���˺����˼fff˺�̚�����˪����������������˪��̪�f���l���˻�ƫ̻l�˻jƨf�ƙl�̊f��{l�̛ll̦���flll����flll����llll����lllf���i�fk��l��lɉ��̩��fj�fff���ƪ��ˊ��i������f�˺���ʬl̪��̉��l�����������������˫�l�������˼�ll�fɼlʩ�������f�ˬ�l��l˛�Ʃ�l̚�ff�˻f�ʙ�lll�����ll�l����l�l�����ffflffff$�I    ;      7      
                       8     �   �����J����      ��     8         �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �f ��        p���� ��   p���� �$ ^h  ��   p   	 ���                  �� �   6   
���(�� x    ����� �    � �$ ^$�� �  �  �� [ 
q~     5���������j � ��� �� � ��� RX� �  �� �       �   d   P���� e����J   g���        f ^�        �� R *      P      ��_��������J���J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  "  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��  DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰ wwwywww�www�www�www�www�www�www����������!��������������������a��������݈����������a������������(-�a������!�-���www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�www�������������������������������������!�����!�-����������!-�����������!������www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�www������m����������݈����������������a݈�����m����!�����������a�-������www�www�www�www�www�www�www�wwwwww�www�www�www�www�www�www�wwwy-��������!�����������������������������������!��������                                          �      �  a r!   f�"""""*��**"*�"�""�""v""*f   "  ""- ��"�"*"-""z"""""����            n   �  "  q  ��                          �  �                                 � gv"!g�vg�vggfvv|�b��r""gb"�vr�rgb��v���g���v���***�*q!q�"!a�!vwfqqr~� qw��q�~~q�����~~~�w~~w�w            �   ~   ��  ~~  �w      v    �                ggj�vvggvvgg!vg�g֪vvg�r�r��⢪rq**gjb�v�q*gjj*vv��gg�z�/�"!�"�*�""*z����qw�~q~ww��q~qwvq�w�`� ��� �w �~p w�p  ��                    �                        lggz�v��g        �       ggbvvrgggavvvqggav� �      ���w!z�w"""�!""*�"! ��        q� q�        `               �        �                      wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p   �   �   	                                       	   �  	   �  	   	   	    �   	�            ����        �   	    �   	    �  	   �  	   �      	   �  	   �  	   �  	   �                   ����   	   	   	   	   	   	   	   	   	   	�  		  	 � 	 	 	  �	  		   �                                           
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  ""   "! " ""            """                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """"! "   "      ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  ""   "! " ""            """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                        � ̻ �ۼͺ�	ۚ����C�˽T;��UJ��ET�35J�D3T�  ̰ ̻	�̻���w���&��wv��wpʨ� ��� ��� ��  "�� .� "�� ��0 "          .  .  "   "             �  �� ʝ ,��+� "" "��CEJ�D5J� J�  �� 
�� �  �� �+� �"" """����    �         ""�"" �  ��                /���"/�  ��                    �                                                                            �               �     "   "                 ���� �                                                   ���                          ����                  �   �� �       �  �  "�  "   "                                                          � ��� ��� ܷz �riwgkww��������"���"��ܽ���̻������������	������J�@T�D                        �   �   �"  "  "  " � � � �  �  ��  ��  "   "   "   "           UJ�@T�DT�TUJ� 5J� �J� �˻�˰ ܩ� ,ʠ "����, �""�"" � ��               /�� "     � �        "   "   "      "   "   "�  �           �   �   �                                                  �               �     "   "                                                                                                                                                                                                                     �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   �   " � ��      �    �   �   �"  ""  !� �� ��  �               �   " ��.�  ��            "  �"     �                       �".��".  ���    �              �  "� "� "/ "�                         ����                               ���                          ����                  �   �� �       �  �  "�  "   "              �  �                        
���	���̜̽�˽�̈ۻ��ۻ�۽��˲"������"���" ��"                "   "   "                 ���       "   "     ����           �  ��� ݼ� w�� b}� ggp wz�����""H�""T�B"UJ�"UJ�@T�DT�TUJ�  ��.�                           5J� �J� �˻ �˰ ʘ� ̪ ˲"�" ""�"" �  ��                /���"/�  ��                    �                                                                            �               �     "   "                                                                                                                                                                                                                        �   �  �  �  	�  �  EH  ET DU CE DD4 DD3 DC0 �3 ɰ �  ,�  +�  "/  ������ � ̹�p�˚��̹���ː�̼�̻���ۜ��۩�ݍ���=��J�ܰT�� EJ�0 EJ� I�  ��  �"  ""  "/  "�� ���                    ̰ ̻ ̻	���̚�wˢ �+���"����"��"  �   �    �   �" �"� "������     �     �� �� ��
��׊��w٪�|��������            "   "   "       �         �        �   �     �       �       "       .      �                    �"  �""� "�                                                                                                                                                                                                                 �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �   �" �!  �  �� �   �                �  �� Ș ��  ��  �     �!� �                                                                                                                                                                                                                          �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �"  "�  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    ��   �   �"  �""��� �   �      �       �                            ""  "".  . �    �                                                                                                                                       	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��                    ""  ."  �"    "   "   .   .                  �  �  �  �                                          "   "                      �    � �  ��                  ���                     �  � �                       � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                        �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���                            "  ""�����"    /   �  �   ��                                �   �                      �".��".  ���    �                    ".  ".  ���              �  �˰ ��� �wp �&                                                                                                                                                                 �  ��� ݼ� wۺ�b}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  �".�".� ���        T   S   C   3   30  30  ;�  ��  ��� 
�" ��" �""/�"" �����                     �   �                      �".��".  ���    �    �� ���  ��                               �  �˰ ��� �wp �&                                                                                                                                                                                  �� �� �� ��  �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H�� UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �݉  ��  ��  ��� ˙� �˼ ��� �ٚ��ک�����J��J� "D�@�D���4���ˮ軽� ̽� ��� ��ٰ�۰"˰""+�""!��"� �                                                  � � �  (�  .   .   )�  )�  �   �   �   �   �   �   �                      �  .   �� ��     �     �  ��  ��  ��  ��� ��� ��� ��˰ɜ˰��˻�̻���������3���DDD�                                �         �  "� "  �  ��                                                                                                                                       	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��                        �          �   � � /  �"" �"  �    "   "   "  �� ��                   �".��".���                                                                                                                                                                                                                                                       2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq �
*� �FC. �> C4.kj �N kr � �B�1 � B�AB�+ 	B�3 �
B� � �B� � � B� �B� � �B� � �cV � �K( � C> �K7 � K!? �K"2 �K%" � K'! �c�@ � c�HN"� �N "� �>� �>
� ��} ��} �  *&~ � )�v?!� �?"
� � � #*Kv � )�v �%*~ � &*Fv �'*8v �  *Gv � )*Gv �  *Av �  *Av � ,*Fv �-*8v �  *Gv �/*8v �  *Gv �  *AvF 
�D r  *Ou �4
� � {  *Ou ~ 6*Ru ~ *}0 )�tM )�tP )�tA  *Gt2<*8tB  *Gt>*<tD *:t � @"�4 �A�" � 
�1D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� � � � � � � � � � � � � � � � � � � � ����������������������������������������������������<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ���������������������������������������������������� � � � � � � � � � � � � � � � � � � � ���������������������������������������������������� � � � � � � � � � � � � � � � � � � � �����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3�������������������������������������������-�N�X�O�Y�Z�G�T��;�[�[�Z�Z�[� � � � � �-�2�3�����������������������������������������#��<�Z�K�\�K��6�G�X�S�K�X� � � � � � � � �-�2�3�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������,�>�0� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�2�3� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 