GST@�                                                           `}�                                                      � ����     �               ����e ����ʴ������������������        Ti     #    ����                                d8<n    �  ?     �P����  �
fD�
�L���"����D"� j   " B   J  jF�"     "�j  " ���
��
�"    
 �j�
�
  
  ��
  �                                                                               ����������������������������������       ��     bbb  411 c c c           	 
       G � ( (                 nhn 1)         8==�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             �h  )*          == �����������������������������������������������������������������������������                                ��  �       n�   @  #   �   �                                                                                '     1nh)n  )�*h    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE  �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    \�M�VA۞@�[��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�M�VA۞@�[��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�M�VA۞@�[��e3�L(@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8\�M�VA۞@�[��e3�L(@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8�M�VK�۞@�[��e3�L(@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8�M�VK�۞@�[��e3�L(@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8�M�VK�۞@�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/   � �8�M]VK�۞@�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8�M]VK�۞@�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8<�M]VK�۞@�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8<�M]VK�۞@�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8<�M]VK�۞@�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8<�M�VK�۞@�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8<�M�VK�۞@�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8<�M�VK�۞@l�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8<�M�VK�۞@l�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8<�M�VK�۞@l�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8<�M�VK�۞@l�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8<�M�VL۞@l�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8 ��M�VL۞@l�\<�e3�L(@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/   � �8 ��M�VL۞@l�\<�e3�L(@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8 ��M�VL۞@l�\<�e3�L(@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8 ��M�VL۞@l�\<�e3�L(@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8 ��M�VL۞@l�\<�e3�L(@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8L�M�VL۞@l�\<�e3�L(@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8L�M�VL۞@l�\<�e3�L(@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8L�M�VL۞@��\<�e3�L(@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8L�M�VL۞@��\<�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�M�VL۞@��\<�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞@��\L�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞@��\L�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞@��\L�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞@��\L�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞@��\L�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞@��\L�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞@��\L�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞@��\L�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞@��\L�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞A�\<�e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞A�\<�e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞A�\<�e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞A�\<�e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞A�\<�e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞A�\<�e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞A�\<�e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞A�\<�e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞A�\<�e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VL۞A�\��e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞A�\��e3�L(@�@no�\�[Ǽ!۳�T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞A�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞A�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞A�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞A�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞K��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞K��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞K��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞K��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞K��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VL۞K��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VK�۞K��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M=VK�۞K��\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8��MMVK�۞K��\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#;P (%2't ��1"t'! ��/    � �8��MMVK�۞K��\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#;P (%2't ��1"t'! ��/    � �8��MMVK�۞K��\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#;P (%2't ��1"t'! ��/    � �8��MMVA۞K��\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#;P (%2't ��1"t'! ��/    � �8��MMVA۞K��\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#;P (%2't ��1"t'! ��/    � �8��MMVA۞L�\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#KP (%2't ��1"t'! ��/    � �8��MMVA۞L�\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#KP (%2't ��1"t'! ��/    � �8��MMVA۞L�\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#KP (%2't ��1"t'! ��/    � �8��MMVA۞L�\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#KP (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ!���T0 k� ���#KP (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8L�NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�NMVA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8L�NMWA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�NMWA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�NMWA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�NMWA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�NMWA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�NMWA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�NMWA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�NMWA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��NMWA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��N=WA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��N=WA۞L�\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��N=WA۞L�]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��N=WA۞L�]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��N=WA۞L�]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�N=WA۞K��]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�N�WA۞K��]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�N�WA۞K��]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�N�WA۞K��]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�N�WA۞K��]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�N�WA۞K��]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�N�WA۞K��]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�N�WA۞K��]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�N�WA۞A�]��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8�N�WA۞A�]��e3�L(@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8�N�WA۞A�]��e3�L(@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8����X<Q���LM+��#3�L,@˃@n�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8����X<Q���LM'��#3�L(@˃@n�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8����\<Q���LM#��#3�L(@˃@n�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8����\<R��LM��#3�L(@˂@n�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8����`;R��LM� #3�L(@˂@n{�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8����`;R��LM��#3�L(@˂@n{�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8����d;R��LM��$3�L$@ς@n{�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8����d;R��LM��$3�L$@ς@n{�[�[��{��T0 k� ���$P (%2't ��1"t'! ��/    � �8����h:R��LM��$3�L$@ς@n{�[�[��{��T0 k� ���$P (%2't ��1"t'! ��/    � �8����h:R��LM��$3�L$@ς@n{�[�[��{��T0 k� ���$P (%2't ��1"t'! ��/   � �8����l:R��LM��$3�L$@ς@n{�[�[��{��T0 k� ���$P (%2't ��1"t'! ��/    � �8����l:R��L=��$3�L @ς@n{�[�[��{��T0 k� ���$P (%2't ��1"t'! ��/    � �8����l9UK��L=��$3�L @ς@n{�[�[��{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8����p9UK��L<����$3�L @ς@n{�[�[��{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8����p9UK��L<����$3�L @ς@n{�[�[��{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8����t9UK��L<����$3�L @ς@n{�[�[��{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8���t9UK��L<����%3�L@ӂ@n{�[�[��{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8���t8UK��D<����%3�L@ӂ@n{�[�[��{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8���x8UK��D<����%3�L@ӂ@n{�[�[��{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8���x8UK��D<����%3�L@ӂ@n{�[�[��{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8���|8UK��D<����%3�L@ӂ@n{�[�[��{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8���|8A��D<����%3�L@Ӂ@n{�[�[��{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8���|7A��E�����%3�L@Ӂ@nw�[�[��{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8����7A��E�����%3�L@Ӂ@nw�[�[��{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8����7A��E�����%3�L@Ӂ@nw�[�[��{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8����7A��E�����&3�L@Ӂ@nw�[�[��{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8����8A��E�����&3�L@Ӂ@nw�[�[��{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8����8A��E���M|&3�L@ׁ@nw�[�[��{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8����8A��E���Mt'3�L@ׁ@nw�[�[��{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8����8A��E���Mp'3�L@ׁ@nw�[�[��{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8����9A��E���Mh'3�L@ׁ@nw�[�[��{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8����9A��E���Md(3�L@ׁ@nw�[�[��{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8� ��9A��D���M\("��L@ׁ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8���:A��D���MX)"��L@ׁ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8���:A��D���MP)"��L@ׁ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8� ͐;A��D���ML*"��L@ׁ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8� ͐<A��D���MD*"��L@ׁ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�$͐<A��D���=@+"��L@ׁ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�$͔=A��D���=8+"��L@ׁ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�$͔>A��D���=4,"��L@ׁ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�$͔>A��D���=0-"��L@ׁ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�$	��?A��D���=(-"��L@ہ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�(
��@A��D���=$."��L@ہ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�(��AA��D���=/3�L@ہ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�(��AA��D���=03�L@ہ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�(��BA��D���=13�L@ہ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�(͐CA��D���=23�L@ہ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�(͐DA��D���M33�L@ہ@nw�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�(͐EA��D���M43�L@ہ@ns�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�$͐FA��D���M 53�L@ہ@ns�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�$͌FA��D���L�63�L@ۀ@ns�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�$݌GA��D���L�73�L@ہ@ns�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�$݈HA��D���<�83�L@ہ@ns�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8� ݈IA��D���<�93�L@ہ@ns�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8� ݄JA��D���<�:"s�L@ہ@ns�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8� ݄JA��D���<�;"s�L@ۂ@ns�[�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��KA��D��<�="s�L@ۂ@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��|LA��D��<�>"s�L@߂@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8� �|MA��E�{�<�?"s�L@߂@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�!�xMA��E�{�<�A"s�L@߃@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�#�xNA��E�t,�B"s�L@߃@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�$tOA��E�p,�C"s�L@߃@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�&pOA��E�p,�E"s�L@߃@ns�[��[��{��T0 k� ���$P (%2't ��1"t'! ��/    � �8�'pPA��E�l,�F"s�L@߄@ns�[��[��{��T0 k� ���$P (%2't ��1"t'! ��/    � �8�)lQA��E�l,�G"s�L@߄@ns�[��[��{��T0 k� ���$P (%2't ��1"t'! ��/    � �8�+lQA��E�h	,�I3�L@߄@ns�[��[��{��T0 k� ���$P (%2't ��1"t'! ��/    � �8�,hRA��Fh,�J3�L@߄@ns�[��[��{��T0 k� ���$P (%2't ��1"t'! ��/    � �8� .hSA��Fh,�L3�L@߄@ns�[��[��{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8��0dSA��Fd,�M3�L@߅@ns�[��[��{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8��1`TA��Fd,�O3�L@߅@ns�[��[��{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8��3`TA��Fd,�P3�L@߅@ns�[��[��{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8��5-\UA��F`,�R3�L@߅@ns�[��[��{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8��6-\VA��F`,�S3�L@߅@ns�[��[��{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8��8-XVAáF`�U3�L@߅@ns�[��[��{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8��:-XWAáF`�V3�L@߆@ns�[��[��{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8��<-TWAáF`�W3�L@߆@ns�[��[��{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8��=-TXAáD�`�Y3�L@߆@ns�[��[��{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8��?-PXAáD�`�Z3�L @߆@ns�[��[��{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��A-PYAáD�`!��\3�L @�@ns�[��[��{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��C-PYAáD�`#��]3�L @�@ns�[��[��{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��E-LZAáD�`%��^3�L @�@ns�[��[��{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��F-LZAáD�`'��`3�L @�@ns�[��[��{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��H-H[AáD�d)��a3�L @�@ns�[��[��{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8��I-H[AàD�d+��b3�L @�@ns�[��[��{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8ݸK-D\AǠD�d,��c3�L @�@ns�[��[��{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8ݴM-D\AǠD�d.��e3�L @�@ns�[��[��{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8ݰN-D]AǠD�h0��f3�L @�@ns�[��[��{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8ݨP-@]AǠD�h2��g3�L @�@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�Q-@^AǠL|h4��h3�L @�@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�S-<^AǠL|l6��i3�L @�@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�T-<_AǠL|l8��j3�L @�@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�V-<_AǠL|l:��l3�L @�@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�W-8`AǠL|p<��m3�L @�@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8݄Y-8`AǠL|p=��n3�L @�@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�|Z-8`AǠL|p?��o3�L @�@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�|Z-0aAǠL|tA��p3�K�@�@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�x[-,bAǠL|tC��q3�K�@�@ns�[��[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�t\-(bAǠL|tD��r3�K�@�@ns�\�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�p]-$cAˠL|xF��s3�K�@�@ns�\�[��{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�l^- dAˠL|xH��t3�K�@�@ns�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�h_-dAˠL|xI��u3�K�@�@ns�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�d`-eAˠL||K��v3�K�@�@ns�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�`a-eAˠL�|L��w3�K�@�@ns�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�Xb-fAˠL�|N��x3�K�@�@ns�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�Tc-gA˟L�|O��y3�K�@�@ns�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�Pd-gA˟L��Q�z3�K�@�@ns�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8�Ld-hA˟L��R�z3�K�@�@ns�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8�Ld- hA˟L��T�{3�K�@�@ns�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8�He,�iA˟L��U�|3�K�@�@no�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8�De,�iA˟L��W�}3�K�@�@no�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8�@f,�jA˟L��X��~3�K�@�@no�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8�<f,�jA˟L��Y��~3�K�@�@no�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8=8f�kA˟L��[��3�K�
@�@no�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8=0g�lA˟L��\���3�K�
@�@no�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8=,g�lAϟL��]���3�K�
@�@no�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8=(g�mAϟL��^��3�K�
@�@no�\�[ü!���T0 k� ���#�P (%2't ��1"t'! ��/    � �8=$g�mAϟL��`��3�K�
@�@no�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�g�nAϟL��a��3�K�
@�@no�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�g��nAϟL��b��~3�K�
@�@no�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�g��oAϟL��c��~3�K�
@�@no�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�g��oAϟL��e|�}3�K�
@�@no�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8�g��oAϟL��f|�}3�K�
@�@no�\�[ü{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8� g��oK�ϟL��g|�}3�K�
@�@no�\�[ü{��T0 k� ���#;P (%2't ��1"t'! ��/   � �8� g��oK�ϟL��h|�}3�K�
@�@no�\�[ü{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8� g�oK�ϟL��h|�}3�K�
@�@no�\�[ü{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8��f�oK�ϟL��i��}3�K�
@�@no�\�[ü{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8��f�oK�ϟL��j��}3�K�@�@no�\�[ü{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8��e�oK�ϟL��j��}3�K�@�@no�\�[ü!˯�T0 k� ���#KP (%2't ��1"t'! ��/    � �8��e�oK�ϟL��k��}3�K�@�@no�\�[ü!˯�T0 k� ���#KP (%2't ��1"t'! ��/    � �8��e�oK�ϟL��l��}3�K�@�@no�\�[ü!˯�T0 k� ���#KP (%2't ��1"t'! ��/    � �8\�d�oK�ϟL��l��}3�L @�@no�\�[ü!˯�T0 k� ���#KP (%2't ��1"t'! ��/    � �8\�d�oK�ϟL��m��}3�L @�@no�\�[ü!˯�T0 k� ���#KP (%2't ��1"t'! ��/   � �8\�c�oK�ϟL��n��}3�L @�@no�\�[ü!˯�T0 k� ���#[P (%2't ��1"t'! ��/    � �8\�c�oK�ϟL��n��}3�L @�@no�\�[ü!˯�T0 k� ���#[P (%2't ��1"t'! ��/    � �8\�c�oK�ϟL�|o��}3�L @�@no�\�[ü!˯�T0 k� ���#[P (%2't ��1"t'! ��/    � �8\�b�oK�ӟL�|o��}3�L @�@no�\�[ü!˯�T0 k� ���#[P (%2't ��1"t'! ��/   � �8\�b�oLӟL�|o��}3�L@�@no�\�[ü!˯�T0 k� ���#[P (%2't ��1"t'! ��/    � �8\�a�oLӟL�xo��}3�L@�@no�\�[ü!˯�T0 k� ���#kP (%2't ��1"t'! ��/    � �8\�a,�oLӟL�xo��}3�L@�@no�\�[ü{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8\�a,�oLӞL�to��}3�L@�@no�\�[ü{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8\�`,�oLӞL�to��}3�L@�@no�\�[ü{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8l�`,�oLӞL�po��}3�L@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8l�`,�oLӞL�poܜ}3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�_,�oLӞL|lpܜ}3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�_,�oLӞL|lpܜ}3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�_,�oLӞL|hpܜ}3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�^,�oLӞL|hpܠ}3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�^,�oLӞL|hpܠ}3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�^,�oLӞL|dpܠ}3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�],�nLӞD�dqܠ|3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�],�nLӞD�dqܠ|3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�],�nLӞD�`q|�|3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�],�nLӞD�`r|�|3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8l�\,�nLӞD�`r|�|3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�\,�nLӞF`r|�|3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�\,�mLӞF`s|�|3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�\,�mLӞF`s|�{3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�[,�mLӞF`t|�{3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�[,�mLӞF`t|�{3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�[,�lLӞE�`u|�{3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�Z,�lLӞE�`u|�z3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�Z,�lLӞE�`v��z3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�Z,�kLӞE�`v��y3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�Z,�kLӞE�`v��y3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�Y,�kLמE�dw��y3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�Y,�jLמE�dw��y3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�Y,�jLמE�dw�x3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�Y,�iLמE�dw�w3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�Y,�iLמE�dw�w3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�X,�iLמE�dw�w3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�X,�hLמE�dw�w3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�X,�hLמE�dw�v3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�X,�gLמE�dw�v3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�X,�gLמB�hwܨu3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8l�W,�fLמB�hwܬt3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�W,�fLמB�lwܬt3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�W,�eLמB�lwܬs3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8l�W,�eK�מB�lwܰr3�L@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8l�W,�dK�מB�lw|�q3�L@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8l�V�dK�מB�pw|�q3�L@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8l�V�cK�מB�pv|�q3�L@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8l�V�cK�מB�pv|�p3�L@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8\�V�bK�מB�pu|�o3�L@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8\�V�bAמB�tu\�o3�L@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8\�U�aAמB�tt\�n3�L@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8\�U��aAמCxt\�m3�L@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8\�U��`AמCxs\�m3�L@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8\�U��`AמC|s\�m3�L@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��U��_K�מC|s\�l3�L@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��T��^K�מC|r\�l3�L@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��T��^K�מC|r\�k3�L@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��T��]K�מC|q\�j3�L@�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8��S��]K�מC�pl�j3�L@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8��S��]K�מC�pl�j3�L@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8��R��\K�מC�pl�j3�L@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8��R��\K�מC�ol�j3�L@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8��Q��[K�מC�ol�j3�L@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8��Q��[K�מC�nl�j3�L@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8�P��ZK�מC�ml�i3�L@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8�O��ZLמC�ml�i3�L@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8�O��ZLמC�ll�i3�L@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8�N��YLמE�k\�h3�L@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8�M��YLמE�j\�h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M��YLמE�j\�h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��L��YLמE�j\�h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��K��YL۞E�i\�h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��K��XL۞E�i\�h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��J��XL۞E�i\�h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��J�XL۞E�i\�h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��I�XL۞E�i\�h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��I�XL۞E�h��h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��I�XL۞B��h��h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H�WL۞B��g��h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H�WL۞B��g��h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H�WL۞B��f��h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H�WL۞B��f��h3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H�WL۞B��e��g3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H\�WL۞B��e��g3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H\�WL۞B��e��g3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H\�WL۞B��e��g3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H\�WL۞B��d��g3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H\�WL۞B��d��g3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��H\�WL۞B��d��g3�L@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�H\�WL۞B��d��g3�L @�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�H\�WL۞B��d��g3�L @�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�H\�WL۞B��d��g3�L @�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�H\�WL۞B��d��g3�L @�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�H\�WL۞B��d��g3�L @�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�H\�WL۞B��d��g3�L @�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�H\�WL۞B��d��g3�L @�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�H\�WL۞B��c��g3�L @�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�H�WL۞B��c��g3�L @�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�H�WL۞B��c��g3�L @�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8L�H�WL۞K��c��g3�L @�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8L�H�WL۞K��b��g3�L @�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8\�H�WL۞K��b��g3�L @�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8\�H�WL۞K��b��g3�L @�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8\�H�WL۞K��b��g3�L @�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8\�H�WL۞K��a��g3�L @�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8\�H�WL۞K��a��g3�L @�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8\�H�WK�۞K��a��g3�L @�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8\�H�WK�۞K��a��g3�L @�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8\�H�WK�۞K��`��g3�L @�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8\�H�WK�۞K��`��g3�L @�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8\�H�WK�۞K��`��g3�L @�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8\�H,�WK�۞K��`��g3�L @�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8l�H,�WA۞K��_��g"s�L @�@no�\�[Ǽ{��T0 k� ���#[P (%2't ��1"t'! ��/    � �8l�H,�WA۞K̨_��g"s�L @�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8l�H,�WA۞K̨_��g"s�L @�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8l�H,�WA۞K̨_��g"s�L @�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8l�H,�WA۞K̨_��g"s�L$@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8l�H,�WA۞K̨^��g"s�L$@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8l�H,�WA۞K̨^��g"s�L$@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8l�H,�WA۞K̬^��g"s�L$@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8l�H,�WA۞K̬^��g"s�L$@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! �/    � �8l�I,�WA۞K̬]��g"s�L$@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8l�I,�WA۞K̬]��g"s�L$@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8|�I,�WA۞K̬]��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8|�I,�WA۞K̬]��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8|�I,�WA۞K̬]��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8|�I,�WA۞K̬]��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8|�J,�WA۞K̬\��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8|�J- WA۞K̬\��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8|�J- XA۞K̰\��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8|�J- XA۞K̰\��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8|�J- XA۞K̰\��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��J-XA۞K̰\��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��J-XA۞K̰[��g3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��J-XA۞K̰[��g"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��J-XA۞K̰[��g"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8 ��J-XA۞K̰[��f"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�K-XA۞K̰[��f"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�K-XA۞K̰[��f"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�K-XA۞K̰Z��f"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�L-XA۞K̴Z��f"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�L-XA۞K̴Z��f"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�L-XA۞K̴Z��f"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8L�L-XA۞K̰Z��e"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8L�L-XA۞K̰[��e"��L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/   � �8\�M-XA۞K̰[��e3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�M-XA۞K̰[��e3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�M-XA۞K̰[��e3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�M-XA۞K̰[��e3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�M-XA۞K̰[��d3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�N-XA۞K̰[��d3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�N-XA۞K̬[��d3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�NXA۞K̬[��d3�L$@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�NXA۞K̬[��d3�L$@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8 ��NXA۞K��[��d3�L$@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8 ��NXA۞K��[��d3�L(@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/   � �8 ��NXA۞K��[��d3�L(@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8 ��NXA۞K��[��d3�L(@�@no�\�[Ǽ{��T0 k� ���$P (%2't ��1"t'! ��/    � �8 ��N�XA۞K��[��d3�L(@�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8�N�WA۞K��[\�d3�L(@�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8�N�WA۞@�[\�d3�L(@�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8�N�WA۞@�[\�d3�L(@�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8�N�WA۞@�\\�d3�L(@�@no�\�[Ǽ{��T0 k� ���#;P (%2't ��1"t'! ��/    � �8�N�WA۞@�\\�d3�L(@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8�N�WA۞@�\\�d3�L(@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8�N�WA۞B��\\�d3�L(@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8�N�WA۞B��\\�d3�L(@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8�N�WA۞B��\l�d3�L(@�@no�\�[Ǽ{��T0 k� ���#KP (%2't ��1"t'! ��/    � �8�N�WA۞B��\l�d3�L(@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8\�N�WA۞B��\l�d3�L(@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8\�N�WA۞B��\l�d3�L(@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8\�N�WA۞B��\l�e3�L(@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8\�N�WA۞B��\l�e3�L(@�@no�\�[Ǽ{��T0 k� ���#kP (%2't ��1"t'! ��/    � �8\�N�WA۞B��\l�e3�L(@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8\�N�WA۞B��\l�e3�L(@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8\�N�WA۞B��\l�e3�L(@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8\�N�WA۞B��\\�e3�L(@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8\�N�WA۞B��\\�e3�L(@�@no�\�[Ǽ{��T0 k� ���#{P (%2't ��1"t'! ��/    � �8\�N�WA۞B��\\�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�N�WA۞B��\\�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�N�WA۞@�\\�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N]WA۞@�\\�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N]WA۞@�\\�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N]WA۞@�\\�e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N]WA۞@�\\�f3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N]WA۞B��\��f3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N�WA۞B��\��f3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N�WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N�WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N�WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N�WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N�WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N�WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N�WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��N]WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M]WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M]WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M]WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M]WA۞B��\��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�WA۞B��[��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�WA۞B��[��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�WA۞B��[��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�WA۞B��[��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�WA۞@�[��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8��M�VA۞@�[��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8\�M�VA۞@�[��e3�L(@�@no�\�[Ǽ{��T0 k� ���#�P (%2't ��1"t'! ��/    � �8                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��,� ]��� �  NO�        ��6G�     NO��6G�                       	 Z�8�         �      ��    8(          W�   > > 
    ��E`q     W��E�     j��               2 Z�8         �`�     ��    @
	"         ��c    	    ���`    ��c���`           	             Z�8         ��     ��   		'           ]n�    	    �-�.     ]n��-�.                        	 Z�8          �     ��   8
           e�     
    .�<�f     e��<�f                       	 Z�8          �`     ��    X

          
j  ��     B ���     
j ���                               ���              <  ��     0 0             \�  $ $       V�
Ә     \��
Ә                          B��          �0     ���   8

�         ��~          j���f    ��~���f                       	 A��           �     ���   0	 	          ��Y�         ~���    ��Y����                         ����          f�     ���   (	"	          ����         ����    �������                           �$         	 J�     ���   H	w         ���          ���    �����                           �$         
 6�     ���   (
         �ܟs ��	      ����    �ܟs���                            �� a               �  ���    0

 2                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         ��s  ��        ���~E    ��s��~E         "                 x                j  �   �   �                             � @@       ���   �r    ��   �X     z                                      .         �                         �6�E���-�< ��
��������������� 	    
             
 �   .�� 5K�B       ��  }` ��  }� �� 0d` �D  d� �� e  � �[� �  \� �D g  �d g  V� g@ �� 0g  �$ g` �D g� 
�\ V  
�\ V  
�| W� 
�\ W� 
�\ W� H� d� 
�| W� 
�\ V� 
�� V� 
�\ W  
�\ W� 
�\ W� 
�\ W� �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� � }`���� � � }`���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����8�� �� �  ������  
�fD
��L���"����D" � j  "  B   J jF�"     "�j  " ��
��
��"     
�j
�� 
  
 �
� �  �  
� ��   ��     ���  �   ��    ��     ���      ����  ��     ���          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �/  '      �� �2 ��        �4 �  ���        �        ��        �        ��        �     �     ��������        ��                         T�) , %	 �                                    �                ����            ������#�%� �    �8 (               22 Dino Ciccarelli     5:33                                                                       1   2     �&
*� �=�� �1�� � c� �) c� �"c� �"c� �B c� �	� �
� �K ~2K n1 � �c� �0 c� �cV � c^ � �K= �K"- �B�. �B�> �C.H � C6@ �B�7 � B�G uk~ z �k� j Ukj q="� z= "� �-"� v- *� �B!"� �B ""� �2#� �2$
� �@  *Kh2&� �2'
� �@  *Kh2)� �2*
� �@  *GhP  *RxX -*K`P  *RxX  *H`X  *H`X  *K`X  *K`X  *K`X  *K`X  *K`8 6*DpP 7*RxX 8*K�X  *K`X  *K`$;*:wD  *AwZ  *AtU  *K �  "P y# 
� �                                                                                                                                                                                                                 �� R   �               $� �     I P E h  ��        
            �������������������������������������� ���������	�
��������                                                                                          ��    �Z�   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E �X 7�  	� �@Y��3����A��                                                                                                                                                                                                                                                                                                                                           @�                                                                                                                                                                                                                                                    T    9 "   ��  4�J      W�  	                           ������������������������������������������������������                                                                                                                                          �  ��              �          ��               	 
     �������� ���� ������������������ ������������� �������� ������������ ��������������������� ����������� � ������������ ������ � �  ������������� ������ ���������������� ��������������������� ���������� ������� �� ����������� �� ������������       	    x                   s     %     ��  .�J      H                             ������������������������������������������������������                                                                                                                                          �  ��                �        P    �          	     ��  ����������   ���� �� ����� ��������������������� ������ ���� ��� ��� ������ �����������������������������  ���� ��������� �������� ������������   ����������������  ������� ������ �������� ��������� ��                                                                                                                                                                                                                                                                                             	          
                   �             


             �  }�                     '�                                          '�                        ��������      	��������������������������������    ����������������������������  '�����  's������������""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" ) J >                                 � �l� �}`                                                                                                                                                                                                                                                                                    1nh)n  )�*h        m      m            k            d      e      m                                                                                                                                                                                                                                                                                                                                                                                                           J �  /#�  >#�  C#�  G#�  EZm< �̎����
����&������I�̞�&�����4 �N x�����        .  �`�? :����          �   & AG� �   "   
              �                                                                                                                                                                                                                                                                                                                                      p N K   �                "         !��                                                                                                                                                                                                                        Y   �� �~ �       �� 8      �������� ���� ������������������ ������������� �������� ������������ ��������������������� ����������� � ������������ ������ � �  ������������� ������ ���������������� ��������������������� ���������� ������� �� ����������� �� ��������������  ����������   ���� �� ����� ��������������������� ������ ���� ��� ��� ������ �����������������������������  ���� ��������� �������� ������������   ����������������  ������� ������ �������� ��������� ��             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    J       8   � ��                       8     �  �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �f ��     �f �$ ^$ �@       �       �     �   n 
� �     �f ��        p���o� H� �    � �$ ^$    ��   0  ��      �   �   ��Ӕ����������J����  ~����    ���     �H   �z � �N ^$         �>         �c   }` �� �� }` �� �$  �8  �� � 8      �       ���� e�����   g��� 	 �     f ^�        ��              ��-,���2�������J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                          �      �  a r!   f�"""""*��**"*�"�""�""v""*f   "  ""- ��"�"*"-""z"""""����            n   �  "  q  ��                          �  �                                 � gv"!g�vg�vggfvv|�b��r""gb"�vr�rgb��v���g���v���***�*q!q�"!a�!vwfqqr~� qw��q�~~q�����~~~�w~~w�w            �   ~   ��  ~~  �w      v    �                ggj�vvggvvgg!vg�g֪vvg�r�r��⢪rq**gjb�v�q*gjj*vv��gg�z�/�"!�"�*�""*z����qw�~q~ww��q~qwvq�w�`� ��� �w �~p w�p  ��                    �                        lggz�v��g        �       ggbvvrgggavvvqggav� �      ���w!z�w"""�!""*�"! ��        q� q�        `               �        �                      wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����   �   �   �   ����                                     	�  		  	 � 	 	 	   	   	   	   	  ��                  ��   	   	   	   	   	   	 	 	 � 		  	�                 �   	    �   	    �   	    �   	   	   �  	   �  	   �  	   �                                      
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  " ! " ""  "!  "" "  """                                                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """"! "   "      ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       """ "!   " ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                      �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �      �                                                                            �               �  �  ��  �   �   �           �     �                                                                                                                                                                                     � 
��	�˽���w��{k��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            �  �  �  ��  �           "! � ����                              � �� ��� ��        �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                  �       �                        �   ��  ���  � �    �                                                                                                                                                     �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �                           � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                    �   ���                            �   �                                                                                                                 �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �                           � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                                                                                                                                                                 �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    4U� 4U� 4U� 3UXP�EX��U����  ��                    �  ��� ݼ� �    �    �   �                     �  �  �   �   �   �                   �   �               �  ��� ݼ� w{� �װ vw�                                                                                                                                                                                         �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                     �� ̽ ̽ ۽ }�  �� 
�� ��� ��� ��� ˼� ��� ��� 	ۉ �8 ��X�� �D �C �3 �0 ��  ��� ˻ �,� ""�"" �  �                        ��  ��  �̰ �˻ �̻���˰�ͻ���� ��� �Ș ��3 ��3 333 D33 330 330 ��� ��� ̰ �� "/   ���  � �� ��           �   ��  � � ��      �    �      �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                                                                                                                                                                                                                                  �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   �   �   �   ˰  ˙  ɪ  ��� ټ� �̰ �̰ ��� ��  ��                              ��          �   �       �    �                     �   �  �  �                �   ��  �   ��  ��  �  �  �   �                   � �������������  �                                                                                                                                                              	   �  �  �� �� ��� �����ɘ�̻9�̼3�̌39��U33=U3: �ET �4E��4ʠ "�" """""������ ���                        �� �� ��� ��� ��w ��p ˚� ̹� �˰ ��� ��  ��  ��  ̻" ��".�2" ��" T�  E�0 4�0���O�  �� ,�  ""/ "!�� ����           �� ����  �       �   �   �                                                   ��                  �                        ���� ��� ����                            ��  ��  ���                                                                                                                                                                                                  	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                       �  ��  ��  ww  ��  vv  w                   �   �                      �������  ���    �                    ��  ��  ���                                                                                                                                                                                                  	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                                                                                                                                                                                                                                               �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �   �"!�����                            �  �� Ș ��  ��  �                                                                                                                                                                                                                                                 �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@  �D�JJN�J��J��J��J��JJD�N�                    �   �          �     	 ��̠       �  �   
�  �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                             "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""����������D��M��M""""����������""""�����ADMA����""""����DD�M�""""��������AD�DM�""""�����������A�A�""""������AD�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��M��M�������D����3333DDDD�DD�M�D�������3333DDDDD�������M�DM�D����3333DDDD��A�M�M���M�����3333DDDDMM������D��D����3333DDDDA�A�A�D��M�D�����3333DDDD�������������D������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�""""��������AA�A �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�ADA�LL��L�D����3333DDDD = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=LL����������D����3333DDDD    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"����������A������ x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx""""�������I�I������ w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww""""�������I��D���I�������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(�D�M�D���M������3333DDDD �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((�D�M�A�����MD�����3333DDDD ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""�����AMAD������ M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M""""������������������ � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�fFfFDfFFfFffdFffff3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DDFFDfFFfdFffff3333DDDD 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5""""wwwwwwwGGD x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x""""wwwwwwqwAqwAwA w w x y�������H���������������������������������H������yxww""""wwwwqwqAwAqAqAq  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(A�A�A�A��LD�����3333DDDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,�A�LDL�L�D�L�����3333DDDD +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+""""wwwwwwDGAD 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5""""wwwwqqDAAq =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=""""wwwwwwwGGwGGwGwGw     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( UQUUQUUQUUQUUUDUUUUU3333DDDD � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � �DEQQUUDUTEUUUU3333DDDD � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � �""""������������������������ ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""�������DAADAI M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M�A�AM�M�DM��M334CDDDD � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�DD����M��DM�����3333DDDD � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�""""wwwwwwDGqGq 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5""""wwwwwwwGwwDGwwwwwwww x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xADAH�DJ�H�H�����3333DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww�H��J�AD�DH�D����3333DDDD + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""�������DD����� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq&
*� �=�� �1�� � c� �) c� �"c� �"c� �B c� �	� �
� �K ~2K n1 � �c� �0 c� �cV � c^ � �K= �K"- �B�. �B�> �C.H � C6@ �B�7 � B�G uk~ z �k� j Ukj q="� z= "� �-"� v- *� �B!"� �B ""� �2#� �2$
� �@  *Kh2&� �2'
� �@  *Kh2)� �2*
� �@  *GhP  *RxX -*K`P  *RxX  *H`X  *H`X  *K`X  *K`X  *K`X  *K`X  *K`8 6*DpP 7*RxX 8*K�X  *K`X  *K`$;*:wD  *AwZ  *AtU  *K �  "P y3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������������������������� �!����� � � �m�n�|�}�c�d�v�w��� � � � � ��������������������������������������"�#�j�k�&�'�(����� � � ������������������ � � � � ��������������������������������������)�*�l�m�n�.�/������#��6�G�X�S�K�X��a��b� � � � ��������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������#��<�Z�K�\�K��6�G�X�S�K�X� � � � � � � � �-�2�3�����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3�������������������������������������������.�O�T�U��-�O�I�I�G�X�K�R�R�O� � � � � �.�/�=����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������=��#�%� � ������������������.�/�=� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�2�3� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            