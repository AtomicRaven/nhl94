GST@�                                                            \     �                                               � ���      �  �           �������J 
 J�������������������        �g      #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"     "�j  " ���
��
�"    
 �j�
�
  
  ��
  F�                                                                              ����������������������������������       ��    =b 0Qb 4 114  4c  c  c      	 
      	   
       ��G �� � ( �(                 �nn 	)1         88�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             F�  ))          == �����������������������������������������������������������������������������                                $�  �   H  ��   @  #   �   �                                                                                '    	�)n1n  )F)�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y�DO  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    ���П�E�c�B�#����|,�c�D�DЧ�cS��P3��T0 k� �C��G�(%2't ��1"t'!  ��" 
   ��� ����Ч�E�c�B�+����|,�k�D��DЧ�cS��P3��T0 k� �C��G�(%2't ��1"t'!  ��" 
   ��� �������E�c�B�3����|,�s�D��DЫ�cW��P
3��T0 k� �O��S�(%2't ��1"t'!  ��" 
   ��� �������E�c�EC����|,���D��Dг�cW��T
3��T0 k� �W��[�(%2't ��1"t'!  ��" 
   ��� �������E�_�EG����|,���D��Dෙc[��T
3��T0 k� �_��c�(%2't ��1"t'!  ��" 
   ��� �������E�_�EO����|,�D��D໘c[��T
3��T0 k� �c��g�(%2't ��1"t'!  ��" 
   ��� �������E�_�EW����|,�D��D࿘S[��T
3��T0 k� �g��k�(%2't ��1"t'!  ��" 	   ��� �������E�_�E_��÷|,�D�D�ØS[��T	3��T0 k� �k��o�(%2't ��1"t'!  ��" 	   ��� �������E�_�Eg��˶|,�D�D�ǙS[��T	3��T0 k� �k��o�(%2't ��1"t'!  ��" 	   ��� ������E�[�Eo��Ӷ|,�D�D�˙S[��T	3��T0 k� �k��o�(%2't ��1"t'!  ��" 	   ��� ������E�[�Ew��۵|,�ÕD� D�ϙS[��T	3��T0 k� �k��o�(%2't ��1"t'!  ��" 	   ��� �����E�[�E{���|,�˖D�,D�әS[��T	3��T0 k� �k��o�(%2't ��1"t'!  ��" 	   ��� �����E�[�E�����|,�ۗD�<D�ߚS[�CT	3��T0 k� �g��k�(%2't ��1"t'!  ��" 	   ��� ��'��#�F[�E������|,��D�HD��SW�CT	3��T0 k� �o��s�(%2't ��1"t'!  ��" 	   ��� ��/��+�F[�E�����|,��D�PD��SW�CT	3��T0 k� �w��{�(%2't ��1"t'!  ��" 	   ��� ��3��3�F[�E�����|,��D�XD��SW�CT	3��T0 k� �{���(%2't ��1"t'!  ��" 	   ��� ��7��;�F_�E�����|,���D�dD��CS�CT	3��T0 k� ������(%2't ��1"t'!  ��" 	   ��� ��;��C�F_�Dݳ���|,��D�lD���CS�CT	3��T0 k� ������(%2't ��1"t'!  ��" 	   ��� ��?��K�Fc�Dݻ��#�|,��D�t D���CO�CT	3��T0 k� ������(%2't ��1"t'!  ��" 	   ��� ��C��W�Fg�D�Ó�+�|,��E| D��CO�CT	3��T0 k� ������(%2't ��1"t'!  ��" 	   ��� ��C��_�Fo�D�˓�3�|,��E�!D��CK��T	3��T0 k� ������(%2't ��1"t'!  ��" 	   ��� ��K��o�Fw�D�ߒ�C�|,�/�E�"D��CG��T	3��T0 k� ������(%2't ��1"t'!  ��" 	   ��� ��K��w�F{�D���K�|,�7�E�#D��CC��T	3��T0 k� ������(%2't ��1"t'!  ��" 	   ��� ��O���F�D���S�|,�?�E��#D��C?��T	3��T0 k� ������(%2't ��1"t'!  ��" 	   ��� ��O����F��D����[�|,�G�E��$E'�C;�3T	3��T0 k� ������(%2't ��1"t'!  ��" 	   ��� ��S����F��D����c�|,�O�E��%E+�C;�3T	3��T0 k� ������(%2't ��1"t'!  ��"    ��� ��T���F��D���s�|,�[�E��&E7�C3~3T	3��T0 k� ����(%2't ��1"t'!  ��"    ��� ��T���F��D���{�|,Bc�E��'E?�C/~3T	3��T0 k� ����(%2't ��1"t'!  ��"    ��� ��T���E���D�#�΃�|,Bk�E��'E�G�C+T	3��T0 k� �� �� (%2't ��1"t'!  ��"    ��� ��T���E���D�+�ދ�|,Bs�E��(E�K�C'T	3��T0 k� ������(%2't ��1"t'!  ��"    ��� ��T���E���D�3�ޓ�|,Bw�E��)E�S�3#�T	3��T0 k� ������(%2't ��1"t'!  ��"    ��� ��T	���E���D�C�ޣ�|,���E�*E�c�3�T	"��T0 k� �� �� (%2't ��1"t'!  ��"    ��� ��T
���E���D�O�ޫ�|,���Er+E�g�3�
�T	"��T0 k� �� �� (%2't ��1"t'!  ��"    ��� ��T���E�� D�W�޳�|,���Er,E�o�3�
�X	"��T0 k� ����(%2't ��1"t'!  ��"    ��� �	�T���E��D�_�޻�|,���Er-E�w�C�
�X	"��T0 k� ����(%2't ��1"t'!  ��"    ��� �	�T���E��D�g��é|,���Er(.E��C�
�X	"��T0 k� ����(%2't ��1"t'!  ��"    ��� �	�T��E��D�{��Ө|,���Er81Eq��C�
�\	"��T0 k� ����(%2't ��1"t'!  ��"    ��� �	�T��E��D����ۨ|,���Er@2Eq��C�
�`	"��T0 k� ��� (%2't ��1"t'!  ��"    ��� �	�T��E��	D�����|,���ErH3Eq��B��
�`	"��T0 k� ��(%2't ��1"t'!  ��"    ��� �	�T�'�E��D�����|,���ErP5Eq��B���`	"��T0 k� ��(%2't ��1"t'!  ��"    ��� �	�T�/�E��D�����|,�ǻD�X6Eq��B���`	3�T0 k� ��(%2't ��1"t'!  ��"    ��� �	�T�?�E�D�����|,�ϾD�d9Eq��B��`	3�	T0 k� � �$(%2't ��1"t'!  ��"    ��� �	�T�G�E�E����|,���D�l:Eq��R��`	3�
T0 k� �(�,(%2't ��1"t'!  ��"    ��� �	�T�S�F�E����|,���D�t;EqûR��d	3�
T0 k� �4�8(%2't ��1"t'!  ��"    ��� �	�T�[�F�EǓ��|,���I�|=EqǼR��d	3�T0 k� �@�D(%2't ��1"t'!  ��"    ��� �	�T�k�F�,Eה�+�!�,���I҈?D�ӿR��d3�T0 k� �P�T(%2't ��1"t'!  ��"    ��� �	�T�s�F�4Eߔ�3�!�,���IҌ@D���Rߓ�d3�T0 k� �X�\(%2't ��1"t'!  ��"    ��� �	�T�{�F�8E��;�!�,���IҔAD���R۔h3�T0 k� �d�h(%2't ��1"t'!  �"    ��� �	�T҃�F�@E��C�!�,���I�BD���Rەh3�T0 k� �l�p(%2't ��1"t'! ��/    ��� �	�Tҗ�F�LE��S�!�,���I�DD���Rәh"s�T0 k� ����(%2't ��1"t'! $�/    ��� �	�T���F�TE��[�!�,���I�ED���RϚh"s�T0 k� 3�����(%2't ��1"t'! ��*    ��� �	�T���F�\D���c�!�,���I�FD���bϜ�l"s�T0 k� 3�����(%2't ��1"t'! ��*    ��� �	�T���F�`D���o�!�,���Er�GD��b˞�l"s�T0 k� 3�����(%2't ��1"t'! ��*    ��� �	�T���F�pD�+���!�,��Er�ID��bǡ�l"s�T0 k� 3�����(%2't ��1"t'! ��*    ��� �	�T���F�tD�3����|,�Er�JD��bã�p"s�T0 k� ������(%2't ��1"t'! �*    ��� �	�T���F�|E�;����|,�Er�KD��b���p"s�T0 k� ������(%2't ��1"t'! ��*    ��� �	�T���F�� E�C����|,�Er�LD��b���t "s�T0 k� ������(%2't ��1"t'!  ��*    ��� �	�P���F��!E�O����|,�Er�MD�#�b��sw�"s�T0 k� ������(%2't ��1"t'!  ��*    ��� �	�P ��F��"E�O����|,+�Er�PD�+�b��s{�3�T0 k� #�����(%2't ��1"t'!  ��*    ��� �P ��F��#E�W����|,/�Er�QEr/�b��s{�3�T0 k� #�����(%2't ��1"t'!  /�*    ��� �P!��F��$E�_����|,7�Er�REr7�2��s�3�T0 k� #�����(%2't ��1"t'!  ��*    ��� �P!��F��%E�c��Ǡ|,#;�Er�TEr;�2��s�3�T0 k� #�����(%2't ��1"t'!  ��*    ��� �L"��F��'E�s��ן|,#G�Er�WErC�2��s��c�T0 k� C�����(%2't ��1"t'!  ��*    ��� �2L#��F��'E{��ߟ!�,#O�Eb�XErG�2��s��c�
T0 k� C�����(%2't ��1"t'!  ��*    ��� �2L#�F��(E����!�,#S�Eb�ZErK�2��s��c�
T0 k� C�����(%2't ��1"t'!  ��*    ��� �2L$�E��)E����!�,#S�Eb�[ErS�2��s��c�	T0 k� C�����(%2't ��1"t'!  ��*    ��� �2H&�E��*E�����!�,#W�Ec _Er[�2��c��c�T0 k� �����(%2't ��1"t'!  ��*    ��� �2H&�E��+E����!�,3[�Ec`Er_�2��c��c�T0 k� �����(%2't ��1"t'!  ��*    ��� �2H'�E��+E����!�,3[�EcbEbc�2��c��c�T0 k� �����(%2't ��1"t'!  ��*    ��� �"H(�E��,E����!�,3[�EcdEbg�"��c��c�T0 k� �����(%2't ��1"t'!  ��*    ��� �"D*�E��,E���'�!�,3[�EcgEbo�"��c��c�T0 k� �����(%2't ��1"t'!  ��*    ��� �"D+�E��-D�è�/�!�,3[�EciEbo�"��c��c�T0 k� �����(%2't ��1"t'!  ��*    ��� �"D,�E��-D�˪�7�|,3_�EckEbs�"��c��c� T0 k� �����(%2't ��1"t'!  ��*    ��� �"D-#�E��-D�ϫ�?�|,3c�ESmEbw�"��c��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �"D/'�E�-D�߭�O�|,3g�ESpEb{�"��c��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �"H0+�E�-D���W�|,3k�ESrEb| "��c��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �"H2�+�E�-D���_�|,3k�EStEb|"��S��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �"H3�/�E�-D���g�|,3o�ESuEb�"��S��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �"H4�3�E� -D����o�|,3s�ESwER�"��S��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �"L6�7�E�(.D����|,3w�ESzER�
"��S��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �"L8�;�E�,/D�����|,3{�ES|ER���S��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �"P9�;�E�0/D�����|,3{�ES}ER���S��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �"P:�?�E�40D�����|,3�ESER���S��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �"T<�?�E�80D�����|,3�ES�ER���S��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �X>�C�E�@1D�#����|,3��ES�C���c��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �X@�C�E�D2F +�0��|,3��EC C���c��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �\A�G�E�D2F /�0��|,3��EB�C���c��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �`B�G�E�H2F 7�0��|,3��EB�~C���c��c��T0 k� �����(%2't ��1"t'!  ��*    ��� �dD�G�E�L3F ;�0è|,3��EB�~C�|��c��c��T0 k� �{���(%2't ��1"t'!  ��*    ��� ��dE�K�E�L3F C�0˩|,3��EB�}C�|��c��c��T0 k� �s��w�(%2't ��1"t'!  ��*    ��� ��lG�K�E�P3F O�0׫|,3��EB�|C�x!�c��c��T0 k� �o��s�(%2't ��1"t'!  ��*    ��� ��pH�K�E�T3D�S�0߬|,3��EB�{C�t#��c��c��T0 k� �o��s�(%2't ��1"t'!  ��*    ��� ��tJ�K�E�T3D�W�0�|,3��EB�zC�p$��c��c��T0 k� �k��o�(%2't ��1"t'!  ��*    ��� ��xK�K�E�T3D�_�0�|,3��EB�yC�p&��	c��c��T0 k� �g��k�(%2't ��1"t'!  ��*    ��� ��|L�K�E�X3D�c� �|,3��C��yC�l'��
c��c��T0 k� �c��g�(%2't ��1"t'!  ��*    ��� ���M�K�ATX3D�k� ��|,3��C��xC�h)��s��c��T0 k� �c��g�(%2't ��1"t'!  ��*    ��� ���N cK�ATX3Epo� ��|,3��C��wC�d*��s��c��T0 k� �g��k�(%2't ��1"t'!  ��*    ��� ���P cK�ATX3Ep{�!�|,3��C��uC�\-��s��c��T0 k� �c��g�(%2't ��1"t'!  ��    ��� ���Q cK�ATX3Ep���|,3��E��tC�X/��s��c��T0 k� �_��c�(%2't ��1"t'!  ��    ��� ���R cK�ATX3Ep����|,3��E��sERT0��s��c��T0 k� �[��_�(%2't ��1"t'!  ��    ��� ���S �K�ATX3Ep����|,3��EҼrERP2��s��c��T0 k� �W��[�(%2't ��1"t'!  ��    ��� ���T �K�ATX3Ep����|,3��EҸqERL3r�s��c��T0 k� �S��W�(%2't ��1"t'!  ��    ��� ���U �K�ATX3Ep���#�|,3��EҰqERD4r�s��c��T0 k� �O��S�(%2't ��1"t'!  �    ��� ��W �K�AT3E��1/�|,3��EҤoER<7r�s��c��T0 k� �G��K�(%2't ��1"t'!  �    ��� ��XK�AP3E��13�|,3��AR�nER88r����c��T0 k� �;��?�(%2't ��1"t'!  ��    ��� ��YK�AP2E��1;�|,3��AR�mER4:�����c��T0 k� �3��7�(%2't ��1"t'!  ��    ��� ��ZK�AP2E��1?�|,3��AR�mER,;����c��T0 k� �/��3�(%2't ��1"t'!  ��    ��� ��[K�AL2E��1C�|,3��AR�lAR(<���w�c��T0 k� �'��+�(%2't ��1"t'!  ��    ��� ��\K�C�L1E��1K�|,3��AR�kAR$>���s�c��T0 k� �#��'�(%2't ��1"t'!  ��    ��� ��]�K�C�H1E��!O�|,3��AR�jAR ?���k�c��T0 k� ����(%2't ��1"t'!  ��    ��� ��^�K�C�D1E��!S�|,3��AR�jAR@��Sg�c��T0 k� ���#�(%2't ��1"t'!  ��    ��� ��_�K�C�D0E��!W�|,3��AR|iARA�  Sc�c��T0 k� �'��+�(%2't ��1"t'!  ��    ��� ��`�K�C�@0E���!_�|,3��ARxhARB�!S[�c��T0 k� �'��+�(%2't ��1"t'!  ��    ��� ���`�G�C�</F ��!c�|,3��ARpgARD�"SS�c��T0 k� �#��'�(%2't ��1"t'!  ��    ��� ��a�G�C�8.F ��!g�|,3��ARlgARE�"SO�c��T0 k� �#��'�(%2't ��1"t'!  ��    ��� ��c�C�C�4-F ��!s�|,3��ARdeARG�$SC�c��T0 k� ����(%2't ��1"t'!  ��    ��� ��c�C�C�0,F � !w�|,3��AR`eAR H�%S;�c��T0 k� ����(%2't ��1"t'!  ��    ��� ��$d�?�C�,,F �!�|,3��AR\dAQ�I�&S3�c��T0 k� ����(%2't ��1"t'!  ��    ��� ��,d�?�C�(+F �!��|,3��ARTcAQ�J�'S+�c��T0 k� ����(%2't ��1"t'!  ��    ��� ��4e�;�C�$*F ���|,3��ARPcAQ�K� 'S#�c��T0 k� �����(%2't ��1"t'!  ��    ��� ��<e7�C� )F ���|,3��ARLbAQ�L�$(C�c��T0 k� ������(%2't ��1"t'!  ��    ��� ��De7�C�(Lp�	��|,3��ARHbAQ�M�()C�c��T0 k� ������(%2't ��1"t'!  ��    ��� ��Lf3�C�'Lp���|,3��ARDaAQ�N�(*C�c��T0 k� ������(%2't ��1"t'!  ��    ��� �sTf/�C�'Lp���|,3��AR@`AQ�O�,*C�c��T0 k� ������(%2't ��1"t'!  ��    ��� �sXf/�C�&Lp���|,3��AR<`AQ�P�0+C�c��T0 k� ������(%2't ��1"t'!  ��    ��� �s`f+�C�%Lq ��|,3��AR8_AQ�Q�4,B��c��T0 k� ������(%2't ��1"t'!  ��    ��� �shf+�C�$Lq��|,3��AR4_AQ�R�8-B�c��T0 k� ������(%2't ��1"t'!  ��    ��� �spf'�C� "Lq��|,3��AR0^AQ�S�8-B�c��T0 k� ������(%2't ��1"t'!  ��    ��� �sxf#�C��!Lq��|,3��AR,]AQ�T�<.B�c��T0 k� �����(%2't ��1"t'! �    ��� �s�f�C��Lq��|,3��AR$\AQ�V�@/bۻc��T0 k� �����(%2't ��1"t'! ��    ��� �s�f�C��Lq���|,3��AR \AQ�W�D0bӻc��T0 k� �����(%2't ��1"t'! ��    ��� ���f�C��Lq���|,3��AR[AQ�X�H1bϺc��T0 k� �����(%2't ��1"t'! ��    ��� ���e�C��Lq���|,3��AR[AQ�Y�L1bǺc��T0 k� ҋ����(%2't ��1"t'!
 ��    ��� ���e#�L��Lq ���|,3��ARZAQ�Y�L2búc��T0 k� �����(%2't ��1"t'! ��    ��� ���e#�L��L�$ ���|,3��ARZAQ�Z�P3b��c��T0 k� �s��w�(%2't ��1"t'! ��    ��� ���d#�L��L�("q��|,3��ARYAQ�[�T3r��c��T0 k� �g��k�(%2't ��1"t'! ��    ��� ���d#�L��L�,#q��|,3��ARYAQ�\�T4r��c��T0 k� �_��c�(%2't ��1"t'! ��    ��� ���c#�L��L�0%q��|,3��ARXAQ�]�X4r��c��T0 k� �S��W�(%2't ��1"t'! ��   ��� ���b#�L��L�4&r�|,3��ARXAQ�]�X5r��c��T0 k� �G��K�(%2't ��1"t'! ��    ��� ���b#�L�L�4'r�|,3��ARWAQ�^�\6r��c��T0 k� �;��?�(%2't ��1"t'! ��    ��� ���a#�L�L�8)r�|,3��AR WAQ�_�`6���c��T0 k� �3��7�(%2't ��1"t'! ��    ��� ���`#�L�L�<*r�|,3��AQ�VAQ�`�`7���c��T0 k� �'��+�(%2't ��1"t'! ��    ��� ���_#�L�L�@+r�|,3��AQ�VAQ�`�d7���c��T0 k� ���(%2't ��1"t'! ��    ��� ���_#�M�L�D-r�|,3��AQ�VAQ�a�d8���c��T0 k� ���(%2't ��1"t'! ��    ��� ���^#�M�L�D.r#�|,3��AQ�UAQ�b�h8���c��T0 k� ���(%2't ��1"t'! ��    ��� ���]"��M�L�H/r+�|,3��AQ�UAQ�c�h9��c��T0 k� �����(%2't ��1"t'! ��    ��� ���\"��M�L�L1r/�|,3��AQ�TAQ�c�l9�{�c��T0 k� �����(%2't ��1"t'! ��    ��� ���["��M�L�P2r3�|,3��AQ�TAQ�d�p:�w�c��T0 k� �����(%2't ��1"t'! ��    ��� �s�Z"��M�
L�P3�7�|,3��AQ�TAQ�e�p:�s�c��T0 k� �����(%2't ��1"t'!  ��    ��� �t Y"��M�	L�T4�?�|,3��AQ�SAQ�e�t;�o�c��T0 k� �����(%2't ��1"t'!! ��    ��� �tW"��M�L�X5�C�|,3��AQ�SAQ�f�t;�k�c��T0 k� �����(%2't ��1"t'!" ��    ��� �tV"��M�L�X6�G�|,3��AQ�RAQ�g�x<�c�c��T0 k� �����(%2't ��1"t'!# ��    ��� �tU"��L�L�\8�K�|,3��AQ�RAQ�g�x<�_�c��T0 k� �����(%2't ��1"t'!$ ��    ��� �tT"��L�L�`9�S�|,3��AQ�RAQ�h�|=�[�c��T0 k� �����(%2't ��1"t'!% ��    ��� �tS"��L�|L�`:�W�|,3��AQ�QAQ�h�|=�W�c��T0 k� �����(%2't ��1"t'!& ��    ��� �tQ"��L�xL�d;�[�|,3��AQ�QAQ�i�>�S�c��T0 k� �����(%2't ��1"t'!' ��    ��� �t P"��L�tL�h<�\ |,3��AQ�QAQ�j�>�O�c��T0 k� �����(%2't ��1"t'!( ��    ��� �t$N"��L�pL�h=�`|,3��AQ�PAQ�j�?�K�c��T0 k� �w��{�(%2't ��1"t'!) ��    ��� �d(M"��L�lL�l>�d|,3��AQ�PAQ�k�?�G�c��T0 k� �k��o�(%2't ��1"t'!* ��    ��� �d,L"��L�h L�l?�h|,C��AQ�PAQ�k�@�C�c��T0 k� �_��c�(%2't ��1"t'!+ ��    ��� �d0J"��L�g�L�p@�l|,C��AQ�OAQ|l�@�?�c��T0 k� �W��[�(%2't ��1"t'!, ��    ��� �d4I"��C�c�L�tA�p|,C��AQ�OAQ|l�@;�c��T0 k� �K��O�(%2't ��1"t'!, ��    ��� �d8G"��C�_�L�tB�t|,C��AQ�OAQxm�A7�c��T0 k� �?��C�(%2't ��1"t'!- ��    ��� �d<F"��C�[�L�xC�x|,C��AQ�NAQxn�A3�c��T0 k� �3��7�(%2't ��1"t'!. ��    ��� �d@D"��C�W�L�xD�||,C��AQ�NAQxn�B/�c��T0 k� �+��/�(%2't ��1"t'!/ ��    ��� �d@B"��C�S�L�|E��|,C��AQ�NAQto�B+�c��T0 k� ���#�(%2't ��1"t'!0 ��    ��� �dDA"��ECO�L�|F��|,C��AQ�MAQto�B+�c��T0 k� � � (%2't ��1"t'!0 ��   ��� �dH?"��ECK�L��G��|,C��AQ�MAQpp�C'�c��T0 k� ��(%2't ��1"t'!1 ��    ��� �4H>"��ECG�L��G��|,S��AQ�MAQpp�C#�c��T0 k� ��� (%2't ��1"t'!2 ��    ��� �4L<"��ECC�L�|H��	|,S��AQ�MAQlq�C�c��T0 k� ����(%2't ��1"t'!2 ��    ��� �4L;"��EC?�L�|H��	|,S��AQ�MAQlq�D�c��T0 k� ����(%2't ��1"t'!3 ��    ��� �4P9"��EC7�L�|I��
|,S��AQ�MAQhq�D�c��T0 k� ����(%2't ��1"t'!3 ��    ��� �4P7"��EC3�L�|I��|,S��AQ�MAQhr�E�c��T0 k�  ���(%2't ��1"t'!4 ��    ��� �dP6"��E3/�L�|J��|,S��AQ�MAQhr�E�c��T0 k�  �	��	(%2't ��1"t'!4 ��    ��� �dT4��E3+�L�|J��|,S��AQ�MAQds�E�c��T0 k�  �
��
(%2't ��1"t'!5 ��    ��� �dT2��E3#�Lq|K��|,S��AQ�MAQds�F�c��T0 k�  ���(%2't ��1"t'!5 ��    ��� �dT0��E3�LqxK��|,S��AQ�MAQ`t�F�c��T0 k�  ���(%2't ��1"t'!6 ��    ��� �dT/��E3�LqxL��|,S��AQ�MAQ`t�F�c��T0 k� ����(%2't ��1"t'!6 ��    ��� �dT/��CC�LqxL��|,S��AQ�MAQ`u�G�c��T0 k� ����(%2't ��1"t'!6 ��   ��� �dT0��CC�LqxM��|,S��AQ�MAQ\u�G��c��T0 k� ����(%2't ��1"t'!7 ��    ��� �TT0R��CC�LqxM��|,S��AQ�MAQ\u�G��c��T0 k� �x�|(%2't ��1"t'!7 ��    ��� �TT0R��CC�FxN��|,S��AQ�MAQ\v�G��c��T0 k� �l�p(%2't ��1"t'!7 ��    ��� �TP1R��CC�FxN��|,S��AQ�MAQXv�H��c��T0 k� �`�d(%2't ��1"t'!8 ��    ��� �TP1R��CC�FxN��|,S��AQ�MAQXw�H��c��T0 k� �T�X(%2't ��1"t'!8 ��    ��� �TP1R��CC�FxO��|,S��AQ�MAQXw�H�c��T0 k� �L�P(%2't ��1"t'!8 ��    ��� ��L2R��CC�FxO��|,S��AQ�LAQTw�I�c��T0 k� �@�D(%2't ��1"t'!8 ��   ��� ��L2R��CR��E�xP��|,S��AQ�LAQTx�I�c��T0 k� �4�8(%2't ��1"t'!9 ��    ��� ��L2R��CR��E�|P��|,S��AQ�LAQTx�I�c��T0 k� �(�,(%2't ��1"t'!9 ��    ��� ��H2R��CR��E�|Q��|,S��AQ�LAQPx�I�c��T0 k� � �$(%2't ��1"t'!9 ��    ��� ��H3R��CR��E�|Qr�|,S��AQ�LAQPy�J�c��T0 k� ��(%2't ��1"t'!9 ��    ��� ��D3R��CR��E��Qr�|,S��AQ�LAQPy�J�c��T0 k� ��(%2't ��1"t'!9 ��    ��� ��D3R��CR��B�Qr�|,S��AQ�LAQLy�Jߪc��T0 k� �� �  (%2't ��1"t'!9 ��    ��� ��D3R��CR��B�Rr�|,S��AQ�LAQLz�Jߪc��T0 k� ��!��!(%2't ��1"t'!9 ��    ��� ��@4R��CR��B�Rr�|,S��AQ�LAQLz�K۪c��T0 k� ��#��#(%2't ��1"t'!9 ��    ��� �4@4R��CR��B�Rr�|,S��AQ�LAQL{�K۪c��T0 k� ��$��$(%2't ��1"t'!9 ��    ��� �4<4R��CR��B�R��|,S��AQ�LAQH{�Kתc��T0 k� ��%��%(%2't ��1"t'!9 ��    ��� �484R��CR��K��R��|,S�AQ�LAQH{�Kתc��T0 k� ��'��'(%2't ��1"t'!9 ��    ��� �484R��Cb��K��R��|,S�AQ�LAQH{�LӪc��T0 k� ��(��((%2't ��1"t'!9 ��    ��� �444R��Cb��K��R��|,S�AQ�LAQD|�Lөc��T0 k� ��)��)(%2't ��1"t'!8 ��    ��� �444R��Cb��K��R��|,S�AQ�LAQD|�Lϩc��T0 k� ��+��+(%2't ��1"t'!8 ��    ��� �404R��Cb��K��R��|,S�AQ�LAQD|�Lϩc��T0 k� ��,��,(%2't ��1"t'!8 ��    ��� �4,4R��Cb��K��S��|,S�AQ�LAQD}�M˩c��T0 k� ��-��-(%2't ��1"t'!8 ��    ��� �4(4R��IR��K��S��|,S�AQ�LAQ@}�M˩c��T0 k� �.��.(%2't ��1"t'!8 ��    ��� �4(4R��IRۿK��S��|,S�AQ�LAQ@}��Mǩc��T0 k� �x0�|0(%2't ��1"t'!7 ��    ��� �4$4R��IR۾K��S��|,S�AQ�LAQ@~��Mǩc��T0 k� �p1�t1(%2't ��1"t'!7 ��    ��� �4 4R��IRۼK��Sr�|,S�AQ�KAQ@~��Néc��T0 k� �d2�h2(%2't ��1"t'!7 ��    ��� �D4R��IR׺K��Ss |,S�AQ�KAQ<~��Nèc��T0 k� �X4�\4(%2't ��1"t'!6 ��    ��� �D3R��Ib׹K��Ss|,S�AQ�KAQ<~��N��c��T0 k� �L5�P5(%2't ��1"t'!6 ��    ��� �D3R��Ib׷K��Ss|,S�AQ�KAQ<��N��c��T0 k� �D6�H6(%2't ��1"t'!5 ��    ��� �D3R��Ib׶K��Ss|,S�AQ�KAQ<��N��c��T0 k� �87�<7(%2't ��1"t'!5 ��    ��� �D2R��Ib״K��S�|,S�AQ�KAQ<��O��c��T0 k� �,9�09(%2't ��1"t'!5 ��    ��� �42R��Ib׳K��S�|,S�AQ�KAQ8��O��c��T0 k� � :�$:(%2't ��1"t'!4 ��   ��� �42R��IRײK��T�|,S�AQ�KAQ8���O��c��T0 k� ;�;(%2't ��1"t'!4 ��    ��� �42R��IRױK��T�|,S�AQ�KAQ8��O��c��T0 k� =�=(%2't ��1"t'!3 ��    ��� �4 1R��IRׯK��T�|,S�AQ�KAQ8��O��c��T0 k�  >�>(%2't ��1"t'!2 ��    ��� �3�1R��IR׮K��T�|,S�AQ�KAQ4��O��c��T0 k� �?��?(%2't ��1"t'!2 ��    ��� �3�1R��IR׭K��T�|,S�AQ�KAQ4��P��c��T0 k� �A��A(%2't ��1"t'!1 ��    ��� �3�0R��Ib׬K��T� |,S�AQ�KAQ4~��P��c��T0 k� ��B��B(%2't ��1"t'!0 ��    ��� �3�0R��Ib׫K��T� |,S�AQ�KAQ4~��P��c��T0 k� ��C��C(%2't ��1"t'!0 ��    ��� �3�0R��IbתK��T�$|,S�AQ�KAQ4~��P��c��T0 k� ��D��D(%2't ��1"t'!/ ��    ��� �3�0R��IbתK��T�(|,S�AQ�JAQ0~��P��c��T0 k� ��F��F(%2't ��1"t'!. ��    ��� �3�/R��IbשK��T�(|,S�AQ�JAQ0}��P��c��T0 k� ޴G��G(%2't ��1"t'!. ��    ��� �3�/R��IRרK��T�,|,S�AQ�JAQ0}��Q��c��T0 k� ��H��H(%2't ��1"t'!- ��    ��� �C�/R��IRקK��T�,|,S�AQ�JAQ0}��Q��c��T0 k� ��J��J(%2't ��1"t'!, ��    ��� �C�/R��IRקK��T�0|,S�AQ�JAQ0}��Q��c��T0 k� ��K��K(%2't ��1"t'!+ ��    ��� �C�.R��IRצK��U�0|,S�AQ�JAQ0}��Q��c��T0 k� ��L��L(%2't ��1"t'!* ��   ��� �C�.R��IRצK��U�4|,S{�AQ�JAQ,|��Q��c��T0 k� �|N��N(%2't ��1"t'!) ��    ��� �C�.R��IbץK��U�8|,S{�AQ�JAQ,|��Q��"���T0 k� �pO�tO(%2't ��1"t'!( ��    ��� �C�.R��IbץK��U�8|,S{�AQ�JAQ,|��R��"���T0 k� �hP�lP(%2't ��1"t'!( ��    ��� �C�.R��IbפK��U�<
|,S{�AQ�JAQ,|��R��"���T0 k� �\Q�`Q(%2't ��1"t'!' ��    ��� �C�-R��IbפK��U�<	|,S{�AQ�JAQ,|��R��"���T0 k� �PS�TS(%2't ��1"t'!& ��    ��� �C�-R��IbפK��U�@|,S{�AQ�JAQ,{��R��"���T0 k� �DT�HT(%2't ��1"t'!% ��    ��� �C�-R��IRףK��U�@|,S{�AQ�JAQ({��R��"���T0 k� �<U�@U(%2't ��1"t'!# ��    ��� �C�-R��IRףK��U�D|,S{�AQ�JAQ({��R��"���T0 k� �0W�4W(%2't ��1"t'!" ��    ��� �C�-R��IRףK��U�D|,S{�AQ�JAQ({��R��"���T0 k� �$X�(X(%2't ��1"t'!! ��    ��� �C�,R��IRףK��U�H|,S{�AQ�JAQ({��S��"���T0 k� �Y�Y(%2't ��1"t'!  ��    ��� �C�,R��IRףK��U�H|,S{�AQ�JAQ({��S��"���T0 k� �Z�Z(%2't ��1"t'! ��    ��� �C�,R��IbףK��U�L|,S{�AQ�JAQ(z��S��"���T0 k� \�\(%2't ��1"t'! ��    ��� �C�,R��IbףK��U�L |,S{�AQ�JAQ(z��S��c��T0 k� �]��](%2't ��1"t'! ��    ��� �C�,R��IbףK��U�S�|,S{�AQ�IAQ$z��S��c��T0 k� �^��^(%2't ��1"t'! ��    ��� �C�+R��IbףK��U�S�|,S{�AQ�IAQ$z��S��c��T0 k� �`��`(%2't ��1"t'! ��    ��� �C�+R��IbףK��V�S�|,S{�AQ�IAQ$z��S��c��T0 k� �a��a(%2't ��1"t'! ��    ��� �C�+R��L�ףK��V�S�|,S�AQ�IAQ$z��S��c��T0 k� �b��b(%2't ��1"t'! ��    ��� �C�+R��L�ףK��V�S�|,S�AQ�IAQ$y��T��c��T0 k� �d��d(%2't ��1"t'! ��    ��� �C�+R��L�ףK��V�S�|,S�AQ�IAQ$y��T��c��T0 k� �e��e(%2't ��1"t'! ��    ��� �C�*R�L�ףK��V�S�!�,S��AQ�IAQ$y��T��c��T0 k� �g��g(%2't ��1"t'! ��    ��� �C�*R�L�ףK��V�S�!�,S��AQ�IAQ y��T��c��T0 k� ��i��i(%2't ��1"t'! ��    ��� �C�*R�L�ףK��V�S�!�,S��AQ�IAQ y��T��c��T0 k� ��j��j(%2't ��1"t'! ��    ��� �C�*R�L�ףK��V�S�!�,S��AQ�IAQ x��T��"���T0 k� ��k��k(%2't ��1"t'! ��    ��� �C�*R�L�ףK��V�S�!�,S��AQ�IAQ x��T��"���T0 k� �tm�xm(%2't ��1"t'! ��    ��� �C�*{�L�ףK��V�S�!�,S��AQ�IAQ x��T��"���T0 k� �hn�ln(%2't ��1"t'!
 ��    ��� �C�){�L�ףK��V�S�!�,S��AQ�IAQ x��U��"���T0 k� �`o�do(%2't ��1"t'!	 ��    ��� �C�){�L�ףK��V�S�!�,S��AQ�IAQ x��U��"���T0 k� �Tq�Xq(%2't ��1"t'! ��    ��� �C�){�L�ףK��V�S�!�,S��AQ�IAQ x��U��"���T0 k� �Hr�Lr(%2't ��1"t'! ��    ��� �C�){�L�ףK��V�W�!�,S��AQ�IAQ x��U��"���T0 k� �<s�@s(%2't ��1"t'! ��    ��� �C�){�L�ףK��V�W�|,S��AQ�IAQx��U��"���T0 k� �4t�8t(%2't ��1"t'! ��    ��� �C�)w�L�ףB�VsW�|,S��AQ�IAQw��U�"���T0 k� �(v�,v(%2't ��1"t'! ��    ��� �C�)w�L�ףB�VsW�|,S��AQ�IAQw��U�"���T0 k� �w� w(%2't ��1"t'!  ,�    ��� �C�(w�L�ףB�VsW�|,S��AQ�IAQw��U�"���T0 k� �x�x(%2't ��1"t'!  ��    ��� �C�(w�L�ףB�VsW�|,S��AQ�IAQw��U�c��T0 k� �z�z(%2't ��1"t'! ��   ��� �C�(w�L�ףB�VsW�|,S��AQ�IAQw��U�c��T0 k� ��{� {(%2't ��1"t'! ��    ��� �C�(w�L�ףE��VsW�|,S��AQ�IAQw��V{�c��T0 k� �|��|(%2't ��1"t'! ��    ��� �C�(w�L�ףE��UsW�|,S��AQ�IAQw��V{�c��T0 k� �}��}(%2't ��1"t'! ��    ��� �3�(s�L�ףE��UsW�|,S��AQ�IAQw��V{�c��T0 k� ���(%2't ��1"t'! ��    ��� �3�("s�L�ףE��UsW�|,S��AQ�IAQv��V{�c��T0 k� Ѐ�Ԁ(%2't ��1"t'! ��    ��� �3�("s�L�ףE��UcW�|,S��AQ�HAQv��V{�c��T0 k� ā�ȁ(%2't ��1"t'! ��    ��� �3�'"s�L�ףE��UcW�!�,S��AQ�HAQv��V{�c��T0 k� �����(%2't ��1"t'! *�    ��� �3�'"s�@�ףE��UcW�!�,S��AQ�HAQv��Vw�c��T0 k� �����(%2't ��1"t'! ��    ��� �3�'"s�@�ףE��TcW�!�,S��AQ�HAQv��Vw�c��T0 k� �����(%2't ��1"t'! ��    ��� �3�'"s�@�ףE��TcW�!�,S��AQ�HAQv��Vw�c��T0 k� �����(%2't ��1"t'! ��    ��� �3�'"s�@�ףE��T3W�!�,S��AQ�HAQv��Vw�c��T0 k� �����(%2't ��1"t'! ��    ��� �3�'"s�@�ףCA�S3W�!�,S��AQ�GAQv��Vw�c��T0 k� L�����(%2't ��1"t'! ��    ��� �3�&"o�@�ףCA�R3W�!�,S��AQ�GAQv��Ww�c��T0 k� Lx��|�(%2't ��1"t'! ��    ��� �3�&"o�@�ףCA�R3S�!�,S��AQ�GAQv��Ws�c��T0 k� Lp��t�(%2't ��1"t'! ��    ��� �3|&"o�@�ףCA�R3S�!�,S��AQ�GAQu��Ws�c��T0 k� Ld��h�(%2't ��1"t'! ��    ��� �3|%"o�AףCA�R3S�!�,S��AQ�GAQu��Ws�c��T0 k� LX��\�(%2't ��1"t'! ��    ��� �3x%"o�AףCA�Q3S�!�,S��AQ�FAQu��Ws�c��T0 k� �P�T(%2't ��1"t'! ��    ��� �3x$"o�AףCA�P3S�|,S��AQ�FAQu��Ws�c��T0 k� �D�H(%2't ��1"t'! ��    ��� �3t$"o�AףCA�O3S�|,S��AQ�FAQu��Ws�c��T0 k� �8�<(%2't ��1"t'! ��    ��� �3p$"o�AףCA�O3S�|,S��AQ�FAQu��Wo�c��T0 k� �0~�4~(%2't ��1"t'! ��    ��� ��l#"o�AףCA�N3S�|,S��AQ�EAQu��Wo�c��T0 k� �$~�(~(%2't ��1"t'!  ��    ��� ��l""k�AףCA�M3S�|,S��AQ�EAQu��Wo�c��T0 k� ,~�~(%2't ��1"t'!  ��    ��� ��h""k�AףCA�L3S�|,S��AQ�EAQu��Wo�c��T0 k� ,}�}(%2't ��1"t'!  -�    ��� ��d!"k�AףCQ�KCS�|,S��AQ�EAQu��Wo�c��T0 k� ,}�}(%2't ��1"t'!  ��    ��� ��` "k�AףCQ�KCS�|,S��AQ�EAQu��Wo�c��T0 k� +�}��}(%2't ��1"t'!  ��    ��� ��\ "k�AףCQ�KCS�|,S��AR DAQu��Wo�c��T0 k� +�{��{(%2't ��1"t'!  ��    ��� ��e?�C`�-D��$}�"|/���E��]AP�'	p�A�`>3�T0 k� ��S��S(%2't ��1"t'!  ��     � < � d3�C`�,D��%}�!|/���E`�]AP�'	p�A�\>3�
T0 k� ��R��R(%2't ��1"t'!  ��     � < ��c+�C`�+D��&��!|/���E`�^AP�'	��A�X>3�
T0 k� ��Q��Q(%2't ��1"t'!  ��     � < ��b�C`�(D��)�� |, ���E`�_AP�'	��A�T>3�	T0 k� ��O��O(%2't ��1"t'!  ��     � < ��a��C`�'D��*�� |,���E`�`AP�'	��A�P>3�	T0 k� ��M��M(%2't ��1"t'!  ��     � < ��`��C`�&D��+�� |,��E`�`AP�'	��A�L>3�T0 k� ��K��K(%2't ��1"t'!  ��     � < ��_���Cp�$D��-�� |,��P�|aAP�'	p�A�H>3�T0 k� ��I��I(%2't ��1"t'!  ��     � <  ��_���Cp�#D��.�| |,��P�xaAP�'	p�A�D>3�T0 k� ��H��H(%2't ��1"t'!  ��     � <����^��Cp�!D��0�| |,��P�xbAP�'	p�A�@>3�T0 k� ��H��H(%2't ��1"t'!  ��     � <����]��Cp� F�1�x|,��P�tcAP�'	p�A�<>3�T0 k� ��G��G(%2't ��1"t'!  ��     � <����\�ߎCp�F�3�t|,���P�tcJ��'	p�A�8>3�T0 k� ��F��F(%2't ��1"t'!  ��     � <����[�ӎE �F�4�t|,���P�pdJ��'P�A0>3�T0 k� ��E��E(%2't ��1"t'!  ��     � <����Z�ˎE �F�6�p|,���P�leJ��'P�A,>3�T0 k� ��D��D(%2't ��1"t'!  ��     � <����Y�ÏE �F�7�p|,���P�leJ��'P�A(>3�T0 k� ��C��C(%2't ��1"t'!  ��     � <����X໏E �F�9�p|,���P�hfJ��'P�A$>3�T0 k� ��B��B(%2't ��1"t'!  ��     � <����W೏E �F�;�l|,���P�hfJ��'P�A>3�T0 k� ��@��@(%2't ��1"t'!  ��     � <����U�E �F�<�l|,���P�dgJ��'��A>3�T0 k� ��?��?(%2't ��1"t'!  ��     � <����T�B�F�>�h|,���P�dgJ��'��A>3�T0 k� ��>��>(%2't ��1"t'!  ��     � <���xS�B�E��?�h|,���P�`hJ��'��A>3�T0 k� ��=��=(%2't ��1"t'!  ��     � <���pR���B�E��A�h|,���P�\hJ��'��A>3�T0 k� ��;��;(%2't ��1"t'!  ��     � <��lP���B�E��C�d|,���P�\iJ��'��A >3�T0 k� ��<��<(%2't ��1"t'!  ��     � <��dO��B�E��D�d|,���P�XjJ��'��A�>3�T0 k� ��<��<(%2't ��1"t'!  ��     � <��`N�s�B�
E��F�`|,���P�XjJ��'��A�>3�T0 k� ��;��;(%2't ��1"t'!  ��     � <��XL�k�B�E��G�`|,���P�TkJ��'��A�>3�T0 k� ��;��;(%2't ��1"t'!  ��     � <��TK�c�B�E��I\|,���P�TkJ��'��A�>3�T0 k� �|:��:(%2't ��1"t'!  ��     � <��PJ�[�B�E��J\|,��P�TlJ� '��A�>3�T0 k� �|9��9(%2't ��1"t'!  ��     � <��HH�S�B�E��KX|,��E`PlJ� '��A�>3�T0 k� �x8�|8(%2't ��1"t'!  ��     � <��DG K�B�E��MT|,��E`LmJ�'��A�>3�T0 k� �t6�x6(%2't ��1"t'!  ��     � <��@E ?�B��E��NT|,��E`LmJ�'��A�>3�T0 k� �l5�p5(%2't ��1"t'!  ��     � <��<D 7�C ��E��P
P|,��E`HnJ�'��A�>3�T0 k� �h3�l3(%2't ��1"t'!  ��     � <��8B /�C ��E��Q
L|,��E`HnJ�'��A	��>3�T0 k� �d2�h2(%2't ��1"t'!  ��     � <��4A '�C ��E��R
H|,��EPDoJ�'��@	��>3�T0 k� �`0�d0(%2't ��1"t'!  ��     � <��0?@�C ��E��S
D|,�ߪEP@pJ�'��@	��>3�T0 k� �\/�`/(%2't ��1"t'!  ��     � <��,>@�C ��E��T
D|,�۪EP<pJ�'��@	��>3�T0 k� �\-�`-(%2't ��1"t'!  ��     � <��,<@�C ��E��U@|,�۫EP8qJ�'��@	��>3�T0 k� �X,�\,(%2't ��1"t'!  ��     � <��(;@�C ��E��V<|,�׫EP4qJ�'��@	��>3�T0 k� �T*�X*(%2't ��1"t'!  ��     � <���$9O��C ��E��W8|,�ӫE@0rJ�'��@	��>3�T0 k� �L,�P,(%2't ��1"t'!  ��     � <���$7O�C ��E��X4|,�ϬE@,rJ�'��@	��>3�T0 k� �H.�L.(%2't ��1"t'!  ��     � <��� 6��C ��E��Y0|,�ˬE@(rEa'0�@	��>3�T0 k� �@.�D.(%2't ��1"t'!  ��     � <��� 4��C ��E��Z-,|,?ǬE@$sEa'0�@	��>3�T0 k� �</�@/(%2't ��1"t'!  ��     � <���3�הC��E��[-(|,?ìE@ sEa&0�@	��>3�T0 k� �8.�<.(%2't ��1"t'!  ��     � <�� /2�ϔC��E��[- |,?��PpsEa&0�@	�|>3�T0 k� �H.�L.(%2't ��1"t'!  ��     � <�� /0�ǕC��E��\-|,?��PptEa&0�A	�x>3�T0 k� �T,�X,(%2't ��1"t'!  ��     � <�� //O��C��E��\-|,?��PptEa&��A	�t>3�T0 k� �\+�`+(%2't ��1"t'!  ��     � <�� /-O��C��E��]
M|,?��PptEa%��A	�p>3�T0 k� �`*�d*(%2't ��1"t'!  ��     � <�� /,O��I0��E��]
M|,﫭PpuEa %��A	�l>3�T0 k� �d(�h((%2't ��1"t'!  ��     � <�� /+O��I0��E��]
M|,吝P�uEa$%��B	�l>3�T0 k� �h'�l'(%2't ��1"t'!  ��     � <�� /)O��I0��E��^
M|,P�uEa$%��B	�h>3�T0 k� �l&�p&(%2't ��1"t'!  ��     � <�� /(O��I0��E��^
M |,P� vEa($��B	�d>3�T0 k� �p$�t$(%2't ��1"t'!  ��     � <�� /'?��I0��E��^
L�|,P��vEa($��C	�`>3�T0 k� �p#�t#(%2't ��1"t'!  ��     � <�� ?&?��I@��E��^
L�|,P��vEa,$��C	�`>3�T0 k� �t"�x"(%2't ��1"t'!  ��     � <�� ?$?{�I@��E��^
L�|,P��vEa,$��C	�\>3�T0 k� �x �| (%2't ��1"t'!  ��     � <�� ? "?k�I@��E��^
\�|,P��wEa0$
� D	�X>3�T0 k� ����(%2't ��1"t'!  ��     � <�� ? !?c�I@��E��^
\�|,P��wEa0$
�D	�X>3�T0 k� ����(%2't ��1"t'!  ��     � <�� ?$ ?[�E ��E��^
\�
|,��P�wEa0$
�D	�T>3�T0 k� ����(%2't ��1"t'!  ��     � <�� ?$?S�E ��E��^
\�
|,�{�P�xEa4$
�D	�T>3�T0 k� ����(%2't ��1"t'!  ��     � <�� ?(?K�E ��E��^
\�	|,�w�P�xEa4$
�E	�P>3�T0 k� ����(%2't ��1"t'!  ��     � <�� ?(?C�E ��C��] l�	|,�s�P�xJ�4$�E	�P>3�T0 k� ����(%2't ��1"t'!  ��     � <�� ?,?;�E ��C��] l�|,�k�P�xJ�4$�E	�P>3�T0 k� ����(%2't ��1"t'!  ��     � <�� ?0?3�E ��C��] l�|,�g�C��yJ�4$� E	�P>3�T0 k� ����(%2't ��1"t'!  �     � <��O0/+�E ��C��\ l�|,�c�C��yJ�4$�$E	�L>3�T0 k� ����(%2't ��1"t'! ��    � ; O4/#�E!�C��\ l�|,�_�C��yJ�4$�,F	�L>3�T0 k� ����(%2't ��1"t'! ��    � : O4/�E!�C��\ l�|,�[�C��yA4$�0F	�L>3�T0 k� ����(%2't ��1"t'! ��    � 9 O8/�E!�C��[ l�|,�W�C��yA4$�8F	�L>3�T0 k� ����(%2't ��1"t'! ��    � 8 O</�E!�C��[ l�|,S�C��yA4$�<F	�L>3�T0 k� ����(%2't ��1"t'! ��    � 7 O</�E!�C��Z l�|,O�C��yA8$�DG	�L>3�T0 k� ����(%2't ��1"t'! ��    � 6 ?@/�E!�C��Z l�|,K�C��yA8$�HG	�L>3�T0 k� ������(%2't ��1"t'! ��    � 5 ?@.��E!�C��Y l�|,G�C��xA8$�PG	�L>3�T0 k� ������(%2't ��1"t'! ��    � 3 ?D.��E!�C��Y l�|,C�C��x@�8$�TG	�P>3�T0 k� ������(%2't ��1"t'! ��    � 1 #?H��E!�C��X l�|,C�C��x@�8$�\G	�P>3�T0 k� ������(%2't ��1"t'! ��    � / &?H��E!�C��W l�|,?�C��x@�8$
�dG
�P>3�T0 k� ������(%2't ��1"t'! ��    � - )/L��E!�C��W l�|,;�C��w@�8#
�hG
�P>3�T0 k� �����(%2't ��1"t'! ��    � + ,/L��E!�C��V l�|,;�C��w@�8#
�pF
�T>3�T0 k� ����(%2't ��1"t'! ��    � ) //P��E!#�C��U l�|,7�C��vCA8#
�xF
�T>3�T0 k� ����(%2't ��1"t'! ��    � ' 2/P.ۯE!#�C��T l�|,�7�C��vCA8#
�|F
�X>3�T0 k� ����(%2't ��1"t'! ��    � % 5/T.۰E!'�C��S l�|,�3�C��uCA8"
��F
�X>3�T0 k� �#��'�(%2't ��1"t'! ��    � # 8/T
.ױE!+�C��S l�|,�3�EO�uCA8"
��E
�\>3�T0 k� �+��/�(%2't ��1"t'! ��    � ! ;/X	.ӲE!+�C��R
�|,�3�EO�tCA8!
��E�`>3�T0 k� �3��7�(%2't ��1"t'! ��    �  >/X.ϳE!/�C��Q
�|,�3�EO|sCA8!
��E�`=3�T0 k� �;��?�(%2't ��1"t'! ��    �  A/\.˴E!3�EL�P
�|,�3�EOxsCA8 
��D�d=3�T0 k� �C��G�(%2't ��1"t'! ��    �  D/\˶E!3�EL�O
�|,�/�EOprCA8
��D�h=3�T0 k� �K��O�(%2't ��1"t'! ��    �  G/`ǷE!7�EL�N
�|,/�E?lqE�8
��C�h=3�T0 k� �S��W�(%2't ��1"t'! ��    �  J/`øE!;�EL�ML�|,3�E?dpE�8
��C�l=3�T0 k� �_��c�(%2't ��1"t'! ��    �  M/dùE!;�EL�LL�|,3�E?`pE�8
��B�p<3�T0 k� �g��k�(%2't ��1"t'! ��    �  P/d��E!?�E<�KL�|,3�E?\oE�8
��B�t<3�T0 k� �o��s�(%2't ��1"t'! ��    �  S/h��E!C�E<�IL�|,3�E?TnE�8
��A�x<3� T0 k� �w��{�(%2't ��1"t'! ��    �  V/h��E!C�E<�HL�|,�3�E?PmE�8
��@�|;3� T0 k� �����(%2't ��1"t'! ��    � 	 Y/h��E!G�E<�G��|,�7�E?LkE�8
��@
��;3� T0 k� ������(%2't ��1"t'! ��    �  [/l��E!K�E<�F��|,�7�E?HjE�4
��?
��;3��T0 k� ������(%2't ��1"t'! ��    �  ]/l ��E!K�CL�D��|,�;�E?@iE�4
��>
��:3��T0 k� ����(%2't ��1"t'! ��    �   _/p ���E!O�CL�C��|,�;�E?<hE�4
��=
��:3��T0 k� ����(%2't ��1"t'! ��    ��� a/s����E!O�CL�B��|,�?�E/8gC�0
��=
��93��T0 k� ����(%2't ��1"t'! ��    ��� c�s����E!S�CL�@��|,�?�E/4eC�0
� <
��83��T0 k� ����(%2't ��1"t'! ��    ��� f�w����E!W�CL�?��|,�C�E/0dC�0
�;
��83��T0 k� ����(%2't ��1"t'! ��    ��� h�{����E!W�CL�=��|,�C�E/,bC�,
�:
��73��T0 k� �ë�ǫ(%2't ��1"t'! ��    ��� j�{����E![�CL�<��|,�G�E/(aC�,
�9
��63��T0 k� �˨�Ϩ(%2't ��1"t'! ��    ��� l�����E!_�CL�:��|,�K�E/$`C�(
� 8
��63��T0 k� �ӥ�ץ(%2't ��1"t'! ��    ��� n�����E!_�CL�9��|,�K�E/$^C�$
�(7
��53��T0 k� �ۢ�ߢ(%2't ��1"t'! ��    ��� p������E!c�CL�7��|,�O�E/ ]C�$
�06
��43��T0 k� ����(%2't ��1"t'! ��    ��� r������E!g�CL�5��|,�S�E/[C� 
�<5
��33��T0 k� ����(%2't ��1"t'! ��    ��� t�����E!g�CL�4��|,�S�E/ZC�

�D4
��23��T0 k� �����(%2't ��1"t'! ��    ��� v�����E!k�C\�2��|,�W�E/XC�	
�L3
��23��T0 k� ������(%2't ��1"t'! ��    ��� x�����E!o�C\�0��|,�[�EWC�
�T2
��13��T0 k� ����(%2't ��1"t'!  ��    ��� {�����E!o�C\�.�� |,�_�EUC�
�\0
��03��T0 k� ����(%2't ��1"t'!  -�    ��� }�����E!s�C\�-���|,�c�ETC�
�d/
��/c��T0 k� ����(%2't ��1"t'!  ��    ��� �����E!s�C\�+���|,�g�ERC��l.
��.c��T0 k� ���#�(%2't ��1"t'!  ��    ��� ������E!w�C\�)���|,�k�EQC��p-
��-c��T0 k� �'��+�(%2't ��1"t'!  ��    ��� �������E!{�C\�'���|,�o�B�PC� �x,
��,c��T0 k� �/��3�(%2't ��1"t'!  ��    ��� �������E!{�C\�%���|,�s�B�NC��Ҁ+
��+c��T0 k� �7��;�(%2't ��1"t'! ��    ��� �������E!�C\�#���|,�w�B�MC���҄*
��*c��T0 k� �?~�C~(%2't ��1"t'! ��    ��� �������E!��C\�!���|,�{�B�KC���Ҍ)
��)c��T0 k� �G|�K|(%2't ��1"t'! )�    ��� �������E!��C\����|,��B�JC���Ґ(
��'c��T0 k� �O|�S|(%2't ��1"t'! ��    ��� �������E!��Cl����|,߃�B�IC���Ҕ'
��&c��T0 k� �W}�[}(%2't ��1"t'! ��    ��� �������E!��Cl����|,B�HC���Ҙ&
� %c��T0 k� �_~�c~(%2't ��1"t'! ��    ��� �������E!��Cl����|,B�FC����%
�$c��T0 k� �g~�k~(%2't ��1"t'!  ��    ��� �������E!��Cl����|,B�EC����$�#c��T0 k� �o�s(%2't ��1"t'!  ��    ��� �������E!��Cl����|,B�DC����#�"c��T0 k� ���(%2't ��1"t'!  ��"    ��� �������E!��I\����|,B�CC����"�!c��T0 k� ы~��~(%2't ��1"t'!  ��"    ��� ������E!��I\���|,留B� @E0��� �c��T0 k� ѓ~��~(%2't ��1"t'!  ��"    ��� ������E��I\���|,頻B�$?E0���� c��T0 k� ћ����(%2't ��1"t'!  ��"    ��� ������E��I\���|,ﳋB�(>E0����$c��T0 k� ������(%2't ��1"t'!  ��"    ��� ������E��E<�	��|,��B�,=E0����$c��T0 k� ������(%2't ��1"t'!  ��"    ��� �����E��E<���|,��B�,<E0����(c��T0 k� ������(%2't ��1"t'!  ��"    ��� �����E��E<���|,ÉB�0;E0�����,c��T0 k� ������(%2't ��1"t'!  ��"    ��� �����E��E<���|,ǉB�4:E0�����,c��T0 k� ������(%2't ��1"t'!  ��"    ��� ����'�E��E<� ��|,ψB�89E0�����0c��T0 k� ������(%2't ��1"t'!  ��"    ��� ����+�E��E<����|,ӇB�@8E0�����0c��T0 k� ����Ð(%2't ��1"t'!  ��"    ��� ��'��/�E��E,�����|,ۇB�D7E0�����4c��T0 k� �Ǒ�ˑ(%2't ��1"t'!  ��"    ��� ��+��7�E�ÎE,�����|,�B�H6E0�����4c��T0 k� �ϕ�ӕ(%2't ��1"t'!  ��"    ��� ��3��;�E�ǎE,�����|,��B�L5E �����4c��T0 k� �ט�ۘ(%2't ��1"t'!  ��"    ��� ��C��G�E�ӏE,�����|,��B�X3E �����8c��T0 k� ����(%2't ��1"t'!  ��"    ��� ��K��K�E�׏E,�����|,���B�\2E �����8c��T0 k� ����(%2't ��1"t'!  ��"    ��� ��S��S�E�ېE,�����|,��B�d1E �����8c��T0 k� ����(%2't ��1"t'!  ��"    ��� ��[��[�E��E,�����|,��B�h0E ����	�8c��T0 k� �����(%2't ��1"t'!  ��"    ��� ��c��_�E��E,�����|,��B�p/E �����<c��T0 k� ������(%2't ��1"t'!  ��"    ��� ��k��g�E��E,�����|,��B�t.E �����<c��T0 k� �����(%2't ��1"t'!  ��"    ��� ��s��o�E��E,�����|,��B�|-E �����<c��T0 k� ����(%2't ��1"t'!  ��"    ��� ����s�E���E,�����|,�'�B߀,E ����<c��T0 k� ����(%2't ��1"t'!  ��"    ��� �����{�Eq��E�����|,�/�B߈+E ��� �<c��T0 k� ����(%2't ��1"t'!  ��"    ��� �������Er�E�����|,�7�Bߐ+E�����<c��T0 k� ����(%2't ��1"t'!  ��"    ��� �������Er�E�����|,�?�Bߘ*E�����<c��T0 k� ����(%2't ��1"t'!  ��"    ��� �������Er�E�����|,�G�Bߜ)E�����<c��T0 k� ���#�(%2't ��1"t'!  ��"    ��� �������Er�E�����|,�O�Bߤ(E������<c��T0 k� �#��'�(%2't ��1"t'!  ��"    ��� �������Er�E�����|,�W�B߬'E������<c��T0 k� �+��/�(%2't ��1"t'!  ��"    ��� �������Er�E�����|,�c�Bߴ'E������<c��T0 k� �/��3�(%2't ��1"t'!  ��"    ��� �������Er'�E�����|,�k�B߼&E������<c��T0 k� �3��7�(%2't ��1"t'!  ��"    ��� �������Er+�E�����|,�s�B��%E�����S<c��T0 k� �;��?�(%2't ��1"t'!  ��"    ��� �������Er/�B������|,�{�B��$I�����S<c��T0 k� �?��C�(%2't ��1"t'!  ��"    ��� �������Er7�B������|,���B��$I�����S<c��T0 k� �C��G�(%2't ��1"t'!  ��"    ��� �������Eb;�B������|,���B��#I�����S<c��T0 k� �7��;�(%2't ��1"t'!  ��"    ��� �������Eb?�B������|,���B��"I����S<c��T0 k� �3��7�(%2't ��1"t'!  ��"    ��� �������EbC�B�����|,���B��"I�����<c��T0 k� �/��3�(%2't ��1"t'!  ��"    ��� �������EbG�B�����|,���E�!I�����<c��T0 k� �+��/�(%2't ��1"t'!  ��"    ��� ������EbK�B�����|,���E  I �����<c��T0 k� �+��/�(%2't ��1"t'!  ��"    ��� ������EbO�B�����|,���EI �����<c��T0 k� �+��/�(%2't ��1"t'!  ��"    ��� �����EbS�B�����|,�ÍEI �����<c��T0 k� �'��+�(%2't ��1"t'!  ��" 
   ��� �����EbS�B�����|,�ˎEI �����<c��T0 k� �'��+�(%2't ��1"t'!  ��" 
   ��� ��'���EbW�B�ǿ�#�|,�ӎE$I �����<c��T0 k� �+��/�(%2't ��1"t'!  ��" 
   ��� ��/���Eb[�B�˽�'�|,�ێE0E�����<c��T0 k� �/��3�(%2't ��1"t'!  ��" 
   ��� ��;��#�ER[�B�Ӽ�+�|,��E�8E��s#��<c��T0 k� �3��7�(%2't ��1"t'!  ��" 
   ��� ��C��/�ER_�B�׺�3�|,��E�@E��s'��<c��T0 k� �;��?�(%2't ��1"t'!  ��" 
   ��� ��K��7�ER_�B�۹�7�|,���E�HE��s+��<c��T0 k� �;��?�(%2't ��1"t'!  ��" 
   ��� ��S��?�ERc�B�߷�?�|,���E�TE��s/��<c��T0 k� �?��C�(%2't ��1"t'!  ��" 
   ��� ��[��G�ERc�B���C�|,��E�\E���s3��@c��T0 k� �C��G�(%2't ��1"t'!  ��" 
   ��� ��k��[�E�c�B���S�|,��D�pE���s;��@c��T0 k� �C��G�(%2't ��1"t'!  ��" 
   ��� ��w��c�E�g�B����W�|,�#�D�xE���s?��@c��T0 k� �C��G�(%2't ��1"t'!  ��" 
   ��� ����k�E�g�B����_�|,�+�DЀE���sC��Dc��T0 k� �G��K�(%2't ��1"t'!  ��" 
   ��� �����s�E�g�B���g�|,�3�DЌDЗ�cG��Dc��T0 k� �G��K�(%2't ��1"t'!  ��" 
   ��� �����{�E�g�B���k�|,�?�DДDЛ�cG��Hc��T0 k� �G��K�(%2't ��1"t'!  ��" 
   ��� ����Ѓ�E�g�B���s�|,�G�DМDЛ�cK��Hc��T0 k� �G��K�(%2't ��1"t'!  ��" 
   ��� ����Џ�E�g�B���{�|,�O�DШDП�cO��Lc��T0 k� �C��G�(%2't ��1"t'!  ��" 
   ��� ����З�E�g�B�����|,�W�D�DУ�cO��Lc��T0 k� �C��G�(%2't ��1"t'!  ��" 
   ��� �                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \��m ]�!�!� � 
��  L   ^ ^	     � ��      �0 س�    ����   	             $�� �          �     ���  8	(
         ��q   � �
	   � ���    ��� ��     ��               J �� �         ��    ���   @
	"          ��F:    
	    �r;    ��F: �r;                      ( 	�� ��        �      ���    		'

           K��  5 5	     pX     K�� pX    ���              �� �          ���    ���  8	
          ��F   � �	    . �	-    ��u �O    �,��               a�� �          ��  %  ���  X
          	`  ��	      B�F�     	`�F�                             ���p              �  ���    0 0            �٢]          V ���    ��� ��    �^              	 C��          H0  �  ��@   8		�          D�)         j �9�     E{ �l    ��"             <��          �     ��@   0
            u�         ~ Ev_     u'h E�`    ���              ��          y�     ��@   (
"
           W�         � ���     W�I ��Y     �              	�� �         	 �P     ��@   H
w          ���        � [,h    ���� [Mi    ���               
 A �         
 �`     ��H   (
         ���k ��
	      � �4�    ���k �4�                              ����             �  ��@    0

 2              I   ��      ���      I ��                                                               �                               ��        ���          ��                                                                 �                          {�]  ��        �����  �� }T����@  ����ߡ                   x        ���     j  �  �
   �                          {    ��        ���       }  ��           "                                                �                          � � � p �� � � E � [ �������   	  
            
  8   y �� $��F       $ �c@ $ d@ D  d` �D �e� �D f� �d  f� ɤ  g  �� g` �D 0x  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ �� 0�  �� 0ʀ �( 0�  �� 0ɀ �h 0�  � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À���� � � }`���� � 
�\ V  
�| V ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���� � �����F  ������  
�fD
��L���"����D" � j  "  B   J jF�"     "�j  " ��
��
��"     
�j
�� 
  
 �
� �  �  
� ����  ��     � �  �   ��    ��     � �      ����  ��     � [          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �"      ��(T ���        � �T ���        �        ��        �        ��        �  
  ��    �
�� |         ��                         T�) , �� ��                                     �                ����            
�� �
���%��  �� ���               22 Christan Ruuttu     4:53                                                                        2  2     �7c� �Oc� �%Kb K"_%K#Zkj^5 kr^ �B� � 	B� � 
B� � � B� � � B� � B� �K � �K � �C. � � C6 � �C7 � �C9 � � C; � �
B�1 �B�0 � B�I � B�) �cV � � c^ � �
c� � � c� � c� �c�p � c�h �	 �
 �	!�! �"� �#�3$"� %"�&"� �'*�Z("� �Z )"� �J*� �J+
� � � ,"O z  "& r  "& r �/": r � 0"A z � 1"P z �  " r � 3"O z � 4"K z � !� r � !� r z7"  r � 8"O z � 9"K z � !� r  "& r � <"O z  "& r �>!� r � "< r                                                                                                                                                                                                                         �� R              @ 
      $ �     W P E [  ��        
            �������������������������������������� ���������	�
��������                                                                                          ��    �v�   ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E   �4, :� �@P���@���@�����                                                                                                                                                                                                                                                                                                                                           @U�                                                                                                                                                                                                                                             
      I    3    ��  4�J      '  	                           ������������������������������������������������������                                                                                                                                          �  ��             �          ��               	 
     ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� �������            5                    %    &      �   .�J      -                              ������������������������������������������������������                                                                        
                                                                     �  ��                P        �    �            	     ��  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���                                                                                                                                                                                                                                                       	                                                              
        �             


           �   }�                                              +                                          ��������    ������������������������������������  +�����������������������������������������������������ww�ww333wwwwwwww�ww�ww�ww�ww333wwww R > / 	                                � ��z" �\                                                                                                                                                                                                                                                                                    	�)n1n  )F)�        m      b      a            l      l            m                                                                                                                                                                                                                                                                                                                                                                                                          0   � ��  � ��  � #��  � #��  EZm*  �N ���(�������������i�����^�����&������������                 x�E : � {          �   & AG� �   �   
              �                                                                                                                                                                                                                                                                                                                                      p N K   �      ��               !��                                                                                                                                                                                                                            Y   �� �� Ѱ��      �� 9      ����������������������������������������� ��� ����� ����������� � �������� �������� ���� ������� �� ������������������� ���������� �������� �� ����� ����������������� ����������������� ��������� ����������������������� ���������  �� ��������� ��  ������������� ���������������  ���� ����� ������ ��� �������� �� �������� ������������������������� ��������������� ����������������������������� ����������� ����������������������������� ���� � ���             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    C      4      }                       8     �   �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �f ��     �f �$ ^$ �@       �       �     �   n 
� �     �f ��        p���� ��   p����      �       �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h  8���( ��  8���( �$ ^$   �  8                  $   ���(�� � ��� �� � ��� �$  � �  �� �  �      �      �����������J   g���        f ^�         ��	��            ��m|�������J���J�������      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                          �      �  a r!   f�"""""*��**"*�"�""�""v""*f   "  ""- ��"�"*"-""z"""""����            n   �  "  q  ��                          �  �                                 � gv"!g�vg�vggfvv|�b��r""gb"�vr�rgb��v���g���v���***�*q!q�"!a�!vwfqqr~� qw��q�~~q�����~~~�w~~w�w            �   ~   ��  ~~  �w      v    �                ggj�vvggvvgg!vg�g֪vvg�r�r��⢪rq**gjb�v�q*gjj*vv��gg�z�/�"!�"�*�""*z����qw�~q~ww��q~qwvq�w�`� ��� �w �~p w�p  ��                    �                        lggz�v��g        �       ggbvvrgggavvvqggav� �      ���w!z�w"""�!""*�"! ��        q� q�        `               �        �                      wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                           �  ��  �� �� ��� ��� +� )� ��  ��  ��  Lɢ Ě� �I�� ��                           "   "    
�� ��� ̼� �����̺�ۻ }�  wg            �   �   �   �   �   ��̷��� ˈ� ��� ��Ȩ�ۊ�����˻� |             ��" ��" ��"       �� �� �� �� ʪ}���w����˚����  ̽  ��  �w  ��  vv  ���"w��"   �  �  �  �  �� 
�w��~˚���   ��  ��  �p  }`  g`  m   }     �  ��  ��  ۽ 
}� 
wv	���ɪ���   �   �   w   �   v   p         �  �� �� ۽ }� �wv
��暪���   �   �   w   �   v   �   �     �  �� �� ۽ }� �wv
��皪���   �   �   w   �   v   p         �  ��  ��  �� �} ��w���������  ̽  �� "�w"����vv� �|� ��    �  ��  ��  �� �� ������������  ��� ���"��|"�}l�wgl ~m� �}    �� �� ͼ �� ʧݼ��w���~�����   ��  ��  �p  }`  g`  m�  }�  �   �   �   �   Ȩ�������                   "   "   "          �  �  �  �  ʧ ��� ��� �����  ��� ��� ��p �}` wg` ~w  �   ˚  �   �                      w`                                �� ���˙�̻�� �� �̰ ��  ��  ��  �P  ��                  ���w��� ��� �̚ �I��˴��  L�    �   �     ��  [�  %�  "�      �� ��  ��  �   �   �   �       p                               ����                             �                              �� �̽ ��� ۽w }�� wvv��uP �� ����                                                            w��"���"��            ���"���"����                          �    "
��"��"�                                               �p    
�� �� �                ��  [�  %�  "�                   �� �̽ ���۽w�}�֪wvv���p��  �   �   �   �                                               ˚� ̹���ˈ�����̻����ۼ̼���˻                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            """ "!   " ""  !"""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  "" "  """ "!  "" "  """           """                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                                       """ "!   " ""  !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                         ��  vv  w                                 �  �  "  �  �     �  �     � � �  �       ڪ��z���
��̚���ɛ������������۸	�݉���˽X���� E�  E�  UX  �   �   
  �� ��� �� ��           �   �   ̰  ̸  ˉ  ��  �E  �T0 �T0 �S3 EC3 T3=�T3�а=؀���� ��  "�""""�""!��!  ��                     �  �  �  w                �   ��  �ڛ�}ک�"   "   "  �� ��                   ����������             ��  �   ��  �                 �   ��  ��  ��  �  �   ��  ��      � �������������  �                                                                                                                                             �   �   �   }�  g�Ȫ��̚���ə��̻ ��� ��  ��  ��  �  I�  DD ED UT UD UD UD DD DL ��  ��  ��  �   "  " �"/��"�   ��  ݰ  w�  mp gp �ת�����ș��˻�˰��� ��� �˰ ̻  ��  ��  DD@ DEH DUH UX UD TD DD  DL ��  ��  ʠ  ,�  "   "" ""���/ "  "  "  ""  �+  ��  �   �     "� .  "+  "�  �  �   �   
      �   �   �        �     �  �           �   �   �                     �  �� �� ��                     ��  ��  ���                                                                                                                                                                                                                �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �        �  ��� ��� ��p �}`
wg`�ww   �   �  �  �  �   �  �  �   �  �                                                �          �       �                        �   ��  ���  � �    �                                ����                  �   �� �       �  �  ��  �   �   �   �                                                 �   �  �  �  ��  ��  C�  U=  UJ  DZ  D  E  �4 
�: ���+��"��""� """ ""   �   �                        ɪ��ɪw̚�p�������������˻��۽��ݸ�̲-ۻ"""�""�2"�@  �C  �D  �T  D@  �   �   �   "�  "     �� �  �                                        ܰ ˻ �ݚ��w{`  g`  w                      �  �  ��"� ��� "                     �        �   �     �       �   �   �   �   �      �                    ��� ���� ��  ���� �                                                                                                                                                                                          �  �� �� wȠm���g���'�̹w ��� ��  ��  ��  ��  ��  ��  I�  C� C3 C4 D4 D4 � ��  ��  ��  �  "  "" �"!"/� �"   "�   ��  ��" {�" }�" wr",z��+�������ݻ���˻� ˼� ��  ˼  ��  ��  ��� DH� DX� D�@ E�  U�  E�  D�  ˸  ��  ��  ,�  ""  ""� ""� !�� � ��                                    �   �   �        "  "  "  ",  "�  �   �   �                 � �� �  �   �   �           �   �   �           �  ��  �                                                                                                                                                                                                                      �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��               �   �   �  �  �  �  �   �   �                                       �  ���          "   "   "                                �   �      ��   �  ��  �  �  �         � �������������  �                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                      �  �� ��  �    � ���                                                                                                                                                                                             	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����            ����  �  �  �  �  ��  �                      � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                        �  ��� ݼ� wۺ�m}ڪggz�p�� 
�� 
�� ��� ��� ˝� ɭ� ʝ ��- ��# �#$ " 8 "$� "���� ��  �        �"��""    ��                       ��  ��� ��� ��� ��� ��� ��� ��� ��ɀ�̔@���@��E@H�T@�TD �D@ DC� C3� �:� �� �"" �"" "�"��"� ��� ��  ��                  ������� ���        T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ���� ��� ����                � ��                    ���� �                                           �   ���                            �   �                                                                                                                 �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �             � ����  �                           �                        ���� ��� ����                                    � �� �  �  �   �   ��  �                            �   ���                            �   �                                                                                                          �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ�����ٺ�����؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� �����  ��� ��  �                                        �� ��                  �          �         �   �  �  �   �               �   �                     �                                                                                                                                                                                                     �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                            @  A   �  D   D                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwwwwwqwwwwDwwG""""wwwwqqAqDAqwqwq""""wwwwwqGAAA""""wwwwwqDDGwDww""""wwwwwwwqqDqG""""wwwwwqDDDG""""wwwwwwwwwAwwwGwwGw""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD��M����������������3333DDDD��A�����A�DMD�����3333DDDDAAMM�D�M�����3333DDDD����DMMDD�M����3333DDDDAMA�����D������3333DDDD�M���DD������3333DDDD�M��M�M�D��DM������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""����������D��M��M""""����������""""�����ADMA����""""����DD�M�""""��������AD�DM�""""�����������A�A�""""������AD�������""""������������������������"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��M��M�������D����3333DDDD�DD�M�D�������3333DDDDD�������M�DM�D����3333DDDD��A�M�M���M�����3333DDDDMM������D��D����3333DDDDA�A�A�D��M�D�����3333DDDD�������������D������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`����������������  `  V    a b c d e f g h i j i i i j i ij i i ij i i ij ihgfedcb(a(((V((`���������������� 
 M k +  l m b n o p q r s t u v u u u v u uv u u uv u u uv utsrqponbml((+(k(M 
���������������� w x M 5 6 y b n z { | } ~  � � � � � � � � �� � � �� � � �� �� � �|{znby(6(5(Mxw���������������� w w x 
 � b � � � � � � � � � � � � � � � � �� � � � � � � � � � � � � � �����b(� 
xww���������������� + � w w � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ����� ��ww�(+���������������� � W  � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � ������ ���((W(����������������� � a � l � � � � � �������� � � � � � � ���������� � � �� �������l(�(a(����������������� �  � y � � � � � � � � � � � � � � � ��� � � ������ � � � � � � � � ������y(�(����������������� = l �  � � � � � � � � � � ��� � � � ��� � ����� � � � ��� � � � ������((�l(=����������������    �  � � � � � � � � � ������ � � � � ����� � � � ������ � � �����((�(( ���������������� x X 5 - � � � � � � � � � � � � � ��� � � � ��� � � � � � � � � � ��� � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����(�xww����������������  � w w � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �����ww�(���������������� �  + � � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� ������(+((����������������� ` m � W � � � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� �����(W(�m(`���������������� M   a � � � � � ��� � � � � � ��� � � � � � � � ��� � � � � � ��� � �� ���(a((M���������������� � 
 � - � � � � � � ����� ���� � � � � � � � � � ����� ���� � � � � ���(-(� 
(����������������� � -    � � � � � � � � ����� � � � � � � � � � � � � � ����� � � � � � ����(( (-(����������������� 5 6  X � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � � � ���(X((6(5���������������� x �  l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���l((�x���������������� w w � � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq7c� �Oc� �%Kb K"_%K#Zkj_6 kr_ �B� � 	B� � 
B� � � B� � � B� � B� �K � �K � �C. � � C6 � �C7 � �C9 � � C; � �
B�1 �B�0 � B�I � B�) �cV � � c^ � �
c� � � c� � c� �c�p � c�h �	 �
 �	!�! �"� �#�3$"� %"�&"� �'*�Z("� �Z )"� �J*� �J+
� � � ,"O z  "& r  "& r �/": r � 0"A z � 1"P z �  " r � 3"O z � 4"K z � !� r � !� r z7"  r � 8"O z � 9"K z � !� r  "& r � <"O z  "& r �>!� r � "< r3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������ �!����������������������������������������������������������"�#�j�k�&�'�(����������������������������������������������������������)�*�l�m�n�.�/����������������������������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E�������������������������������������������������������������������������������������������������������������������������������������1�G�S�K���\�K�X���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �����������������������������������������"��4�K�X�K�S�_��;�U�K�T�O�I�Q� � � � � � �-�2�3�����������������������������������������$��<�Z�K�\�K��B�`�K�X�S�G�T� � � � � � � �.�/�=�������������������������������������������-�N�X�O�Y�Z�G�T��;�[�[�Z�Z�[� � � � � �-�2�3�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������.�/�=� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������-�2�3� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                