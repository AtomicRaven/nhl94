GST@�                                                           �o�                                                      R���      �  ��           ���2�������J�����������h�������        �g     #    ����                                d8<n    �  ?     B����  �
fD�
�L���"����D"��   " `  J  jF��    "�j "����
��
��     �j�� 
   ��
  �                                                                               ����������������������������������      ��    bb QQb  114 44c c   c         		 

       	   
       ��G �   ( (                 nnn ))1         888�����������������������������������������������������������������������������������������������������������������������������?=  00  54  81                        
     
                ��  4�  �  ��                  YE            : �����������������������������������������������������������������������������                                   3       �   @  &   �   �                                                                                 '       )n)n1n  YE    ��   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� IE 3 �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������     ��A^��AS|]�aA��zZ��V�Ph,D�|�s �v3��T0 k� ����Í&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��zZ��VTi,D�|�s �v3��T0 k� ����Ì&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��zZ��VXj,D�|�s �u3��T0 k� �Ì�ǌ&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��zZ��V\k,D�{�s �u3��T0 k� �Ì�ǌ&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��zZ��V`k,D�{�s �u3��T0 k� �ǋ�ˋ&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��zZ��Vdl,@�{�s �u3��T0 k� �ǋ�ˋ&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��zZ��Vhm,@�{�s �u3��T0 k� �ˊ�ϊ&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��zZ��Vln,@�z�s �u3��T0 k� �ˊ�ϊ&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��zZ��Vpo,@�z�s �u3��T0 k� �ω�Ӊ&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��zZ��V�to,@�z�s �u3��T0 k� �ω�Ӊ&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��zZ��V�|p,@�yxs �u3��T0 k� �Ӊ�׉&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��{Z��V��q,@,y�ps �u3��T0 k� �ӈ�׈&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��{Z��V��q,@,y�hs �u3��T0 k� �׈�ۈ&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��{Z��V��r,@,y�`s �t3��T0 k� �׈�ۈ&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��{Z��V��r,@,y�Xs �t3��T0 k� �ۇ�߇&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��{Z��V��s,@,y�Ps �t3��T0 k� �ۇ�߇&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��{Z��V��s,@ y�Hr �t3��T0 k� �߇��&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��{Z��V��s,@ y�@r �t3��T0 k� �߆��&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��{Z��V��t,@ y�8r�t3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��{Z��V��t,@ x�0r�t3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��{Z��V��t,@ x�(r�t3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��{Z��V��t,@Lx� r�t3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��{Z��V|�t,@Lx�r�t3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��{Z��V|�t,@Lx�r�t3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��{Z��V|�t,@Lx�r��t3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��V|�t,@Lx� r�|t3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��V|�t,@�w��r�xt3��T0 k� �����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��V|�s,@�w��r�tt3��T0 k� �����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��V|�s,@�w��r�ps3��T0 k� �����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��V|�s,@�v��r�ls3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��V|�r,@�v��r�hs3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��V|�r@�u��r�ds3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��V|�q@� u��r�`s3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��Vl�q@� t��r�Xs3��T0 k� �����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��Vl�p@�$t�r�Ts3��T0 k� �����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�bA��|Z��Vm o@�$s�r�Ps3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�bA��|Z��Vmo@�(r�r�Hs3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�bA��|Z��Vmn\@�,r�r�Ds3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�bA��|Z��Vmm\@�0q�r�@s3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��|Z��Vml\@�0p�r�8s3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��|Z��Vmk\@�4p�r�4s3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��|Z��Vmk\@�8o�r�,s3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��Vmj\@�<o|r�(s3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��Vmi\@�@ntr� s3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��V]h\@�Dmlr�s3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��V]g\@�Hmdr�s3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��V] f\@�Ll\r�s3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��V] e\@�TlTr s3��T0 k� ��&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��V] d\@�XkLr  r3��T0 k� ��&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��V] c\@�\kDr�r3��T0 k� ��&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��V]$c\<�`j<r�r3��T0 k� ��&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��V]$b\<�hi4r�r3��T0 k� ��#&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��ASx]�cA��}Z��V�$a\<�li,r�r3��T0 k� ��#&�1D"3Q	2�4#Q  ��_    � +�8 ��A^�ASx]�cA��}Z��V� `\<�ph$r�r3��T0 k� ��#&�1D"3Q	2�4#Q  ��_    � +�8 ��A^�ASx]�cA��}Z��V� _\<�xgq�r3��T0 k� �#~�'~&�1D"3Q	2�4#Q  ��_    � +�8 ��A^�ASx]�cA��}Z��V� _\<�|gq�r3��T0 k� �#~�'~&�1D"3Q	2�4#Q  ��_    � +�8 ��A^�ASx]�cA��}Z��V� ^\<��f�q�r3��T0 k� �'~�+~&�1D"3Q	2�4#Q  ��_    � +�8 ��A^�ASx]�cA��}Z��V ]\<��e�r�r3��T0 k� �'~�+~&�1D"3Q	2�4#Q  ��_    � +�8 ��A^�ASx]�bA��}Z��V \\<��d�r�r3��T0 k� �'~�+~&�1D"3Q	2�4#Q  ��_    � +�8 ��A^�ASx]�bA��}Z��V \\<ܔc� s�r3��T0 k� �+~�/~&�1D"3Q	2�4#Q  ��_    � +�8 ��A^�ASx]�bA��}Z��V[\<ܜb��s�r3��T0 k� �+~�/~&�1D"3Q	2�4#Q  ��_    � +�8s�eR�#�D�S�T6B��Y|/����r�q	#��W�#����T0 k� �k��o�&�1D"3Q	2�4#Q  ��    ��� s�dR�#�D�_�\7B���Y|/����r�q	#��_�#����T0 k� �w��{�&�1D"3Q	2�4#Q  ��    ��� s�cR�#�D�g�d7B���Y|/����r�p c��g�#����T0 k� ���&�1D"3Q	2�4#Q  ��    ��� s�bR�#�D�s�l7B��Y|/����r�p c��o�#����T0 k� ��~��~&�1D"3Q	2�4#Q  ��    ��� s�bR�#�D�{��t8B��Y|/����r�o c��w�#����T0 k� ��~��~&�1D"3Q	2�4#Q  ��    ��� s�aR�#�O����|8B��Y|/����r�n c��������T0 k� ��~��~&�1D"3Q	2�4#Q  ��    ��� s�`R��O�����8B��Y|/����r�m c���������T0 k� ��~��~&�1D"3Q	2�4#Q  ��   ��� s�^R��O�����9B�+�Y|/�q��r�l c���������T0 k� ��~��~&�1D"3Q	2�4#Q  ��    ��� ��]R��O�����9B�3�Y|/�q��b�k ����������T0 k� ��~��~&�1D"3Q	2�4#Q  ��    ��� ��[R��O�����9B�;�Y|/�q��c j ����������T0 k� ��~��~&�1D"3Q	2�4#Q  ��    ��� ��ZR��O�����9B�C�Y|/�q��ci ����������T0 k� ��~��~&�1D"3Q	2�4#Q  ��    ��� ��YR��O�����9B�K�Y|/�r�ch ����������T0 k� ����&�1D"3Q	2�4#Q  ��    ��� �XR��O�����9B�S�Y|/�r�cg ����������T0 k� ����&�1D"3Q	2�4#Q  ��    ��� �UR��O�����9B�c�Y|/�r�ce��ϗ�����T0 k� ����&�1D"3Q	2�4#Q  ��    ��� �TR��O�����9B�k�Y|/�r#�c d��חC����T0 k� ����&�1D"3Q	2�4#Q  ��    ��� �RR��O���p�9B�s�Y|/�r+�c$c��ۘC����T0 k� ����&�1D"3Q	2�4#Q  ��    ��� �$QR��O���p�9B�{�Y|/�r3�c(b���C����T0 k� ������&�1D"3Q	2�4#Q  ��    ��� �,OR��O��p�9Bރ�Y|/�r;�c,a���C����T0 k� �����&�1D"3Q	2�4#Q  ��    ��� �0NR��O��p�9B���Y|/�bC�S0`S�C�C����T0 k� ����&�1D"3Q	2�4#Q  ��    ��� �<KR��O��q8B���Y|/�bS�S8]S�C��C�"���T0 k� ����&�1D"3Q	2�4#Q  ��    ��� �@IR��O���8B���Y|/�b[�S<\S�D�C�"��T0 k� ����&�1D"3Q	2�4#Q  ��    ��� �HHR��O���7B���Y|/�bc�S<[S�D�C�"��T0 k� ���#�&�1D"3Q	2�4#Q  ��    ��� �LFR��O�'�� 7B���Y|/�bg��@Z��D�C�"��T0 k� �'��+�&�1D"3Q	2�4#Q  ��    ��� �TDR��O�/��(7B���Y|/�bo��DY��D�C�"��T0 k� �+��/�&�1D"3Q	2�4#Q  ��    ��� �\AR��O�;��85B���Y|/�b{��HW��D#�C�"��T0 k� �7��;�&�1D"3Q	2�4#Q  ��    ��� �d?R��E�C��@5B���Y|/�2��HV���D+���"��T0 k� �?��C�&�1D"3Q	2�4#Q  ��    ��� �h>R��E�K��D4B���Y|/�2���HU���D/���"��T0 k� �C��G�&�1D"3Q	2�4#Q  ��    ��� �l<R��E�K��L3B���Y|/�2���LT���D7���"��T0 k� �K��O�&�1D"3Q	2�4#Q  ��    ��� �t:R��E�O��T3B���Y|/�2���LS����;�����T0 k� �K��O�&�1D"3Q	2�4#Q  ��    ��� �|7R��E�[��`1B���Y|/�2���LQ����C�����T0 k� �S��W�&�1D"3Q	2�4#Q  ��    ��� ��5R��Erc��h0B���Y|/�2���LQ����G�����T0 k� �W��[�&�1D"3Q	2�4#Q  ��    ��� ��3R��Erg��l/B��Y|/�2���LP����G�����T0 k� �W��[�&�1D"3Q	2�4#Q  ��    ��� ��0R��Erg��|-I�Y|/�2���LN����O�����T0 k� �_��c�&�1D"3Q	2�4#Q  ��)    ��� ��.R��Erk���,I�Y|/�b���LM����O�����T0 k� �_��c�&�1D"3Q	2�4#Q  ��)    ��� ��,R��E�o�q�+I#�Y|/�b���HL����S�����T0 k� �c��g�&�1D"3Q	2�4#Q  ��)    ��� ��*R��E�s�q�*I'�Y|/�b���HK���tW�����T0 k� �g��k�&�1D"3Q	2�4#Q  ��)    ��� ��'R��E��q�'I/3�Y|/�b���DJ���t[�����T0 k� �k��o�&�1D"3Q	2�4#Q  ��)    ��� ��%R��E��q�&I/;�Y|/�b���DI���t[���"��T0 k� �k��o�&�1D"3Q	2�4#Q  ��)    ��� ��#R��F��q�%I/?�Y|/�b���@H��t_�	s�"��T0 k� �k��o�&�1D"3Q	2�4#Q  ��)    ��� ��!R��F��q�#I/C�Y|/�b��@G��tc�	s�"��T0 k� �o��s�&�1D"3Q	2�4#Q  ��)    ��� ��R��F��q� IO�Y|/�b��<F��tg�	s�"��T0 k� �s��w�&�1D"3Q	2�4#Q  ��)    ��� ��R��F��a�IS�Y|/�b��8E��tg�	s�"��T0 k� �s��w�&�1D"3Q	2�4#Q  ��)    ��� ��R��F��a�IW�Y|/�R��4D��tk�	��"��T0 k� �w��{�&�1D"3Q	2�4#Q  ��)    ��� ��R��F��a�I[�Y|/�R��0C��tk�	� "��T0 k� �w��{�&�1D"3Q	2�4#Q  ��)    ��� ���R��F��a�I/g�Y|/�R��(B��do�	�"��T0 k� �k��o�&�1D"3Q	2�4#Q  ��)    ��� ���R��E���a�I/k�Y|/�R��(A��do�	�"��T0 k� �_��c�&�1D"3Q	2�4#Q  �)    ��� ���R��E���a�I/k�Y|/�R��$@{�ds�	s��T0 k� �S��W�&�1D"3Q	2�4#Q  ��/    ��� ���R��E���a�I/o�Y|/�R��@�w�ds�	s��T0 k� �C��G�&�1D"3Q	2�4#Q  ��/    ��� ���R��E���a�Iw�Y|/�R��>�g�dw�	s��T0 k� �+��/�&�1D"3Q	2�4#Q  ��/    ��� ���R��E�����I{�Y|/�R��>�_�$w�	s��T0 k� ���#�&�1D"3Q	2�4#Q ��/    ��� �	ԄR��E�����I�Y|/�R��=�S�${�	�	��T0 k� ����&�1D"3Q	2�4#Q ��/    ��� �	ԄR��E�����I�Y|/�R��<�K�${�	�
��T0 k� ����&�1D"3Q	2�4#Q ��/    ��� �	Ԅ R��E����
I��Y|/�R�� <�C�${�	�
��T0 k� ������&�1D"3Q	2�4#Q ��/    ��� �	ԇ�R��E���I/��Y|/�R���:�3��	���T0 k� �۪�ߪ&�1D"3Q	2�4#Q ��/    ��� �	ԇ�R��E���I/��Y|/�R���:�3���	s��T0 k� �Ϭ�Ӭ&�1D"3Q	2�4#Q ��/    ��� �	��R��E���I/��Y|/�R���9�/���	s��T0 k� �í�ǭ&�1D"3Q	2�4#Q  ��/    ��� �	��R��E���I/��Y|/�S��8�/���	s��T0 k� ������&�1D"3Q	2�4#Q  ��/    ��� �	��R��E#���I/��Y|/�S���8�+���	s��T0 k� ������&�1D"3Q	2�4#Q  ��/    ��� �	��R��E7��� B���Y|/�S���7�'���	���T0 k� ������&�1D"3Q	2�4#Q  ��/    ��� �	ԇ�R��E�?����B���Y|/�S���6�'���	���T0 k� ������&�1D"3Q	2�4#Q  ��/    ��� �	ԇ�R��E�G����B���Y|/�S���5�'���	���T0 k� �s��w�&�1D"3Q	2�4#Q  ��/    ��� �	ԇ�R��E�O����B���Y|/�S��5�'���	���T0 k� �g��k�&�1D"3Q	2�4#Q  ��/    ��� �	ԇ�R��E�[�a��B���Y|/�S��4�#���	�d�T0 k� �[��_�&�1D"3Q	2�4#Q  ��/    ��� �	ԇ�R��E�c�a��B���Y|/�S��4����	sd�T0 k� �O��S�&�1D"3Q	2�4#Q  ��/    ��� �	��R��E�k�a��B���Y|/�S��3����	sc��T0 k� �?��C�&�1D"3Q	2�4#Q  ��/    ��� �	��R��E�w�a��B���Y|/�S��3����	sc��T0 k� �3��7�&�1D"3Q	2�4#Q  ��/    ��� �	��R��E��a��B���Y|/�S��2����	sc��T0 k� �'��+�&�1D"3Q	2�4#Q  ��/    ��� |	��R��E���a��B���Y|/����1����	�c��T0 k� ����&�1D"3Q	2�4#Q  ��/    ��� w	ԇ�R��E���a��B���Y|/����1����	�c��T0 k� ����&�1D"3Q	2�4#Q  ��/    ��� x	ԇ�R��E���a��B���Y|/����|0����	�c��T0 k� ������&�1D"3Q	2�4#Q  ��&    ��� y	ԇ�R��E���Q��B���Y|/����t0����	�c��T0 k� ������&�1D"3Q	2�4#Q  ��&    ��� z	ԇ�R��E���Q��B���Y|/����l/r���	�c��T0 k� ������&�1D"3Q	2�4#Q  �&    ��� {	ԇ�R��QS��Q��B���Y|/�c��X.r���Sc��T0 k� �׽�۽&�1D"3Q	2�4#Q  ��&    ��� |	��R��QS��Q��B���Y|/�c��P.q��4��Sc��T0 k� �ϻ�ӻ&�1D"3Q	2�4#Q  ��&    ��� }	��R��QS��Q��B���Y|/�c��H-q��4��Sc��T0 k� �Ǻ�˺&�1D"3Q	2�4#Q  ��&    ��� }	��R��QS��Q��B���Y|/�c��@-a��4��Sc��T0 k� �ù�ǹ&�1D"3Q	2�4#Q  ��&    ��� }	��R��QS��Q��I��Y|/�c��8-a��4��Sc��T0 k� ����ø&�1D"3Q	2�4#Q  ��&    ��� }	��R��QS����I��Y|/�c��0,a��4���c��T0 k� ������&�1D"3Q	2�4#Q  ��&    ��� }	ԇ�R��QS����I��Y|/�c� +a��4���c��T0 k� ������&�1D"3Q	2�4#Q  ��&    ��� }	ԇ�R��Qc����I��Y|/�c�+a��4���c��T0 k� ������&�1D"3Q	2�4#Q  ��&    ��� }	ԇ�R��Qc����I��Y|/�s�*a��4���c��T0 k� ������&�1D"3Q	2�4#Q  ��&    ��� }	ԇ�R��Qc����I/��Y|/�r��*a��4���c��T0 k� ������&�1D"3Q	2�4#Q  ��&    ��� }	ԇ�R��Qc����I/��Y|/�r���*a��4���c��T0 k� ������&�1D"3Q	2�4#Q  ��&    ��� |D��R��Qc���w�I �Y|/�r���)a��4���c��T0 k� ������&�1D"3Q	2�4#Q  ��&    ��� {D��R��Qc���s�I �Y|/�r�Q�)a��D���c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� zD��R��Qc��Qk�I �Y|/�r�Q�(Q��D���c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� yD��R��Qs��Qg�I�Y|/�R�Q�(Q��D��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� xD��R��Qs��Q_�I�Y|/�R�Q�(Q��D��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� w ��R��Qs��QS�I�Y|/�R߮Q�'Q��Dw��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� v ��R��Qs��QK�I�Y|/�RۮQ�'Q��Dw��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� u ��R��Qs��QC�I �Y|/�R׭Q�&Q��Ds��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� s ��R��Qs��Q;�I �Y|/�RϭQ�&Q��Do��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� q ��R��Qs��Q7�I �Y|/�RˬQ�&Q��Dk��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� o d��R��Qs� Q/�I �Y|/�RëQ�%Q��Dg��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� m d��S�Qs� Q'�I �Y|/�R��A�%Q��dg��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� k d��S�Qs�A�I#�Y|/�R��A�%A��dc��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� i d��S�Qs�A�I#�Y|/�B��A|$A��d_��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� g d��S�Qs�A�I#�Y|/�B��At$A��d[��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� eD��S�Qs�A�I#�Y|/�B��Al$A��dW��c��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� cD��S�Qs�@��I'�Y|/�B��A\$A�dO�� c��T0 k� �{���&�1D"3Q	2�4#Q  ��6    ��� aD��S�Qs�@��I '�Y|/�B��AT$Aw�dK�� c��T0 k� �s��w�&�1D"3Q	2�4#Q  ��6    ��� _D�S�Qs�@��I '�Y|/�B��AH$Ao�dG��$c��T0 k� �k��o�&�1D"3Q	2�4#Q  ��6    ��� ]D�U��Qs�@��I '�Y|/�B��A@$Ak�TC��$c��T0 k� �c��g�&�1D"3Q	2�4#Q  ��6    ��� [��U��Qs����I '�Y|/�B�A8$Ac�T;��$c��T0 k� �_��c�&�1D"3Q	2�4#Q  ��6    ��� Y��U��Qs����I '�Y|/�w�A0$A[�T7��(c��T0 k� �O��S�&�1D"3Q	2�4#Q  ��6    ��� W��U��Qs����@`'�Y|/�s�1($AW�T3��(c��T0 k� �C��G�&�1D"3Q	2�4#Q  ��6    ��� U�{�U��Qs����@`'�Y|/�k�1 $1O�T/��,c��T0 k� �;��?�&�1D"3Q	2�4#Q  ��6    ��� S�{�U��Qs����@`'�Y|/�c�1$1G��'��0c��T0 k� �/��3�&�1D"3Q	2�4#Q  ��6    ��� Q�{�U��Qs�@��@`'�Y|/�[�1$1C��#��0c��T0 k� �#��'�&�1D"3Q	2�4#Q  ��6    ��� O�w�U��Qs�@��@`'�Y|/�W�1%1;����4c��T0 k� ����&�1D"3Q	2�4#Q  ��6    ��� M�w�U��Qs�@��@�'�Y|/�O���%17����8c��T0 k� ����&�1D"3Q	2�4#Q  ��6    ��� K�w�U��Qs�@��@�'�Y|/�G���%A/����8c��T0 k� ����&�1D"3Q	2�4#Q  ��6    ��� I�s�A��Qs�@��@�'�Y|/�?���&A+����<c��T0 k� ����&�1D"3Q	2�4#Q  ��6    ��� G�o�A��Qs�	@�@�'�Y|/�/���&A�����Dc��T0 k� ������&�1D"3Q	2�4#Q  ��6    ��� E�o�A��Qs�	0w�@�'�Y|/�+���'A�����Hc��T0 k� ����&�1D"3Q	2�4#Q  ��6    ��� C�k�A��Qs�	0o�@�'�Y|/�"#���'A����Lc��T0 k� ����&�1D"3Q	2�4#Q  ��6    ��� A�k�Es�Qs�
0g�A '�Y|/�"���(A����Pc��T0 k� ����&�1D"3Q	2�4#Q  ��6    ��� ?�k�Es�Qs�
0g�A #�Y|/�"���(A����Tc��T0 k� �߻��&�1D"3Q	2�4#Q  ��6    ��� =�g�Es�Qs�
0g�A �Y|/�"���)A��ߵ�Xc��T0 k� �׼�ۼ&�1D"3Q	2�4#Q  ��6    ��� :�g�Es�Qs�0c�A �Y|/�"���)@��S۵�\c��T0 k� �ϼ�Ӽ&�1D"3Q	2�4#Q  ��6    ��� 8�g�Es�Qs�0_�A �Y|/�!����*P��SӴ�`c��T0 k� �ǽ�˽&�1D"3Q	2�4#Q  ��6    ��� 6�g�Ec�Qs�0[�E��Y|/�!���*P�S˴�`c��T0 k� ������&�1D"3Q	2�4#Q  �6    ��� 1�g�Ec�Qs� [�E��Y|/�a���+P�Só�dc��T0 k� ������&�1D"3Q	2�4#Q ��?    ��� ,�c�Ec�Qs� W�E��Y|/�a���+P�S���hc��T0 k� ������&�1D"3Q	2�4#Q ��?    ��� '�c�Ec�Qs� S�E��Y|/�a۰��,P�S���h3��T0 k� ������&�1D"3Q	2�4#Q ��?    ��� "�c�Ec�Qs� S�E��Y|/�aӱ�x,0۪S���l3��T0 k� ������&�1D"3Q	2�4#Q ��?    ��� �c�C��Qs� O�E��Y|/�a˱�p-0׫C���p3��T0 k� �{���&�1D"3Q	2�4#Q ��?    ��� �_�C��Qs��O�E���Y|/�aò�h-0ӬC���p3��T0 k� �o��s�&�1D"3Q	2�4#Q ��?    ��� �_�C��Qs��K�E���a�/�q���`.0ϬC���p3��T0 k� �_��c�&�1D"3Q	2�4#Q ��?    ��� �[�C��Qs��K�E���a�/�q���T.0˭C���t3��T0 k� �S��W�&�1D"3Q	2�4#Q ��?    ��� 	�[�C��Qs��G�E���a�/�q���L/0ǮC���t3��T0 k� �G��K�&�1D"3Q	2�4#Q ��?    ��� �W�C��Qs��G�Eo��a�/�q���D00��C��t3��T0 k� �;��?�&�1D"3Q	2�4#Q ��?    ��� �S�C��Qs� G�Eo��a�/�q���<0 ��Cw��x3��T0 k� �/��3�&�1D"3Q	2�4#Q ��?    ������S�C���Qs� G�Eo��a�/�����41 ��Co��x3��T0 k� ���#�&�1D"3Q	2�4#Q ��?    ������O�C���Qs� C�Eo��a�/�����,1 ��Cg��x3��T0 k� ����&�1D"3Q	2�4#Q ��?    ������K�C���Qs� C�Eo��a�/�����$2 ��C_��x3��T0 k� ����&�1D"3Q	2�4#Q ��?    ������G�C��Qs� C�E���a�/�����2 ��CW��x3��T0 k� ������&�1D"3Q	2�4#Q ��?    ������G�C��Qs�C�E���a�/�����3 ��3S��x3��T0 k� ������&�1D"3Q	2�4#Q ��?    ������C�C��Qs�C�E���a�/��{��3 ��3K��x3��T0 k� ������&�1D"3Q	2�4#Q ��?    ������?�C��Qs�G�E���Y|/��w��4 ��3C��x3��T0 k� ������&�1D"3Q	2�4#Q	 ��?    ������;�C��Qs�G�E���Y|/��s���4 ��3;��x3��T0 k� ������&�1D"3Q	2�4#Q	 ��?    ������7�C�ۯQs�G�E���Y|/��k���5 ��33��x3��T0 k� ������&�1D"3Q	2�4#Q	 ��?    ������/�C�ׯQs��G�F��Y|/��g���5���3+��x3��T0 k� ������&�1D"3Q	2�4#Q	 ��?    ������+�C�ӰQs��K�F��Y|/��_���6���3'��x3��T0 k� ������&�1D"3Q	2�4#Q	 ��?    ������'�C�ϰQs��K�F��Y|/��[���6���3��x3��T0 k� ������&�1D"3Q	2�4#Q	 ��?    ������#�C�ǱQs��K�F��Y|/��W���7���3��x3��T0 k� ������&�1D"3Q	2�4#Q	 ��?    �������C�òQs��O�F��Y|/��O���8���3��x3��T0 k� �{���&�1D"3Q	2�4#Q	 ��?    ������C�Qs��O�D߻�Y|/��K���8���#��x3��T0 k� �o��s�&�1D"3Q	2�4#Q	 ��?    ������D��Qs��O�D߻�Y|/��G�ϼ9���#��x3��T0 k� �c��g�&�1D"3Q	2�4#Q	 ��?    ������D��Qs��S�D߷�Y|/��?�ϴ9���"���x3��T0 k� �W��[�&�1D"3Q	2�4#Q	 ��?    ������D��Qs��S�D߷�a�/��;�Ϭ:���"���x3��T0 k� �G��K�&�1D"3Q	2�4#Q	 ��?    ������D��Qs��W�D߷�a�/��7�Ϥ:���"��x3��T0 k� �;��?�&�1D"3Q	2�4#Q	 ��?    �������D��Qs��W�D߳�a�/��3�Ϝ;���"��x3��T0 k� �/��3�&�1D"3Q	2�4#Q	 ��?    �������D��Qs��W�D߳�a�/��+�ϔ;���"��x3��T0 k� � �$&�1D"3Q	2�4#Q	 ��?    �������D��Qs��W�E���a�/��'�ό<���"��x3��T0 k� ��&�1D"3Q	2�4#Q	 ��?    �������D��Qs��W�E���a�/��#�τ<���"ߵ�x3��T0 k� ��&�1D"3Q	2�4#Q	 ��?    �������D�Qs��[�E���a�/����|=���"۶�x3��T0 k� ����&�1D"3Q	2�4#Q ��?    �������Dw�Qs��[�E���a�/����t=���"׷�x3��T0 k� ��	��	&�1D"3Q	2�4#Q ��?    �������Ds�Qs��[�E���a�/����l>���ӷ�x
3��T0 k� ����&�1D"3Q	2�4#Q ��?    �������Dk�Qs��[�E��a�/����d>���ϸ�x
3��T0 k� ����&�1D"3Q	2�4#Q ��?    �������Dc�Qs��[�E��a�/����\?���˹�x
3��T0 k� ����&�1D"3Q	2�4#Q ��?    �������D[�Qs��[�E��Y|/����X?���˹�x
3��T0 k� ����&�1D"3Q	2�4#Q ��?    �������DS�Qs��[�E��Y|/�����P@���Ǻ�x
3��T0 k� ����&�1D"3Q	2�4#Q ��?    �������DK�Qs��[�E��Y|/�����H@���û�x
3��T0 k� ����&�1D"3Q	2�4#Q ��?    �������DC�Qs��[�E��Y|/�����@A����ü�x
3��T0 k� ����&�1D"3Q	2�4#Q ��?    �������D;�Qs��[�E��Y|/�����8A�������x
3��T0 k� ����&�1D"3Q	2�4#Q ��?    �������D/�Qs��[�E��Y|/�����0B�������x
3��T0 k� �x�|&�1D"3Q	2�4#Q ��?    �������D'�Qs��_�E��Y|, ����$B�������x
3��T0 k� �l�p&�1D"3Q	2�4#Q ��?    �������D�Qs��_�E��Y|, ����C�������x
3��T0 k� �` �d &�1D"3Q	2�4#Q ��?    ����}��D�Qs��_�E��Y|, ����C�������x
3��T0 k� �T"�X"&�1D"3Q	2�4#Q ��O    ����z�{�C��Qs��[�E��Y|,����D������Cx
3��T0 k� �H$�L$&�1D"3Q	2�4#Q ��O    ����w�s�C��Qs��[�E��Y|,����D������Cx
3��T0 k� �<&�@&&�1D"3Q	2�4#Q ��O    ����t�k�C���Qs��[�Eo��Y|,л���E������Cx
3��T0 k� �,(�0(&�1D"3Q	2�4#Q  ��O    ����p�_�C���Qs��[�Eo��Y|,г���E������Cx
3��T0 k� � +�$+&�1D"3Q	2�4#Q  ��O    ����m�W�C��Qs��[�Eo��Y|,����FЗ����Cx
3��T0 k� �-�-&�1D"3Q	2�4#Q  ,�O    ����j�O�C��Qs��[�Eo��Y|,����FЗ���� x
3��T0 k� �/�/&�1D"3Q	2�4#Q  ��O    ����g�G�C�ۿQs��W�Eo��Y|,�����GЗ�B�� x
3��T0 k� ��1� 1&�1D"3Q	2�4#Q  ��O    ����d�?�C�ӿQs��W�Eo��Y|,�����GГ�B�� x
3��T0 k� ��3��3&�1D"3Q	2�4#Q  ��O    ����a�7�C�˿Qs��W�Eo��Y|,�����GГ�B�� x
3��T0 k� ��5��5&�1D"3Q	2�4#Q ��O    ����^�/�C���Qs��S�Eo��Y|,�����HЏ�B�� x
3��T0 k� ��7��7&�1D"3Q	2�4#Q ��O    ����[�#�C��Qs��S�Eo��Y|,�{�޸HЏ�B�� cx
3��T0 k� ��9��9&�1D"3Q	2�4#Q ��O    ����X��C��Qs��O�Eo��Y|,0s�ްIЋ�B�� cx
3��T0 k� ��;��;&�1D"3Q	2�4#Q ��O    ����V��C��Qs��O�Eo��Y|,0k�ިIЋ�B�� cx
3��T0 k� ��=��=&�1D"3Q	2�4#Q ��O    ����T��C��Qs��K�Eo��Y|,0c�ޠJЋ�B�� cx
3��T0 k� ��?��?&�1D"3Q	2�4#Q ��O    ����R��C��Q���G�Eo��Y|,0[��JЇ�B�� cx
3��T0 k� ��A��A&�1D"3Q	2�4#Q ��O    ����P���C��Q���D Eo��Y|,0S��JЃ�B��Cx
3��T0 k� ��C��C&�1D"3Q	2�4#Q ��O    ����N���C��Q���@Eo��Y|,0K��J��R��Cx
3��T0 k� �|E��E&�1D"3Q	2�4#Q ��O    ����L���C��Q���<E_��Y|,0C��|K�{�R��Cx3��T0 k� �pG�tG&�1D"3Q	2�4#Q ��O    �  �J���C�w�Q���8E_��Y|,P;��tK�w�R��Cx3��T0 k� �dI�hI&�1D"3Q	2�4#Q ��O    � �H���C�o�Q���4E_��Y|,P3��lK�s�R��Cx3��T0 k� �XK�\K&�1D"3Q	2�4#Q ��O    � �G���C�g�Q���0E_��Y|,P+��dK�o�R��Cx3��T0 k� �LM�PM&�1D"3Q	2�4#Q ��O    � �F���C�[�Q���,E_��Y|,P#��\K�h "��Cx3��T0 k� �@O�DO&�1D"3Q	2�4#Q ��O    � �E��C�S�Q���(
E_�Y|,P��PK�d"��Cx3��T0 k� �0Q�4Q&�1D"3Q	2�4#Q ��O    � 
�D��DK�U#��$E_{�Z�,P��HK�`"��Cx3��T0 k� �$S�(S&�1D"3Q	2�4#Q ��O    � �C��DC�U#�� E_t Z�,	P�>@KP\"��Cx3��T0 k� �U�U&�1D"3Q	2�4#Q ��O    � �B��D;�U#��E_pZ�,	_��>8KPX"��Cx3��T0 k� �W�W&�1D"3Q	2�4#Q ��O    � �A��D3�U#��E_lZ�,	_��>0KPP"��Sx3��T0 k� � Z�Z&�1D"3Q	2�4#Q  ��O    � �@��D+�U#��C�hZ�,
_��>(KPL"��Sx3��T0 k� ��\��\&�1D"3Q	2�4#Q  ��O    � �?��D#�U#��C�`Z�,
���> JPH��Sx3��T0 k� ��^��^&�1D"3Q	2�4#Q  ��O    � �>��D�U#��C�\Z�,
���>JP@	��Sx3��T0 k� ��`��`&�1D"3Q	2�4#Q  ��O    � �=��D�U#��C�XZ�,
���>JP<
��Sx3��T0 k� ��b��b&�1D"3Q	2�4#Q  /�O    � �<��D�U#�� C�T
Z�(���>JP4��Sx3��T0 k� ��d��d&�1D"3Q	2�4#Q  ��O    � �;��D ��@c���E�PZ�(���=�I�0��Sx3��T0 k� ��f��f&�1D"3Q	2�4#Q  ��O    � �:��D ��@c���E�HZ�(��=�I�("��Sx3��T0 k� ��h��h&�1D"3Q	2�4#Q  ��O    � �9��D��@c���E�DZ�(��=�I�$"��Sx3��T0 k� ��j��j&�1D"3Q	2�4#Q  ��O    �  �8��D��@c��E�@Z�(��=�H�"��Sx3��T0 k� ��l��l&�1D"3Q	2�4#Q  ��O    � !�8��D��@c��E�8Z�(��M�H�"��Sx3��T0 k� ��n��n&�1D"3Q	2�4#Q  ��O    � "�8��D��@���E�4Z�(��M�H�"��cx3��T0 k� �xp�|p&�1D"3Q	2�4#Q  ��O    � #�8{�D��@���E�0Z�$��M�G�"��cx3��T0 k� �lr�pr&�1D"3Q	2�4#Q  ��O    � $�8s�D��@���E�(Z�$��M�G� "��cx3��T0 k� �`t�dt&�1D"3Q	2�4#Q  ��_    � %�8Bk�D��@��� D?$Z�$��M�F����cx3��T0 k� �Pv�Tv&�1D"3Q	2�4#Q  ��_    � &�8Bg�D��@���!D? Z�$�w��F����cx3��T0 k� �Dx�Hx&�1D"3Q	2�4#Q  ��_    � '�8B_�D��A��"D?Z�$�o��E����cx3��T0 k� �8z�<z&�1D"3Q	2�4#Q  ��_    � (�8BW�D��A��#D?Z�$�g��E���cx 3��T0 k� �,|�0|&�1D"3Q	2�4#Q  ��_    � )�8BO�D��A��$D?Z�$�[��D���cx!3��T0 k� � ~�$~&�1D"3Q	2�4#Q  ��_    � *�8BK�C���A��%D?Z�(�S��D���	Sx#3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8BC�C���A��&D? Z�(�K��C���	Sx$3��T0 k� ����&�1D"3Q	2�4#Q  �_    � +�8B;�C��E���'A� !Z�(_C�m|C�� b�	Sx%3��T0 k� ���� �&�1D"3Q	2�4#Q  *�_    � +�8B3�C�w�E���(A��#Z�,_;�mtB�� b�		Sx&3��T0 k� �����&�1D"3Q	2�4#Q  -�_    � +�8B+�C�o�E���)A��$Z�,_3�mlA�� b�
	Sx(3��T0 k� ����&�1D"3Q	2�4#Q  ��_    � +�8'�APg�E���*A��&Z�,_+�mdA� b��x)3��T0 k� �؂�܂&�1D"3Q	2�4#Q  ��_    � +�8�AP_�E��_�+A��'Z�0_#�m\@� b��x*3��T0 k� �Ђ�Ԃ&�1D"3Q	2�4#Q  ��_    � +�8�APW�E��_x+A��(Z�4_�mT?����x,3��T0 k� �ā�ȁ&�1D"3Q	2�4#Q  ��_    � +�8�APO�E��_p,A��*Z�4_�mL?����x-3��T0 k� ̸����&�1D"3Q	2�4#Q  ��_    � +�8�APG�E��_l-A��+Z�8_�mD>����x.3��T0 k� ܬ����&�1D"3Q	2�4#Q ��_    � +�8�AP?�AS�_d.A��,Z�<^��m<=����x03��T0 k� ܠ����&�1D"3Q	2�4#Q ��_    � +�8��AP;�AS�_`/A��.Z�<^��]4<| ���x13��T0 k� ܔ��&�1D"3Q	2�4#Q ��_   � +�8��AP3�AS�_X0A��/Z�@N��],<x!���x23��T0 k� ܈��&�1D"3Q	2�4#Q ��_    � +�8��AP+�AS�_T0A��0a<@N��]$;p!���x33��T0 k� �|~��~&�1D"3Q	2�4#Q ��_    � +�8��AP#�AS�_L1A��1a<D N��]:h"���x43��T0 k� �p~�t~&�1D"3Q	2�4#Q ��_    � +�8��AP�AS�_H2A��2a<H!N��]:d#���x63��T0 k� �d}�h}&�1D"3Q	2�4#Q ��_    � +�8��AP�AS�_@3A��4a<H"N��9\#���x73��T0 k� �X}�\}&�1D"3Q	2�4#Q ��_    � +�8��AP�AS�_<4A��5a<L#N��8T$��!�x83��T0 k� �P|�T|&�1D"3Q	2�4#Q ��_    � +�8��AP�AS�_84A��6a<L%N���8P%��#�x93��T0 k� �D|�H|&�1D"3Q	2�4#Q  ��_    � +�8��AP�AS�_05A��7a<P&N���7/H%¬%�x:3��T0 k� �8{�<{&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�_,6A��8a<T'N���6/D&¬'�x;3��T0 k� �,{�0{&�1D"3Q	2�4#Q  ��_   � +�8��A_��AS�_(6A��9a<T(N���6/<&°)�x<3��T0 k� � z�$z&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�_ 7A��:a<X)����5/8'°+�x=3��T0 k� �z�z&�1D"3Q	2�4#Q  ��_   � +�8��A_��AS�_8A��;aLX*����5/0(°-�x>3��T0 k� �y�y&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�_8A��<aL\+����4/,(°/�x?3��T0 k� �y� y&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�_9A��=aL\,���4/$)´1�x@3��T0 k� �x��x&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�_:A��>aL`-�w��3/ )´3�xA3��T0 k� �x��x&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�_:A��?aL`.�k�,�2/*´5�xB3��T0 k� �w��w&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�_;A��@aLd/�c�,�2/*´7�xC3��T0 k� �w��w&�1D"3Q	2�4#Q  *�_    � +�8��A_��AS�_ <A��AaLd0�[�,�1/+Ҵ9�xD3��T0 k� ��u��u&�1D"3Q	2�4#Q  /�_    � +�8��A_��AS�^�<A��BaLh1�S�,�1/+Ҵ;�xE3��T0 k� ��s��s&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�^�=A��CaLh2�K�,�1/,Ҵ=�xF3��T0 k� �r��r&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�^�>A��DaLh3�C�,�1/ ,Ҵ>�xG3��T0 k� �p��p&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�^�>A��EaLh4�;�,�0.�-Ұ@�xH3��T0 k� �n��n&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�^�?A�|FaLd5�3�,�0.�-�B�xI3��T0 k� ��l��l&�1D"3Q	2�4#Q  ��_    � +�8��A_��AS�^�?A�|GaLd6�+�,�/.�.�D�xI3��T0 k� ��k��k&�1D"3Q	2�4#Q  ��_    � +�8�A_��AS�^�@A�xHaLd7�#�,�/.�.�F�xJ3��T0 k� ��i��i&�1D"3Q	2�4#Q  ��_    � +�8{�A_��AS�^�@A�tIaLd8��,�/.�/�G�xK3��T0 k� ��g��g&�1D"3Q	2�4#Q  ��_    � +�8w�A_��AS�^�AA�pIaL`9��,�..�/�I�xL3��T0 k� ��e��e&�1D"3Q	2�4#Q  ��_    � +�8s�A_��AS�^�AA�pJaL`:N�,�..�0�K�xM3��T0 k� ��c��c&�1D"3Q	2�4#Q  ��_    � +�8o�A_��AS�^�BA�lKaL`;M��,�-.�0�L�xM3��T0 k� ��a��a&�1D"3Q	2�4#Q  ��_    � +�8k�A_��AS�^�CA�hLaL`<M��,�-.�1�N�xN3��T0 k� ��_��_&�1D"3Q	2�4#Q  ��_    � +�8g�A_��AS�^�CA�dMaL\=M��,�-.�1�O�xO3��T0 k� �|]��]&�1D"3Q	2�4#Q  ��_    � +�8c�A_��AS�^�DA�dMaL\=M��,�,.�1�Q�xP3��T0 k� �|[��[&�1D"3Q	2�4#Q  ��_    � +�8_�A_�AS�^�DA�`NaL\>M��,�,.�2�S�xP3��T0 k� �xY�|Y&�1D"3Q	2�4#Q  ��_    � +�8[�A_{�AS�^�EA�\OaL\?M��,�+.�2�T�xQ3��T0 k� �tW�xW&�1D"3Q	2�4#Q  ��_    � +�8W�A_w�AS�^�EA�\PaLX@M��,�+.�3�V�xR3��T0 k� �pT�tT&�1D"3Q	2�4#Q  ��_    � +�8S�A_s�AS�^�FA�XPaLXA=��,�+.�3�W�xS3��T0 k� �pR�tR&�1D"3Q	2�4#Q  ��_    � +�8O�A_o�AS�^�FA�XQaLXB=��,�*.�4�X�xS3��T0 k� �lP�pP&�1D"3Q	2�4#Q  ��_    � +�8K�A_k�AS�^�FA�TRaLXB=��,�*.�4�Z�xT3��T0 k� �lN�pN&�1D"3Q	2�4#Q  ��_    � +�8K�A_g�AS�^�GA�PSaLXC=��,�*.�4�[�xU3��T0 k� �lL�pL&�1D"3Q	2�4#Q  ��_    � +�8G�A_c�AS�^�GA�PSaLTD=��,�).�5�]�xU3��T0 k� �hJ�lJ&�1D"3Q	2�4#Q  ��_    � +�8C�A__�AS�^�HA�LTaLTEM��,�).�5�^�xV3��T0 k� �hH�lH&�1D"3Q	2�4#Q  ��_    � +�8?�A_[�AS�^�HA�LUaLTEM��,�).�5�|_�xW3��T0 k� �hF�lF&�1D"3Q	2�4#Q  ��_    � +�8;�A_W�AS�^�IA�HUaLTFM��,�(.�6�xa�xW3��T0 k� �hD�lD&�1D"3Q	2�4#Q  ��_   � +�8;�A_S�AS�^�IA�DVaLTGM��,�(.�6�tb�xX3��T0 k� �hB�lB&�1D"3Q	2�4#Q  ��_    � +�87�A_O�AS�^�IA�DVaLPHM��,�(.�6lc�xY3��T0 k� �hA�lA&�1D"3Q	2�4#Q  ��_    � +�83�A_O�AS�^�JA�@WaLPHM�,�'.�7hd�xY3��T0 k� �h?�l?&�1D"3Q	2�4#Q  ��_    � +�8/�A_K�AS�^�JA�@XaLPIMw�,�'.�7df�xZ3��T0 k� �h=�l=&�1D"3Q	2�4#Q  ��_    � +�8/�A_G�AS�^�KA�<XaLPJMs�,�'.�7`g�xZ3��T0 k� �h;�l;&�1D"3Q	2�4#Q  ��_    � +�8+�A_C�AS�^�KA�<YaLPJ]k�,�&�8Xh�x[3��T0 k� �h9�l9&�1D"3Q	2�4#Q  ��_    � +�8'�A_?�AS�^�KA�8YaLPK]g�,�&�8Ti�x[3��T0 k� �h8�l8&�1D"3Q	2�4#Q  ��_    � +�8#�A_;�AS�^�LA�8ZaLLL]_�,�&�8Pj�x\3��T0 k� �h6�l6&�1D"3Q	2�4#Q  ��_    � +�8#�A_;�AS�^�LA�4[aLLL][�,�&�9Hl�x]"���T0 k� �h4�l4&�1D"3Q	2�4#Q  ��_    � +�8�A_7�AS�^�MA�4[aLLM]S�,|%�9Dm�x]"���T0 k� �h2�l2&�1D"3Q	2�4#Q  ��_    � +�8�A_3�AS�^�MA�0\aLLN]O�,|%�9<n�x^"���T0 k� �h0�l0&�1D"3Q	2�4#Q  ��_    � +�8�A_/�AS�^�MA�0\aLLN]G�,|%�|:8o�x^"���T0 k� �h.�l.&�1D"3Q	2�4#Q  ��_    � +�8�A_/�AS�^�NA�,]aLLO]C�,x$�x:0p�x_"���T0 k� �h-�l-&�1D"3Q	2�4#Q  ��_    � +�8�A_+�AS�^|NA�,]aLHO];�x$�t:,q�x_"���T0 k� �h+�l+&�1D"3Q	2�4#Q  ��_   � +�8�A_'�AS�^xNA�(^aLHP]7�x$�p;$r�x`"���T0 k� �h)�l)&�1D"3Q	2�4#Q  ��_    � +�8�A_#�AS�^xOA�(^aLHQ]/�x$�l;s�xa"���T0 k� �h'�l'&�1D"3Q	2�4#Q  ��_    � +�8�A_#�AS�^tOA�$_aLHQm+�t#�h;t�xa"���T0 k� �h&�l&&�1D"3Q	2�4#Q  ��_    � +�8�A_�AS�^tOA�$_a<HRm'�t#�d;u�xb"���T0 k� �h$�l$&�1D"3Q	2�4#Q  ��_    � +�8�A_�AS�^pPA�$`a<HRm�t#�`<v�xc"���T0 k� �h"�l"&�1D"3Q	2�4#Q  ��_    � +�8�A_�AS�^pPA� `a<HSm�\t#�\<w�xd3��T0 k� �h �l &�1D"3Q	2�4#Q  ��_    � +�8�A_�AS�^lPA� aa<DSm�\p"�T<�x�xe3��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8�A_�AS�^hQA�aa<DTm�\p"�P<�y�te3��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A_�AS�^hQA�ba<DTm \p"�L=�z�tf3��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A_�AS�^dQA�ba<DUm\p"�D=��{�tg3��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A_�AS�^dQA�ca<DUm \p"�@=��|�ph3��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A_�AS�^`RA�ca<DVl�\l!�<=��}�ph3��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A_�AS�^`RA�ca<DVl�\l!�4>��}�li3��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A_�AS�^\RA�dZ�DV|�	\l!�,>��~�lj3��T0 k� �h�l&�1D"3Q	2�4#Q  ��_   � +�8 ��A_�AS�^\SA�dZ�@V|�\l!�(>���hk3��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A_�AS�^XSA�eZ�@V|�\h!� >ἀ�dk3��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^XSA�eZ�@V|�\h �?ᴀ�dl"s��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^TSA�fZ�@V|�\h �?��`m"s��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^TTA�fZ�@V|�\h �?��\m"s��T0 k� �h
�l
&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^TTA�fZ�@V|�h �?��Xn"s��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^PTA�gZ�@V|�d �?��Xo"s��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^PTA�gZ�@V��d�@�~�To"s��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^LUA�gZ�@V��d�@�~�Pp"s��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^LUA�hZ�<V��d�@�~�Lq"s��T0 k� �h�l&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^HUA�hZ�<V��d�@|~�Hq"s��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^HUA�hZ�<V��d�@t}�Dr"s��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^HUA�iZ�<Vܼ!`�Ap}�@s"s��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^DVA�iZ�<Vܸ#`�Ah}�8s3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^DVA� jZ�<Vܸ%`�Ad}�4t3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^DVA� jZ�<Vܴ&`�A\}�0t3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^@VA� jZ�<Vܰ(`]�AX|�,u3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^@WA��jZ�<Vܬ)`]�BP|(u3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^<WA��kZ�<Vܨ+\]�B!L| v3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^<WA��kZ�8Vܤ,,\]�B!D|w3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^<WA��kZ�8Vܤ.,\]�B!@|w3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^8WA��lZ�8V�0,\]�B!8{x3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^8XA��lZ�8V�1,\]xB!4{x3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^8XA��lZ�8V�2,\]pC!0{y3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^4XA��mZ�8V�4,\]hC!({ y3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^4XA��mZ�8V�5,XM`C!${�z3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^4XA��mZ�8V�7,XMXC! {�z3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^0XA��mZ�8V�8,XMPC!z�{3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^0YA��nZ�8V�9,XMHD!z�{3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^0YA��nZ�8V�;,XM@D!z�|3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^,YA��nZ�8V�<,XM4D!z�|3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^,YA��nZ�8V�=,XM,E!z�|3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^,YA��oZ�8V�?,XM$E! z�}3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^,ZA��oZ�4V�|@,TMF �y�}3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^(ZA��oZ�4V�xA,TMF �y�~3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^(ZA��oZ�4V�xB,TMG �y�~3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^(ZA��pZ�4V�tC,TMG �y�3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^(ZA��pZ�4V�tE,TL�H �y�3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^$ZA��pZ�4V�pF,T<�H �y�3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^$ZA��pZ�4V�lG,T<�I �y☀3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^$[A��qZ�4V�lH,T<�I �x␀3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^ [A��qZ�4V�hI,T<�J �x�3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^ [A��qZ�4V�hJ,P<�K �x�3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^ [A��qZ�4V�dK,P<�L �x�x3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^ [A��rZ�4V�dK,P<�M �x�p3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^ [A��rZ�0V�dL,P<�N �x�h~3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^[A��rZ�0V�dL,P<�O �x�\~3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^\A��rZ�0V�dL,P<�P �w�T~3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^\A��rZ�,V�dL,P<�Q �w�L~3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^\A��sZ�,V�dM,P<�Q �w�D}3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^\A��sZ�,V�dM,PܤR �w�<}3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^\A��sZ�(V�dM,PܠS �w�4}3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^\A��sZ�(V�`M,LܜU �w�,}3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^\A��sZ�$V�`M,LܘV �w�$|3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^\A��sZ�$V�\N,LܔW �w�|3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^]A��tZ� V�\N,LܐX �w�|3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^]A��tZ� V�\N,L܌Z �v�|3��T0 k� �k��o�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^]A��tZ�V�XN,L܈[ �v� |3��T0 k� �o��s�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^]A��tZ�V�XN,L܄\ �v��{3��T0 k� �o��s�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^]A��tZ�V�TN,L܄]�v��{3��T0 k� �o��s�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^]A��uZ�V�TNL܀^�v��{3��T0 k� �o��s�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^]A��uZ�V�PNL�|_�v��{3��T0 k� �s��w�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^]A��uZ�V�POL�xa�v�{3��T0 k� �s��w�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^^A��uZ�V�POL�tb�v�{3��T0 k� �s��w�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^^A��uZ�V�LOH�ld�v�z3��T0 k� �w��{�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^^A��uZ�V�LO\H�le��u�z3��T0 k� �w��{�&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^^A��vZ�V�HO\H�hf��u�z3��T0 k� �{���&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^^A��vZ�VLHO\H�dg��u�z3��T0 k� �{���&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^^A��vZ�VLDO\H�`h�|u�z3��T0 k� �����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^^A��vZ�VLDP\H�`i�xu�y3��T0 k� �����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^^A��vZ�VLDP\H�\j�tu�y3��T0 k� �����&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^^A��vZ�VLDP\H�Xk�pu�y3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^_A��vZ�VLDP\H�Tl�lu�y3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS�^_A��wZ� VLDP\H�Tm�huxy3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^_A��wZ� VLDQ\H�Pm�dupy3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^_A��wZ� V<@RH�Ln�`uhx3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^_A��wZ��V<@RH�Lo�Xu!`x3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^_A��wZ��V<@SH�Hp�Tt!\x3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^_A��wZ��V<<TH�Dq�Pt!Tx3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^_A��wZ��V<<UH�Dr�Lt!Lx3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^_A��xZ��V<<UD�@s�Dt!Hx3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^_A��xZ��V,<VD�<s�@t!@x3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^_A��xZ��V,<WD�<t�8t!<x3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^_A��xZ��V,<XD�8u�4t!4w3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^`A��xZ��V,<YD�8v�,t!0w3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^`A��xZ��V,<ZD�4w�(t!(w3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^ `A��xZ��V,<[D�0w� t!$w3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^ `A��xZ��V,<\D�0x�t!w3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^ `A��xZ��V<]D�,y t!w3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^ `A��yZ��V<^,D�,z t!w3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^ `A��yZ��V<_,D�(z t!w3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^ `A��yZ��V@`,D�({  t!v3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^ `A��yZ��V@a,D�$|�t! v3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^ `A��yZ��V@b,D�$|�s �v3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|^ `A��yZ��VDc,D� }�s �v3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�`A��yZ��V�Dd,D� ~�s �v3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�`A��yZ��V�He,D�}�s �v3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�`A��yZ��V�Lf,D�}�s �v3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8 ��A^��AS|]�aA��yZ��V�Lg,D�}�s �v3��T0 k� ������&�1D"3Q	2�4#Q  ��_    � +�8                                                                                                                                                                            � � �  �  �  d A�  �K����   �      6 \��� ]� 4 3 8 ����    �	   �  T�    ��  ]     <��   	             � �          �       ���   0	&
         ��[?         �����    ��Z�����     �e   	                 <�        �     ���   (	           �U       ���     �U ��?      ��              	   ��        �     ���   0
           bK�           �{W�     b�F�{�%    �&��   	             A�$          0     ���   H
$
          }�n          /�q�     }՛�qb     ���                  ��$           �     ���   0
3            V�. ��     C���     V�.��4>      ��                      ���w                ���    P		 5              [��  � �     W�G�     \=�H�    �W��             g Z�8         �P�     ��`  (
	           �    
	   k�ޤ      ���]    ����             2  Z�8         ��     ��H   8	 

          b��  M M    �'g     c�$�%�    ��             -	 Z�8         � �  �	  ��@  		�           s�%  > >       ��~�x     s'���e�    ��S             
 Z�8         	 6 �     ��@  0
3
          r��  A ]
	     ���MT     r����L�    ���                , Z�8         
  p�    ��@  H


         ���� ��
	      � ��Q    ���� ��Q                              ���]                 ��@    		 5 	                 ��      �                                                                           �                               ��        ���          ��                                                                 �                         �~N�  ��        ��
��  W��~i��
Xi  W��n�                   x                j  �   �   �                         �~    ��        ��      �~  �           "                                                 �                           �� ��{�q���G��'�~�� ����
�  
         	      
  B   ��� ��B       3� �o� 4� p� B� q  #� `j� $d k� &� s@���J ����X ���� ����  ����. ����< ����J ����X � 
�< V� 
� W  
�| W  @� 0u� A v@ A$ v` D� s` �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� � }����� ����� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����8�� +�� �  ������  
�fD
��L���"����D"� �  " `   J jF��    "�j "���
��
���     �j��  
  �
� �  �  
� ����  ��     � |  �    V   ��     ���           ��     ��          � ��   �    ��        LL     �    ��        MM     �    ��        a�         �    ��  �_	 5       �� � �  ���        � � �  ���        �        ��        �        ��        �    �     �x>����        ��                         T�) ,  ����                                      �                 ����            �� ~���&��   +�8��               18 Denis Savard                                                                                     6  5      � KC0&KD(� �� �ck �$ cs � �c. � c�& �	cW$ � 
cc, �K/G � K7W �C/ � C#7 �c�@ � c�P tJ� � � J� �E"�#E "�55"�5*�*$"� �$ "� �� �
� � �*;u �)�u*=u0*}8 *M]X  *LMP  *SeP  *SeX #*LMP  *SeH %*QMP &*PeX  *IM(*}8 )*E]0**}P +*DeX ,*HmX  *LMX  *LMX /*HmX  *LM 1"' |  "+ | � 3"K �-  "! | � 5"F � � 6"B � � 7"Q �  8" �@  "F � � :"B � ;"Q � <" �S  "F � >"K �0 !� |                                                                                                                                                                                                                         �� P         �     @ 
        �     Y P E k  ��                    ������������������������������������� ���������	�
���������                                                                                          ��    �^�� ��������������������������������������������������������   �4, E� B 9�� �  ۂ �@ @$��@����@����@���A(��&�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     '    ��  �D�J      Te  	                           ������������������������������������������������������                                                                                                                                       ���� ��                                             �������������������������� ������� ����� ����������������� ��������������� � ������������� �����������  ���� ��� ���������������� � ����� ���������������������� � ������ ��� ������������������ ��������� �� ������������ � ��                                   V    '    �� �\�J     0�                             ������������������������������������������������������                                                                                                                                         ��<�  � J�                                           ����������������������������� �� ����� � ��������� ��������������� ����������� ������������ ��������������� ���������������� �� ������������������������� ���������������������  ����������� �������������� ������������� ��������                                                                                                                                                                                                                                                                                                                         �              


             �  }�         ����          J7����  W  K����������������������������������������������������������������������������  �  [�  c�               Y                                                      ""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" : D 7                                  � ��� �o�                                                                                                                                                                                                                                                                                      )n)n1n  YE        k      k                              k      k                                                                                                                                                                                                                                                                                                                                                                                                         > �  >�  J�  <�  
�  Fa�  �̞�T�̞�x��0�+��� |����|��H�,�̞������                      �� r        $   �   & QW  �   �                  �                                                                                                                                                                                                                                                                                                                                        K K    �                       !��                                                                                                                                                                                                                            Z   �� �~ ���      �� \     �������������������������� ������� ����� ����������������� ��������������� � ������������� �����������  ���� ��� ���������������� � ����� ���������������������� � ������ ��� ������������������ ��������� �� ������������ � ������������������������������� �� ����� � ��������� ��������������� ����������� ������������ ��������������� ���������������� �� ������������������������� ���������������������  ����������� �������������� ������������� ��������             $����������������˪�������������������������������������f��ff��ff�������̺�ff�fffffffffffffffffff����ƹ��ffʻfff�fffjffffffffffff��������������������ʺ��l���f˪������������������������������������������������������������������fff�fff�fff�ffk�ffi�ff��ff��ff�ffffffff�fff�x�����w��xx�������wfffffff�ffff�fffww��ww�x����wx��fk��ff��ff��ffʹffj��fʪ�f�ˊ�k������������ʚ��������������������������������������������˫��ʫ��ff��fl��fl��ff̫fff�ffʬ�f���f�����������wu���w��l������f����W��������xww��Wy�l����x������k���W�fi���j���j���f����˘�����y�y�y����������������������������������������������������ʻ����ʫɚ�����l���ƨ�lƘ�j���k���̜i���j���kxx���wx������wx������������ƈx����������������wW����w�������������������������z����������˫��̺������������������������������������������������������������ʺ������k������������������������������������������x�j���˙�x�˘��̩�x������x���xx�x������x������wx���˫��ʫ����������˪�����ʻ��������������������������������������ʻ�ʻ�����ʪ̫����˺��������������������˪�����f���k��f��fǶW�g���k���̻���f������������������x�������˩f̺�����uw�����w��x�wXx��˪�����������l����l���i��ƹx�f�������������������ʫUW��UUU�UUUX      7      4   � �~                       4     �  �����J����'      ��     ��      �            �   �   �      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��   ( ����  �� �� �    � �N ^$   ��B   (  ��   )  �1   �   ��Ҍ����������J����  ��    # ��     F�  ��    ���   ����� >�������J J�������   �����   i ��   ��     ��   �� �� �z  ���� �$ ^$   �   ��   	  ��  �� �� o� �� �� �z o� 3� �$ 0 �  ��R  �      �  ��   �������2����  g���        f ^�         ��� +            ��Z���2�������J����  ��      y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N���wwwtwwwtwwwtww~Dww�wwH4wwH4wwH4�wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwwwwww�wwwGwwwGwwwGwwwNwwwDwwwDwwwwwwwwwwwwwwwNwww��ww8Gww8Gww8GwwwtwwwtwwwtwwwtwwwtwwwtGwwwGwwwGww~H4w~D�ww��wwwdwwwvwwwtwwwdwwwv8Nww�Nww��ww�wwwwwwwgwwwwwwwwwwwwwwtwwwdwwwvwfwtvwfdc337eUUTEUUTGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���Dwww��wwD�ww�GwwDGww�GwwDGww�Gwwgwwwwwwwwwwwgwwwwwww3333UUUUUUUU         D �  H4wwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNww�DwwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c      ������������  9�  	�  �  �  �   �   9   9                  �����������ߚ�����������	������ 9�� �� ��  9�  �   9       ����������������������������8���      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0       ��� ��  �   8                ����������������8��� 8��  ���������������������������������8���                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���w           N  �� 8@ DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    8888����������������������������8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w  H4 H4H4 D�  ��   d    DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0       ����������������������������������������������������������������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8�����������������������8��� 8��  �    ����������������������������3:������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                      ��������������������������������                                8@  8@ 8N �N ��     `      d    d       d  DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   �   ��� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5    �  �  ���������  	�  	�  	��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53  �������������������w~욪��"""��""��""�r""rb""gb""w"""""""̹���˜��̽���ͻ�ۧ�̺�w̚�~�����"""��""��""�r""rb""gb""wU""�CR"���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#2"��""��""�r""rh�"gk�"wU�"�CR"�#2"��""��""�r""rh�"gk�"wU�"�CR"������������ۻ������_��SU  U5  �����۽�ۻ�۽�۽��������        ��������������۽��������        ~���~���~���~���~���~���~���~���̋��̛��˘�̽����8���U8���S3۹��"̚�"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"UuW�UvW�UgW�UTW�UWg�www�������������wwwCGww34ww33wws3wwt33333333��""��""��""+�""""""""""""""""""                             ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                      wwwwwwwwwwwwwwwwwwww3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UUUGwwwWwwwTwwwTwwwWGwwWGwwWGwwWt3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               �DDE�fDMffDMffDMffDD3333UUUUUUUUwwWtwwWtwwWwwwWwwwWw3333ff6fff6fwwwwgwwwGwwwGwwwFwwwtwwwtwwwvgwwffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0tDDtTDDtDDDDDDIDDD��3333UUUUUUUUffVfffVfffVfffVfffVfwwgwDDgw��gwuuwwsvwwsgwwsT��sWl�sVw�sUG�sUg�uUUU|UUU|UUU|UUU|�UU|�gw|���|���#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�swwwswwwswwwEwwwFwwwE333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP U3U�ۻۻ�ۻݻ�۽ݽ������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  B  @  @  @                                                    !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3                                                    @ B   @  @   B   @ `   P                                                ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfffFfDvFfDDDv����    `       a   fff d                                                                4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffdfffdfffffff                                                                ����������������������������DDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDffUUddUUffUTddUDffwDf�D�f�D�ffD�DDDDgwwtGwwtDwwtDwwtDwwt�Dwt�DGtfUDIUUDDU�TMU�DMeUDDefDDffDDffDDTDDtDDDtDDDDDDDDDDDDDDDDDDDDDDDtffDDddDDdfDDffDDfFDJffDIfDDJdDDGDDGtDwwtDGwtDGwt�GwtzGwt�Dwt�DGt"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD���������������������������������������������������������������������������������������                      �  9� ��  P                             3333333333333333333333333333333333333DD34DD34��33��33��33��37ww37wrsww!wwwqwwwqwwwqwwwqwwwwDwwtGs3www�www�wwwwws7wws7wws7wws7wws7wws7wws7wws7www7www7www3ww3333333333DD34DD34DC33D�33��33>�37ww37wwswwwwwwwwwwwwwwwwwwwwwwwDwwtGww37ww�ww~�7www7wws7wws7wws7wws7wws7wws7wws7wws3www37ww33ww3333UUUUwwwwwwwwwwwwwwwwwwwwwwwwwwww�"""+�""���"��̲r'&"wvv"��r"��""�����˚��̸���̽��̌̽��̽�˻��˻""")�""���"����}�&"wvv"��r"��""���̋��̛��˘�̽����8��۪8���3۹"̑"ܹ�"���"���"��""˞""˸""�5S=��S��Y3���S���"���"���+���-���"���"ع����������=��"۹�"���"��""��""��""+�""""""""""""""""""wwwCGww34ww33wws3wwt33333333                                                  U  T   T   T     T UDUDDUDDDDDDDDDDDDDDDP   E�  DU� DDU�DDDUDDDDDDDDDDDD                UP  E�  E   E                                           ���U�UTD�DDDDDDTDD TDD   �   U_ DEU�DDDUDDDDD��DZT�DDDDDDDDDDDDTDDDDDDDDUTU�����DDDDDDDDDDDEDDDEDDDDTUTU�Ԫ���Z_   P   � �U�UTDUDDDDUTD�DT��D        U_��DEU_DDD_DDDPDDE�DDE  �DD DD DD �DD �UD  �U       DZTDEDDDDE�DDE�DDE�TDDT�DE�TE���DDTU�ZD���������DDTDD��ZT�T���ZTDDE��D��T�T��DUTTT��Z��TQTDDUTD�DDDTDDD�DDDDDDE�DD_TDE�DD_ DDP DDP DD_ DU_ U�  �                                       TE�DDD�UUU                    ���DDDUUUTD  D  D  D  D  U��D�TDDDDEUUDP  DP  DP  DP  UP  TDE�DDDPUUU_                                                    wwwwtDDDt""$t"""t"w"t"w"t"w"t""$wwwwtDGtD"GtD"GtD"GtD"GtD"GtD"GtwwwwDDDD"D"""D"""DD""Gt""Gt""Gt"wwwwDDDD"B"""B""DDD"GwD"GwB$GtB$wwwwDwww$www$wwt$wwtGwwtGwwwwwwwwwwwtDDDD�DLL�D���D�D�D�t�D�t�D�wwwwDDww��Gw��Gww�Gww�Gww�Gww�Gwt"""t"w"t"w"t"w"t"""t""$tDDDwwwwD"GtD"GtD"GtD"DDD""$D""$DDDDwwww"Gt""Gt""Gt""Gt""Gt""Gt"DGtDwwwwGt"DGD"DGB$GGB$DGB""GB""GDDDwwwwwwwwwwwwwwwwDwww$www$wwwDwwwwwwwt�D�t�D�t�D�t�D�t�D�t�DMtDDDwwwww�Gww�Gww�Gww�Gw��Gw��GwDDwwwwww���������������333wwwwUZ��UZ��UZ��UZ��UZ��3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ�#UZ�#UZ�#UZ�#UZ�#3333wwwwUZ"#UZ"#UZ"#UZ"#UZ"#3333wwwwUR"#UR"#UR"#UR"#UR"#3333wwwwU""#U""#U""#U""#U""#3333wwwwR""#R""#R""#R""#R""#3333wwww"""#"""#"""#"""#"""#3333wwww���������������333wwww��"��"��"��"��"333wwww��"��"��"��"��"333wwww�""�""�""�""�""333wwww�""�""�""�""�""333wwww"""""""""""""""333wwww"""""""""""""""333wwww                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "!  "! " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��               "!  " ! " "" """ "!   " ""                                                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """ "!    " ""            """                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                                     �   �   w   b   g     
�  �� �� �� �̻ ������ɨ�-�ݼ-ݍ�"Չ� X���DDX�TCZES3�T3�@ ��"��"�� ""� �"/��/��        �   ��  ��  ��  {�  wp  ��� ���������̻��̽��̽���ؚ��ڨ��؛˻��˸� ��  �C  D0  3   0   0   �   �   �    �  /   ���                     2�  2   1   �                  �    � .� .  �� 	  
  �  ",  ""  �"   "                      �"  �"  �      �         "   "   �                       ".  ".  ���                    � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                         	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��  T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ��"� �"� ����            �   �   �   D   E�  U�  UO                         "  "  "    �   �   .   .�   �       �                                                                                                                                      ̰ �ˉ",ɩ""��""��"/���    ���̻��̻�����w��rg���&z��wڻ��H�̹������̻�̿�˿ ��� ����      "   "   "   "  �" �� �ȯ D�� TD� UC�U3�TD4ETE�4EU���E                    �  �  "� � �� �ɫDKˏET��UX��U�� T�  H�      "   "   "   "�  /�  �   �   ̻����ߪ����� �                         �  � ��� ��  �   �ˀ ��� ����������+� ""��"�""��"/� ����                                     �"  �"  �                  �  ".��".� ��             "   "   "�  �                            �   ���                            �   "    �                                                                                             	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��   �� �̽���ݪ۽w�}�&��vv���p���                             ��                     �   �                      �".��".  ���    �  �   �   �   �  �  �  �  �  ���                                                                                                                                                                                             �� ��� ��� ww� &'� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                               " "/ �/� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  &'  vv  w                �                        ��"� �"� ����                            ".  ".  ���                 ��                               �   ���                            �   "                                                                                                                     �� �����ݼڜ��ک��ک��z�	��� 
�� 
�� 	�� ̘ ɪ  ��  �  �� �� ������������ ���  � � � �� "� "��"�/ ��                      �   ��  ��  �̰ ��� ��˰�̻��̻���������ˉ�U��EP�ET �I� ٕ  �D� �L� ��� ��" ����/�"�"�""�����                         ��� �"" ��" �""��"��"  �!� "    �  .        .   �          �     �       �              !   "  �  �!  �"  �"  �                   �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  "   "                                                                      �  �� 
�� ɨ�˻�+�""� "�  .    �  �  �   �  E  E  U  D  D  �   �   �   �   "  "  �" �"   �                    �gz���������˻����̽��̽��̰��˰�������@DDDDTDDTUDET�@EU^@ETD�TD�DL D� �  ��  �   ,   "   "/ �"��������           �    �   �   ̰  ��  ݚ� ��  �"� "   ""  ""       @   H   H   D   D   L   �   �   �   ��  .�"." "."   /�  �  �              � ��         �� �� �� g} &' vw     �     "   "                   ��   �  ��  �  �  �         � ".��".��/����  �                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� &'��vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   "   "�  "�  ��  ��    ""  ""       @   H   H   D   D   L   �   �   �   ��  .�"." "."   /�  �  �              � ��         �� �� �� g} &' vw                     ".  ".  ���     ��   �  ��  �  �  �         � ".��".��/����  �                                                                                                                                         ˰ ̻ ̻ �� {�  �� 
�� ��� ��� ������
���	��ܻ̍ݻ���"� 8"  8  �  D�  H�  X�  ��  �   �          "  "     �                        ��  ��� �̺�̻����ۻ�˽��̽��̝ ̙� �30 �EP �U@ �T0 EC0 T3  C:  K�  �"  �"/ ����˽� �"� "" �""� � �� ��      �   �  .�  ."  �            �   �"  ""  !� �� ��  �               �   " ��.�  ��                                                    �               �     "   "               ���                                                �   ���                            �   "                                                                                                    � 
��	�˽���w��rb��gg�Ͷw��ۻ+=�"D3
.�4
DE��E �� 	��  ��  ʠ  ��  "   "  " �"�� ���    �   ٜ  ک� ��� ��� ��� �ۜ��٩�3;� C"� �"- ��  "��  �   "  �"/�� �� � ��     �            .  .     �   �            ��  ��                                �  "� "     �   �            �   "   "  "             �  ��  ��  ww  &'  vv  w                �                        ��"� �"� ����            ����  �  �  �  �  ��  �                      � �� �                  �  � �                       � �� �                 ��� "   "   "   "        ��   .  .  "  "  �   �             �  �                                  �� �� ���
��ۘ�g}˷&'̶vw��g{�� �˰ "   "�  .       �  �  "   "                           ��  ��� ʜ� ʩܰ��͹��͹������̄���Dݻ�E���E	��U̚3E��34̰�   �      �   �          �   �   X�  X�  U�  UH  T�  K�  ��� ڬ� ۻ� +�" """ """ �"" ��"/����� ��   .   .   ��                        �          �   � � /  �"" �"  �    "   "   "  �� ��                   �".��".���                            �   ��  "   "   �   "  "  "   �                                                                                                                                                                                     �  �  �� 	� 
� ɩ �� 蘰 ��� ��������  ��  �   �      �  �   �   �         ��� ݼۼ����))������؜������ ��� 3���34ۍ�5��������ݘ ��������������������� �������� ����    �   ��  ��� ݻ� �ۘ ��� ɩ� ��� ]�S ڌ0 ��  ��� ��� ��� ������������������������������� ����"  �". �.  �                                        �� ��                  �          �         �   �  �  �   �               �   �               � . "/��/ ��                                                                                                                                                                                             2  %  2P  % P0 # R00 S�� :�� Y� :�0 Y�*�5Y�U """####RP00000000000000��������00005555UUUU""""####0002#0002#0002#0000��������00005555UUUU 2:� #	� :�#	�P:�	�P:�%	� Z� %	� 2Z� 9� *�                                                                                                                 �� 
22  0 
3  0 
2 �0 
23 �" 
02 � 
00 � 
00 � 
00 � *003�"000#0000# 000# 000" 00 "  0  ""    ����2222000000000000000022220000000000000000000000000000000000000000""""    ����2223000200020002000222220002#0002#0002#0002#0002#0002#0002#0002#0002#0002""""                                                                                                                                                                                    D@ DD D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I��""""�������AD�I�""""����������������I���I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�I��I��I��I���I�����3333DDDD���D�I�DD�����3333DDDDAIA�II��I�D����3333DDDDI����D��DI����3333DDDDA�A�A����D������3333DDDDI��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDDI���I���I���������������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""����������A��I��I""""����������IAIA""""�������DI���""""������DI�I�""""�����A�DA�I��I�""""�������A��AA""""�������DD�I""""������D��""""��������I���I���I���I���"""$���4���4���4���4���4���4������������������333DDD��M��M��M��M���M����3333DDDDMAMAMMMM�M�M����3333DDDD���D�M�DD�����3333DDDDM�M�M�M��M�D����3333DDDD�M��M��M��M���M�����3333DDDDD�����MD��M����3333DDDDDM����DD�����3333DDDDADAM�M�M�D�����3333DDDDM���M�������DD������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                        """�"""�                                             � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��                              ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   �"" �""       �  �     �  � "�� "�                                " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        �             ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      �  �                      �""��""��           �   �                         �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                                  �   �   �   ��" ��"                        ".� ".�                                   �                 � ���и���݊��    �   �   �   ��""�""                        "�  "�              DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                                  �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      �""�""" "          ����            �   �       �   �                   �   �  �  �wqqwqwqDwqDGwwwwww3333DDDDADAwAwADwtGwwww3333DDDD � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(�GwDGwqwDDwtwwww3333DDDD �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(�""""����������A��I��I = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=""""�����A�DA�I��I�    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( """"��������I���I���I���I��� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(XxMAMAMMMM�M�M����3333DDDD w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xwwD�����MD��M����3333DDDD  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���4���4���4���4���4���43334DDDD �  + � � � � � � � � � � ��	� � � ��� � � � � � � � � � � ��	� � � ��� �� ����(+((�""""wwwwqqqqwGwGGG ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`""""wwwwwwqqDAwG M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M������������������333DDD � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(�M��M��D��M����������3333DDDD � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(�DD��D�M��D����3333DDDD 5 6  X � �F � � � � � ����� � ����������� � ����� � � � � ��	F ��(X((6(5""""������DH�H� x �  l � �G � � � � � � � � � � ������������� � � � � � � � � � ��	G ��l((�x""""�������H�H��D w w x y ������H���������������������������������H�����yxww""""��������H��H��H��H�  � + w�������I�J�K�L�M�N�O � � � � � � � � � � � � � � � � � � � ��O�N�M�L�K�J�I������w(+�(DD������L��DL����3333DDDD , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A e ��A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,L�A�AAD��DL�����3333DDDD +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�] � ځ]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+���4���4���4L��4L��4���43334DDDD 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U �h�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5""""���������M�MMM =  U ,     !d�P���e�f�g�!�!�!�k�!�!�!�l�!�!�!�!�k�!�!�!�l�!�!�!�g�f�e���P)d((( ((,(U((=""""�������A��AA     =  U , N ,�-�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�p�-(,(N(,(U((=((( ��������������333DDD � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � �I��I����������������3333DDDD � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � ���A���I��I���I�����3333DDDD m � �!�A�A� � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`""""������������������������  � �!�AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M""""������D�D��� 
 � �!�AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(�""""������������������������ - � �!�!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(�wqwwqwwwwwqwwwDwwww3333DDDD 69�:���  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5qqwwwDDwtGwwww3333DDDD x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�xwww4www4www4www4www4www43334DDDD w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww""""wwwwwwqwwwqwqwq + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+""""wwwwwwwDwGwA � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(��A�L�L�L��L���333DDDLDD�L��L��L���L����3333DDDDA�A�A�A��LD�����3333DDDD�����ADDLD����3333DDDDADA�A�A��LD����3333DDDD�A�ALD��DL������3333DDDDDLL��LDD�D����3333DDDD�A�LDL�L�D�L�����3333DDDDLD�L�L�L��L�����3333DDDDA�A�A�A�LD�D����3333DDDDL4DL4�L4�L4��L4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD""""(���(���(���(���(���(���""""������������������������""""��������������������""""�����ADAHA�A""""��������H�A�A�A""""����DDD�AHA""""�������ADH""""������HDAD�H��""""����������D�����������""""������������������������"""$���4���4���4���4���4���4(���(���(���(���(���(���#333DDDD������������������������3333DDDD���������������������3333DDDD�A�AHH�DH��H�3333DDDD�A�AHH�DDH�����3333DDDDDHH��HDD�D����3333DDDDAD��D�DH������3333DDDDD������H�DH�D����3333DDDD��������������D�������3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwwwwwwwwwwwwwwwwwww""""wwwwwqqDDqwwww""""wwwwwwqwDqq""""wwwwwwDGqGq""""wwwwwwwwwwwwwwwwwww""""wwwwwqGADAGqAwq""""wwwwwqwDDwq""""wwwwwqGADDqwqG""""wwwwwwwwwwwwwwwwwwwwwwww"""$www4www4www4www4www4www4������������������333DDD������������������������3333DDDD�������D�DDH����3333DDDDADAH�H��H�D����3333DDDDH�H�H�H��H�D����3333DDDD����������D��DH����3333DDDDA��A�H����DD����3333DDDD�A��DH��DD����3333DDDD�DHA��HH���DD����3333DDDD������������������������3333DDDD���4���4���4���4���4���43334DDDD""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUUUUUUUUUUUUUUUUUUU""""UUUUQQADDEUUQU""""UUUUUUADUQUUQUU""""UUUUUUQUUQUUQUUQUUQ""""UUUUUUQUUUQDUQEUQU""""UUUUUUUEEQEQE""""UUUUQUQEQEQEQE""""UUUUQUEDDEUUQU""""UUUUUUUUUUUUUUUUUUUUUUUU"""$UUU4UUU4UUU4UUU4UUU4UUU4(���(���(���(���(���(���#333DDDD������������������������3333DDDD�A���HHH�DD�����3333DDDD�����������D������3333DDDD���������H��H��D����3333DDDD�������H�DH�D����3333DDDD�HD�H�D�������3333DDDD�H�HHHDD�H����3333DDDD�A���HHH�DD�����3333DDDD KC0&KD(� �� �ck �$ cs � �c/ � c�' �	cW% � 
cc- �K/G � K7W �C/ � C#7 �c�@ � c�P tJ� � � J� �E"�#E "�55"�5*�*$"� �$ "� �� �
� � �*;u �)�u*=u0*}8 *M]X  *LMP  *SeP  *SeX #*LMP  *SeH %*QMP &*PeX  *IM(*}8 )*E]0**}P +*DeX ,*HmX  *LMX  *LMX /*HmX  *LM 1"' |  "+ | � 3"K �-  "! | � 5"F � � 6"B � � 7"Q �  8" �@  "F � � :"B � ;"Q � <" �S  "F � >"K �0 !� |3333DDDDAqAqAqAqGDwDwwww3333DDDDqAqGqGqGwDtGwwww3333DDDDGDwDwwGwwGwwtGwwww3333DDDDAwqAwqqwqqwqwDwwwwww3333DDDDwqwAAADDDwwwww3333DDDDGDGwGwGDwtGwwww3333DDDDDwqGwqwwqwwwDwwwwww3333DDDDwww4www4www4www4www4www43334DDDD"""������������������""""������������������������""""�����I�DA�I��I�""""�������DI���""""������DIAD""""�������AD�I�""""��������AA�A�""""�������ADI��I����������������������������������"""$���4���4���4���4���4���4������������������333DDD�����������������������������������D�I�DD�����3333DDDDAIA�II��I�D����3333DDDD��������������������������������I��I��I��I��I�D�����3333DDDDI����D��DI����3333DDDD��������������������������������""""%UUU%UUU%UUU%UUU%UUU%UUU""""UUUUUUEEQQQQQ��������������������������������""""UUUUUUQEDADUQEUQ""""UUUUQUUDEQUQ��������������������������������""""UUUUUQQADAQQ""""UUUUUUUAUQEE��������������������������������qwDwGwDwwtGwwwww3333DDDDADAGqGqtGwDwwww3333DDDD��������������������������������wqwDqGwDDwwwww3333DDDDGqqqwwtDDwwww3333DDDD��������������������������������DwwqwwGDwtGwwww3333DDDDwww4www4www4www4www4www43334DDDD��������������������������������""""��������AAAHA""""�������DDA��H���������������������������������""""���������DAAAq""""�����ADHA��H���������������������������������"""$���4���4��4��4H�4H�4�����������������333DDD��������������������������������M�M��AADMDDM����3333DDDDDAMAMAMA�M�M����3333DDDD��������������������������������M�M�M�M�DM�D����3333DDDD�M����������D����3333DDDD������������������������������������������������������������""""-���-���-���-���-���-���""""������������������������ �
�
�
�
�
�
�����������������������""""�������A��A�A""""�������A��A�A��� �
�
�
�
�
�
�=�[�H�Y�Z��V�M��[�O�L��2�H�T�L������""""������MDDMA��M""""��������������������������� �
�
�
�
�
�
�����������������������������������������������3333DDDD�DD�H�H����3333DDDD��� �
�
�
�
�
�
������������������������A�A�A�A��HD����3333DDDDAHHD�H��H���H������3333DDDD��� ��%��:�L�S�S�L��0�R�S�\�U�K���������8�>�7���������������������������3333DDDD���4���4���4���4���4���43334DDDD��� ����>�L�L�T�\��=�L�S�H�U�U�L��������>��<���""""������A�D��I��""""�������D����� ��$��/�L�U�P�Z��=�H�]�H�Y�K���������>��<���""""��������A��A�A""""������IDDAA��A��������������������������������"""$���4���4���4���4���4���4������������������������3333DDDD�����������������������������������������������������AA�DDD����3333DDDD�DALA�A��D������3333DDDD� ��	���&������������������ �8�>�7���"���A�ALL�DDL�����3333DDDDDL����������DD������3333DDDD� �ơǡȡɡʡˡ̤��������������� ��������""""'www'wq'w'qA'qG'q""""wwwwwqwqwqwAwAw� �͡ΡϡСѡҡӤ��������������� �>��<���!��""""wwwwqAGADwqwwqw""""wwwwwwqwDqq��������������������������������""""wwwwwwwwwGwwGwwqwwq""""wwwwwwqqqqqq"""$www4www4www4www4www4www4,�,�D,�����������DDA�A�AA�LDD����3333DDDD��������ALLDDL����3333DDDD��A�������DD����3333DDDD���L��L��L����D�����3333DDDDADAL�L��L�D����3333DDDDLA�L�L��L�D����3333DDDD�A���LLL�DD�����3333DDDD��������������������3333DDDD�DLDD�L�L�����3333DDDD���4���4��4|�4�|�4���43334DDDD"""������������������""""������������������������""""�������DA�A�A""""�������I�I�DI�II�""""������D""""������IADD���I""""��������D��""""�������I��I�I�I�""""�������A�D�II�I""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""wwwwwwwwwwwwwwwwww""""wwwwwwDGAD""""wwwwwGGtGwGw""""wwwwqADGAGwqGwq""""wwwwqDDDwwwq""""wwwwqAADqq""""wwwwqwqwAwAwqw""""wwwwqwAAAAqA""""wwwwwqwqDDAAAQ""""wwwwqqAqAqqA"""$www4www4www4www4www4www4UUUUUUUUUUUUUUUUUU333DDDAEEDUEUUEUUTEUUUUUU3333DDDDEUEUEUEUTEUTUUUU3333DDDDEUQEUQEUQEUQEUUDUUUU3333DDDDUUAUUUUUUTDDUUUU3333DDDDqTAUAAUDDDUUUU3333DDDDqUAUEEQUUDDUUUU3333DDDDADAAQAUEDUTUUUU3333DDDDQUQUUEQEUDDUUUU3333DDDDAAAQAQAQEDUDUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            