GST@�                                                            \     �                                               `(         ��5             �i  2�������J����������    ����        �      #    ����                                d8<n    �  ?     |�����  �
fD�
�L���"����D"� j   " B   J  jF�"    B�jl �  �
����
�"    
 �j,� B ��
  ��                                                                              ����������������������������������      ��    ??= 000 554 881                  

    

             ��� 44� � ���                 YYn 	         ::�����������������������������������������������������������������������������������������������������������������������������o=  0  o4   1  +      '           �                    	�  7�  V�  	�                  �  	          : �����������������������������������������������������������������������������                                ��  �       ��   @  #   �   �                                                                                'w w  YY	n  	�    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    T5I���K�	��)�Y|/�Db��D�N����hErG�s�+T0 k� ��A��AeA�s B1e 'Q  ��    �  mS�5I���[�	��) �Y|/�Db��D|N����`ErK�s�,T0 k� ��D��DeA�s B1e 'Q  /�    �  hS�5C���g�	��) �Y|/�Db��DtN����`D�O�s�,T0 k� ��E��EeA�s B1e 'Q  ��    �  cS�5C���o�	��) �Y|/�Db��DpN����\D�O�s�-T0 k� ��G��GeA�s B1e 'Q  ��    �  ^S�5C���w�	��* �	Y|/�Eb��DhN����XD�S�s�-T0 k� �xH�|HeA�s B1e 'Q  ��    �  ZS�5C�����	��* �	Y|/�Eb�DdN����TD�W�s�-T0 k� �lJ�pJeA�s B1e 'Q  ��    �  VS�5C�����	��* xY|/�Eb�DXN����PF[�s�.T0 k� �XM�\MeA�s B1e 'Q  ��    �  R��5C��s��	��+ pY|/�Eb�DPN��LF_�s�.T0 k� �LN�PNeA�s B1e 'Q  ��    �  P��5C�s��	��+ lY|/�Eb�	DHN��LFc�s�.T0 k� �4O�8OeA�s B1e 'Q  ��    �  N��5C�s��	��+ dY|/�Eb�DDN��HFg�s�.T0 k� �$N�(NeA�s B1e 'Q  ��    �  L��6C�së	��,XY|/�Eb�D4N��DFo�s�.T0 k� �M�MeA�s B1e 'Q  ��   �  J�6CРs˪	��,PY|/�Eb�Ab,N ��DFs�s|/T0 k� ��M� MeA�s B1e 'Q  ��    �  G�6CДsө	��-HY|/�Eb|Ab$N ��@D�w�x.T0 k� ��M��MeA�s B1e 'Q  ��    �  D�7CЈsۨ	�|-@Y|/�EbxAbN ��@
D�{�t.T0 k� ��M��MeA�s B1e 'Q  ��    �  A�7C�|s�	�x.<Y|/�ERtAbN {�@	D��t.T0 k� ��M��MeA�s B1e 'Q  ��    �  >�7C�|s�	�t.(Y|/�ERhE�N k�<D҇�l-T0 k� ��M��MeA�s B1e 'Q  ��    �  ;�8C�ts��	�p. Y|/�ER`E��N c�<Er��h-T0 k� ��M��MeA�s B1e 'Q  ��    �  8�8C�lt�	�l/Y|/�ER\E��N [�<Er��h,T0 k� ��M��MeA�s B1e 'Q  ��    �  5�8C�dd�	�h/Y|/�ERT!E��N S��<Er��d,T0 k� ��M��MeA�s B1e 'Q  ��    �  2�9C�\d�	�d/�Y|/�ERP#E��N K��@Er��d+T0 k� ��M��MeA�s B1e 'Q  ��    �  /�9C�Td�	�\/�Y|/�ERH%EA�N C��@ Er��`*T0 k� ��H��HeA�s B1e 'Q  ��    �   ,�:C�Dd'��T0��Y|/�C�<(EA�N7��C�Er��\)T0 k� ��D��DeA�s B1e 'Q  ��    � ! )�:C�<d+��P0��Y|/�C�8*EA�N/��G�D���3\(T0 k� ��B��BeA�s B1e 'Q  ��    � " &�:C�8 d3��H1o�Y|/�C�0,EA�N'��G�D���3\'T0 k� ��@��@eA�s B1e 'Q  ��7    � # $�x;C�0 d7��D1o�Y|/�C�(.EA�N��G�D���3\&T0 k� ��?��?eA�s B1e 'Q  ��7    � $ "�t;C�(!d?��@1o�Y|/�C�$/EA�M��K�D���3\%T0 k� ��>��>eA�s B1e 'Q  ��7    � %  �d;C�"dG��41o�Y|/�C�3EA�M��O�D���3\#T0 k� �l;�p;eA�s B1e 'Q �7    � % \<C�"dK��,2o�Y|/�C�4Ga�M���S�D���3`"T0 k� �`:�d:eA�s B1e 'Q ��?    � % T<C�#dS��(2o�Y|/�C�6Ga�L���W�D���3`!T0 k� �P9�T9eA�s B1e 'Q �?    � % L<C�#TO�@ 2	��Y|/�AR 8Ga�L_���[�A��3` T0 k� �D7�H7eA�s B1e 'Q �?    � % H<C��#TK�@3	��Y|/�AQ�9GaxL_���[�A���3`T0 k� �86�<6eA�s B1e 'Q ��?    � % @=C��$TK�@3	��Y|/�AQ�;GapL_���_�A���3dT0 k� �,5�05eA�s B1e 'Q ��?    � % 4=C��$TG�@3	��Y|/�AQ�<GalL_���c�A���3dT0 k� �4� 4eA�s B1e 'Q ��?    � % ,=C��%TC�@4	��Y|/�AQ�>GqdK_���g�A���3dT0 k� �2�2eA�s B1e 'Q ��?    � % $=E��%TC�@ 4	��Y|/�AQ�?Gq\K_���g�A���3dT0 k� �1�1eA�s B1e 'Q ��?    � % >E��&D?�O�5	ϜY|/�AQ�AGqTK_���k�A���3hT0 k� ��0��0eA�s B1e 'Q ��?    � % >E��&D;�O�5	ϘY|/�AQ�BGqLK_���o�A���3hT0 k� ��/��/eA�s B1e 'Q ��?    � % >E��'D7�O�6	ϔY|/�AQ�CGqHK_���o�A���3hT0 k� ��-��-eA�s B1e 'Q ��?    � % >E��'D3���6	ϐY|/�AQ�EG�@J_�� s�A���3hT0 k� ��,��,eA�s B1e 'Q ��?    � % �?E��(D/���7	όY|/�AQ�FG�8J_�� w�A���3lT0 k� ��+��+eA�s B1e 'Q ��?    � % �?E��)�+���8	��Y|/�AQ�HG�0J_�� w�A���3lT0 k� ��*��*eA�s B1e 'Q	 ��?    � % �?E��)�'���8	��Y|/�AQ�IG�,J_�� {�A���3lT0 k� ��(��(eA�s B1e 'Q	 ��?    � % �?E�*�#���9	��Y|/�AQ�JG�$J_�� �A���3lT0 k� ��'��'eA�s B1e 'Q	 ��?    � % �@E�+��O�:	��Y|/�AQ�KG� J_�� �A���3pT0 k� ��&��&eA�s B1e 'Q
 ��?    � % �@E�+��O�;	�|Y|/�AQ�MG�I_{� ��A���3pT0 k� ��%��%eA�s B1e 'Q
 ��?    � % �@E��,��O�;	�xY|/�AQ�NG�I_s� ��A���3pT0 k� �t#�x#eA�s B1e 'Q
 ��?    � % �@E��,��O�<	�xY|/�AQ�OG�I_k� ��A���3pT0 k� �h"�l"eA�s B1e 'Q ��?    � % �@E��-��O�=	�tY|/�AQ�PG�I_c� ��A�� 3tT0 k� �X!�\!eA�s B1e 'Q ��?    � % �AE��.��O�>	�tY|/�AQ�RG� I_[� ��A��3tT0 k� �L �P eA�s B1e 'Q ��?    � % �AE��/��?�?	�pY|/�AQ�SG��I_W� ��A��3tT0 k� �@�DeA�s B1e 'Q ��?    � % �AE��/��?�@	�pY|/�AQ�TG��H_O� ��A��3tT0 k� �0�4eA�s B1e 'Q ��?   � % �AE��0���?�B	�lY|/�AQ|UG��H_G� ��A��3tT0 k� �$�(eA�s B1e 'Q ��?    � % �AE��1���?�C	�lY|/�AQxVG��H_?� ��A��3xT0 k� ��eA�s B1e 'Q ��?    � % �BE�|2���?�D	�lY|/�AQtWG��H_7� ��A��3xT0 k� ��eA�s B1e 'Q ��?    � % "�BE�x3��?�E	�hY|/�AQpXG��H_/� ��A��	3x
T0 k� ��� eA�s B1e 'Q ��?    � % "xBFt4��?|G	�hY|/�AQhYG��H_'� ��A� 
3x
T0 k� ����eA�s B1e 'Q ��?    � % "pBFl6��?tH	�hY|/�AQdZG��H_� ��A�3x	T0 k� ����eA�s B1e 'Q ��?   � % "lBFh7��?pI	�hY|/�AQ`[G��G_� ��A�3|T0 k� ����eA�s B1e 'Q ��?    � % "dBFd8��?hK	�hY|/�AQ\\G��G_� ��A�3|T0 k� ����eA�s B1e 'Q ��?    � % "\CF`9�/dL	�hY|/�AQX]A �G_� ��A�3|T0 k� ����eA�s B1e 'Q ��?    � % "XCF\;ߞ/`N	�hY|/�AQT^A �G_� ��A�3|T0 k� ����eA�s B1e 'Q ��?    � % "PCFX<۟/XO	�hY|/�AQP_A �G^�� ��A�3|T0 k� ����eA�s B1e 'Q ��?    � % "HCFT=ן/TQ	�hY|/�AQL`A �G^�� ��A�3|T0 k� ����eA�s B1e 'Q ��?    � % DCFP?ӟ/PR	�hY|/�AQHaA �G^�� ��A�3�T0 k� ����eA�s B1e 'Q	 ��?    � % <CFL@Ӡ/LT	�hY|/�AQDbA �G^�� ��A�3�T0 k� �|��eA�s B1e 'Q	 ��?    � % 8DFLBϠ/HUOhY|/�AQ@cA �F^�� ��A�3�T0 k� �l
�p
eA�s B1e 'Q	 ��?    � % 0DE�HCˠ/DWOhY|/�AQ<dA �F^�� ��A�3�T0 k� �`	�d	eA�s B1e 'Q ��?    � % ,DE�DDǡ/@YOhY|/�AQ8eA �F^�� ��A�3�T0 k� �T�XeA�s B1e 'Q ��?    � % $DE�DFá/<ZOhY|/�AQ4fA �F^�� ��A�3�T0 k� �D�HeA�s B1e 'Q ��?    � %  DE�@Gá/8\OhY|/�AQ0gA �F^�� ��A�3�T0 k� �8�<eA�s B1e 'Q ��?    � % DE�@H��8] hY|/�AQ,gA �F^�� ��A�3� T0 k� �,�0eA�s B1e 'Q ��?    � % EE�@J��4_ hY|/�AQ(hA �F^�� ��A�3� T0 k� � �$eA�s B1e 'Q ��?    � % �EE�@K��0a hY|/�AQ$iA �F^�� ��A� 3��T0 k� ��eA�s B1e 'Q ��?    � % �EE�<L��0b hY|/�AQ jA �F^�� ��A� 3��T0 k� � � eA�s B1e 'Q ��?   � % �EB�<M��,d hY|/�AQkA �E^�� ��A�$3��T0 k� ������eA�s B1e 'Q ��?    � % ��EB�<O��,e ohY|/�AQkA �E^�� ��A�$3��T0 k� ������eA�s B1e 'Q ��?    � % ��EB�<P��(g ohY|/�AQlA |E^�� ��A�$3��T0 k� ������eA�s B1e 'Q ��?    � % �EB�<Q��(h ohY|/�AQmA xE^�� ��A�( 3��T0 k� ������eA�s B1e 'Q ��?    � % �EB�<R��$j ohY|/�AQnA tE^�� ��A�(!3��T0 k� ������eA�s B1e 'Q ��?    � % �FB�@S��$k ohY|/�AQnA pE^{� ��A�,"3��T0 k� ������eA�s B1e 'Q ��?    � % �FB�@T��  l�hY|/�AQoA pE^s� ��A�,"3��T0 k� ������eA�s B1e 'Q ��?    � % �FB�@V��  n�hY|/�AQpA lE^k� ��A�,#3��T0 k� ������eA�s B1e 'Q ��?    � % �FB�DW��  o�l Y|/�AQqA hE^g� ��A�0$3��T0 k� ������eA�s B1e 'Q  ��?    � % �FB�DX�� p�l Y|/�AQ qA dE^_� ��A�0%3��T0 k� ������eA�s B1e 'Q  ,�?    � % !�FB�HY�� r�l Y|/�AP�rA `D^W� ��A�0&3��T0 k� �w��{�eA�s B1e 'Q  ��?    � % !�FB�HZ�� s�l Y|/�AP�sA \D^O� ��A�4&3��T0 k� �k��o�eA�s B1e 'Q  ��?    � % !�FB�L[�� t�p!Y|/�AP�sA \D^K� ��A�4'3��T0 k� �_��c�eA�s B1e 'Q  ��?    � % !�GB�L\�� v�p!Y|/�AP�tA XD^C� ��A�4(3��T0 k� �O��S�eA�s B1e 'Q ��?    � % !�GB�P]�� wp!Y|/�AP�tA TD^;� ��A�8(3��T0 k� �C��G�eA�s B1e 'Q ��?    � % !�GB�T^�� xt"Y|/�AP�uA PD^3� ��A�8)3��T0 k� �7��;�eA�s B1e 'Q ��?    � % !�GB�X_�� yt"Y|/�AP�vA PD^/� ��A�8*3��T0 k� �+��/�eA�s B1e 'Q ��?    � % !�GB�X`�� zx#Y|/�AP�vA LD^'� ��A�<*3��T0 k� ����eA�s B1e 'Q ��?   � % !�GB�\a�� {x#Y|/�AP�wA HD�� ��A�<+3��T0 k� ����eA�s B1e 'Q ��?    � % �GB�`b�� }|$Y|/�AP�xA DD�� ��A�<,3��T0 k� ����eA�s B1e 'Q ��?    � % �GB�db�� ~|$Y|/�AP�xA DD�� ��A�@,3��T0 k� ������eA�s B1e 'Q ��?    � % �GB�hc�� �%Y|/�AP�yA @D�� ��A�@-3��T0 k� ������eA�s B1e 'Q ��?    � % �GB�ld�� ��%Y|/�AP�yA <D�� ��A�@.3��T0 k� ������eA�s B1e 'Q ��?    � % �HB�te� ��&Y|/�AP�zA <C]�� ��A�@.3��T0 k� ������eA�s B1e 'Q ��?    � % �HB�xf� �'Y|/�AP�zA 8C]�� ��A�D/3��T0 k� ������eA�s B1e 'Q ��?    � % �HB�|g{� �'Y|/�AP�{A 4C]�� ��A�D03��T0 k� ������eA�s B1e 'Q ��?    � % �HBπh�{� �(Y|/�AP�{A 4C]�� ��A�D03��T0 k� ������eA�s B1e 'Q ��?    � % �HBψh�{� �)Y|/�AP�|A 0C]�� ��A�D13��T0 k� ������eA�s B1e 'Q ��?    � % �HBόi�w�  ~�)Y|/�AP�|A ,C]�� ��A�H13��T0 k� ������eA�s B1e 'Q ��?    � % �|HBϐj�w�  ~�*a�/�AP�}A ,C��� ��A�H23��T0 k� �����eA�s B1e 'Q ��?    � % �xHBϘk�s�  ~��+a�/�AP�}A (Cݿ� ��A�H23��T0 k� �s��w�eA�s B1e 'Q ��?    � % �tHBϜl�s� �~��+a�/�AP�~A (Cݳ� ��A�H33��T0 k� �k��o�eA�s B1e 'Q ��8    � % �lHE��l�o� �}��,a�/�AP�~A $Cݧ� ��A�L33��T0 k� �c��g�eA�s B1e 'Q ��8    � % �hHE��m�o� �}��-a�/�AP�A  Cݛ� ��A�L43��T0 k� �W��[�eA�s B1e 'Q ��8    � % �dIE��n�k� �}��-a�/�AP�A  Cݏ� ��A�L43��T0 k� �O��S�eA�s B1e 'Q  ��8    � % �\IE��n�k� �}��.a�/�AP��A C�� ��A�L53��T0 k� �C��G�eA�s B1e 'Q  ��8    � % �XIE��o�g� �}��.a�/�AP�A C�s� ��A�P53��T0 k� �7��;�eA�s B1e 'Q  ��8    � % �TIE��p�g� �|��/a�/�AP�A C�g� ��A�P63��T0 k� �+��/�eA�s B1e 'Q  /�8    � % �LIE��q�c� �|��/a�/�AP�A C�[� ��A�P63��T0 k� ���#�eA�s B1e 'Q  ��8    � % �HIE��q�_� �|��0a�/�AP�A C�S� ��A�P73��T0 k� ����eA�s B1e 'Q  ��8    � % �@IE��r�[� �|��1Y|/�AP�A B�G� ��A�T73��T0 k� ����eA�s B1e 'Q  ��8    � % �<IE��s�[� �|ϰ1Y|/�AP�~A B�;� ��A�T83��T0 k� ������eA�s B1e 'Q  ��8   � % �4IE��s�W� �{ϴ2Y|/�AP�~A B�/� ��A�T83��T0 k� ������eA�s B1e 'Q  ��8    � % �,IE��t�S� �{ϴ2Y|/�AP�~A B�#� ��A�T93��T0 k� ������eA�s B1e 'Q  ��8    � % �(IE��t�O� �{ϸ3Y|/�AP�~A B�� ��A�T93��T0 k� ������eA�s B1e 'Q  ��8    � % � IE��u�K� �{ϸ3Y|/�AP�}A B�� ��A�X:3��T0 k� ������eA�s B1e 'Q  ��8    � % �IE�u�G� �{ϼ4Y|/�AP�}A B�� ��A�X:3��T0 k� ������eA�s B1e 'Q  ��8    � % AJE�u�C� �zϼ4Y|/�AP�}A B��� ��A�X;3��T0 k� ������eA�s B1e 'Q  ��8    � % AJE�v�?� �z��5Y|/�AP�}A B��� ��A�X;3��T0 k� ������eA�s B1e 'Q  ��8    � % AJE�v�;� �z��5Y|/�AP�}A  B��� ��A�X;3��T0 k� ������eA�s B1e 'Q  ��8    � % @�JE�$v�7� �z��6Y|/�AP�|A  B��� ��A�\<3��T0 k� ������eA�s B1e 'Q  ��8    � % @�JE�,v�3� �z��6a�/�AP�|A  B��� �A�\<3��T0 k� ������eA�s B1e 'Q  ��8    � % @�KE�4v�/� �z��6a�/�AP�|A�B��� �A�\=3��T0 k� ������eA�s B1e 'Q  ��8    � % @�KE�<v�+� �y��7a�/�AP�|A�B��� �A�\=3��T0 k� ������eA�s B1e 'Q  ��8    � % @�LE�Dv�'� �y��7a�/�AP�|A�Bܷ� ��A�\=3��T0 k� �w��{�eA�s B1e 'Q  ��8    � % @�LE�Lv�#� �y��7a�/�AP�{A�B\�� ��A�\>3��T0 k� �o��s�eA�s B1e 'Q  ��8    � % @�LE�Tv�� �y��7a�/�AP�{A�B\�� ��A�`>3��T0 k� �g��k�eA�s B1e 'Q  ��8    � % ��ME�\v�� �y��7a�/�AP�{A�C\�� ��A�`>3��T0 k� �[��_�eA�s B1e 'Q  ��8    � % ��NE�\v�� �y��7a�/�AP�{A�C\�� ��A�`?3��T0 k� �S��W�eA�s B1e 'Q  ��8    � % ��NE�`u�� �x��7a�/�AP�{A�C\�� ��A�`?3��T0 k� �K��O�eA�s B1e 'Q  ��8    � % ��OE�dt�� �x��7a�/�AP�{A�C\�� ��A�`?3��T0 k� �C��G�eA�s B1e 'Q  ��8    � % ��OE�ht�� �x��7a�/�AP�{A�D\{� ��A�`@3��T0 k� �;��?�eA�s B1e 'Q  ��8    � % 	p�OE�hs��� �x��8Y|/�AP�|A�D\s� ��A�d@3��T0 k� �3��7�eA�s B1e 'Q  ��8    � % 	p�PE�lr��� �x��8Y|/�AP�|A�D\k� ��A�d@3��T0 k� �+��/�eA�s B1e 'Q  ��8    � % 	p�PE�pq��� �x��8Y|/�AP�|A�D\c� ��A�dA3��T0 k� �#��'�eA�s B1e 'Q  ��8    � % 	p�PE�tp��� �x��8Y|/�AP�|A�D\[� ��A�dA3��T0 k� ����eA�s B1e 'Q  ��8    � % 	p�PE�to��� �w��8Y|/�AP�|A�E\S� ��A�dA3��T0 k� ����eA�s B1e 'Q  ��8    � % 	��QE�xn��� �w��8Y|/�AP�|A�E\O� ��A�dB3��T0 k� ����eA�s B1e 'Q  ��8    � % 	��QE�xm�����w��8Y|/�AP�|A�E\G� ��A�dB3��T0 k� ����eA�s B1e 'Q  ��8    � % 	�|QE�|l�����w��8Y|/�AP�|A�E\?� ��A�hB3��T0 k� �����eA�s B1e 'Q  ��8    � % 	�xQE�|k�����w��8Y|/�AP�|A�E\7� ��A�hC3��T0 k� ������eA�s B1e 'Q  ��8    � % 	�pQE�|j�����w��8Y|/�AP�}A�F\/� ��A�hC3��T0 k� ������eA�s B1e 'Q  ��8    � % 	plQE��i�����w��9Y|/�AP�}A�F\+� ��A�hC3��T0 k� ������eA�s B1e 'Q  ��8    � % 	phQE��h»���w��9Y|/�AP�}A�F\#� ��A�hD3��T0 k� ������eA�s B1e 'Q  ��8    � % 	pdQE��g³���w��9Y|/�AP�}A�F\� ��A�hD3��T0 k� ������eA�s B1e 'Q  ��8    � % 	p`QK��f¯���v��9Y|/�AP�}A�F\� �A�hD3��T0 k� ������eA�s B1e 'Q  ��8    � % 	p`QK��e§���v��9Y|/�AP�}A�G\� �A�hD3��T0 k� ������eA�s B1e 'Q  ��8    � % 	�\QK��d�����v��9Y|/�AP�}A�G\� �A�lE3��T0 k� ������eA�s B1e 'Q  ��8    � % 	�XQK��b�����v��9Y|/�AP�}A�G\� �A�lE3��T0 k� ������eA�s B1e 'Q  ��8    � % 	�TQK��a�����v��9Y|/�AP�}A�G[�� �A�lE3��T0 k� ������eA�s B1e 'Q  ��8    � % 	�TQK��`�����v��9Y|/�AP�}A�G[�� �A�lE3��T0 k� ������eA�s B1e 'Q  ��8    � % 	�PQK��_�����v��9Y|/�AP�}A�G[�� �A�lF3��T0 k� ������eA�s B1e 'Q  ��8    � % 	pLQK��^����v��9Y|/�AP�~A�H[�� �A�lF3��T0 k� ������eA�s B1e 'Q  ��8    � % 	pLQK��]�w���v��9Y|/�AP�~A�H[�� �A�lF3��T0 k� ������eA�s B1e 'Q  ��8    � % 	pHQK��\�o���u��:Y|/�AP�~A�H[�� �A�lF3��T0 k� ������eA�s B1e 'Q  ��8    � % 	pHQK��[�g���u��:Y|/�AP�~A�H[�� �A�pG3��T0 k� ������eA�s B1e 'Q  ��8    � % 	pHQK��Z�c���u��:Y|/�AP�~A�H[�� �A�pG3��T0 k� ������eA�s B1e 'Q  ��8    � % 	�DQK��Y�[���u��:Y|/�AP�~A�H[�� �A�pG3��T0 k� ������eA�s B1e 'Q  ��8    � % 	�DQK��Y�S���u��:Y|/�AP�~A�I[�� �A�pG3��T0 k� ������eA�s B1e 'Q  ��8    � % 	�DQL �X�K���u��:Y|/�AP�~A�I[�� �A�pH3��T0 k� �����eA�s B1e 'Q  ��8    � % 	�DQL �W�G���u��:Y|/�AP�~A�I[�� �A�pH3��T0 k� �{���eA�s B1e 'Q  ��8    � % 	�@QL �V�?���u��:Y|/�AP�~A�I[�� �A�pH3��T0 k� �w��{�eA�s B1e 'Q  ��8    � % 	p@QL �U�7���u��;Y|/�AP�~A�I[�� �A�pH3��T0 k� �s��w�eA�s B1e 'Q  ��8    � % 	p@QL �T�/���u��;Y|/�AP�~A�I[�� �A�pH3��T0 k� �k��o�eA�s B1e 'Q  *�8    � % 	p@QL �S�+���u��;Y|/�AP�~A�I[�� �A�pI3��T0 k� ;k��o�eA�s B1e 'Q  ��8    � % 	p@QL �S�#���u��;Y|/�AP�A�J[�� �A�tI3��T0 k� ;c��g�eA�s B1e 'Q  *�8    � % 	p@QL �R����t��<Y|/�AP�A�J[�� �A�tI3��T0 k� ;c��g�eA�s B1e 'Q  .�8    � %  @QL �Q����t��<Y|/�AP�A�J[�� �A�tI3��T0 k� ;_��c�eA�s B1e 'Q  ��8    � %  @QL �P����t��<Y|/�AP�A�J[�� �A�tI3��T0 k� ;_��c�eA�s B1e 'Q  ��8    � %  @QL �O����t��<Y|/�AP�A�K[�� �A�tJ3��T0 k� �_��c�eA�s B1e 'Q  ��8    � %  @QL �N�� ��t�<Y|/�AP�A�K[�� �A�tJ3��T0 k� �c��g�eA�s B1e 'Q  ��8    � %  @QL �M����t�<Y|/�AP�A�L[�� �A�tJ3��T0 k� �c��g�eA�s B1e 'Q  ��8    � %  @QL �L����t�=Y|/�AP�A�L[�� �A�tJ3��T0 k� �c��g�eA�s B1e 'Q  ��8    � %  @QL �L����t�=Y|/�AP�A�L[�� �A�tK3��T0 k� �c��g�eA�s B1e 'Q  ��8    � %  @QL �K����t�=Y|/�AP�A�M[�� �A�tK3��T0 k� �c��g�eA�s B1e 'Q  ��8    � %  @QL �J����t�=Y|/�AP�A�M[�� �A�xK3��T0 k� �c��g�eA�s B1e 'Q  ��8    � % P@QL �J��
��t�=Y|/�AP�A�N[�� �A�xK3��T0 k� �c��g�eA�s B1e 'Q  ��8    � % P@QL �I����t�>Y|/�AP�A�N[�� �A�xK3��T0 k� �g��k�eA�s B1e 'Q  ��8    � % P@QL �H����t�>Y|/�AP�A�N[�� �A�xK3��T0 k� �g��k�eA�s B1e 'Q  ��8    � % P@QL �G����s�>Y|/�AP�A�O[�� �A�xL3��T0 k� �g��k�eA�s B1e 'Q  ��8    � % P@QL �G����s�?Y|/�AP��A�O[�� �A�xL3��T0 k� �g��k�eA�s B1e 'Q  ��8    � % P@QL �F����s�?Y|/�AP�A�P[�� �A�xL3��T0 k� �k��o�eA�s B1e 'Q  ��8    � % P@QL �F����s�@Y|/�AP�A�P[�� �A�xL3��T0 k� �k��o�eA�s B1e 'Q  ��8    � % P@QL �E����s�@Y|/�AP�A�P[�� �A�xL3��T0 k� �k��o�eA�s B1e 'Q  ��8    � % P@QL �D����s�@Y|/�AP�A�Q[�� �A�xL3��T0 k� �k��o�eA�s B1e 'Q  ��8    � % P@QL �D����s�@Y|/�AP�~A�R[�� �A�xL3��T0 k� �k��o�eA�s B1e 'Q  ��8    � % P@QL �C����s�AY|/�AP�~A�R[�� �A�xM"s��T0 k� �o��s�eA�s B1e 'Q  ��8    � % P@QL �C����s�AY|/�AP�~A�S[�� �A�xM"s��T0 k� �o��s�eA�s B1e 'Q  ��8    � % P@QL �B�x��s�BY|/�AP�~A�S[�� �A�|M"s��T0 k� �o��s�eA�s B1e 'Q  ��8    � % P@QL �A�p ��s�BY|/�AP�}A�S[�� �A�|M"s��T0 k� �o��s�eA�s B1e 'Q  ��8    � % P@QL �A�l"��s�BY|/�AP�}A�T[�� �A�|M"s��T0 k� �o��s�eA�s B1e 'Q  ��8    � % P@QL �@�d#��s/�BY|/�AP�}A�U[�� �A�|M"s��T0 k� �s��w�eA�s B1e 'Q  ��8    � % P@QL �@�\%��s  CY|/�AP�}A�U[�� �A�|M"s��T0 k� �s��w�eA�s B1e 'Q  ��8    � % P@QL �?�T'��s  DY|/�AP�}A�V[�� �A�|N"s��T0 k� �s��w�eA�s B1e 'Q  ��8    � % @QL �?�P(��s DY|/�AP�|A�V[�� �A�|N"s��T0 k� �s��w�eA�s B1e 'Q  ��8    � % @QL �>�H*��s EY|/�AP�|A�W[�� �A�|N"s��T0 k� �s��w�eA�s B1e 'Q  ��8    � % @QL �>�@,��s EY|/�AP�|A�W[�� �A�|N"s��T0 k� �w��{�eA�s B1e 'Q  ��8    � % @QL �=�8-��s FY|/�AP�|A�X[�� �A�|N3��T0 k� �w��{�eA�s B1e 'Q  ��8    � % @QL �=�4/ �r FY|/�AQ |A�X[�� �A�|N3��T0 k� �w��{�eA�s B1e 'Q  ��8    � % DQK�<�,1 �r FY|/�AQ {A�X[�� �A�|N3��T0 k� �w��{�eA�s B1e 'Q  ��8    � % DRK�<�$3 �r GY|/�AQ {A�Y[�� �A�|N3��T0 k� �w��{�eA�s B1e 'Q  ��8   � % DRK�;� 4 �r GY|/�AQ {A�Y[�� �A�|O3��T0 k� �{���eA�s B1e 'Q  ��8    � % HRK�;�6 �r�GY|/�AQ {A�Z[�� �A�|O3��T0 k� �{���eA�s B1e 'Q  ��8    � % HSK�:�8 �r�HY|/�AQ {A  Z[�� �A�|O3��T0 k� �{���eA�s B1e 'Q  ��8    � %  LSK�:�9 �r�HY|/�AQzA  [[�� �A�|O3��T0 k� �{���eA�s B1e 'Q  ��8    � %  LSEР:�; �r�IY|/�AQzA  [[�� �A�O3��T0 k� �{���eA�s B1e 'Q  ��8    � %  PTEМ9��= �r�IY|/�AQzA  \[�� �A�O3��T0 k� �{���eA�s B1e 'Q  ��8    � %  PTEМ9��> �r� IY|/�AQzA  \[�� �A�O3��T0 k� �����eA�s B1e 'Q  ��8    � %  TUEМ8��@ �r� JY|/�AQzA  \[�� �A�O"���T0 k� �����eA�s B1e 'Q  ��8    � %  TUEМ8��A �r� JY|/�AQzA  ][�� �A�P"���T0 k� �����eA�s B1e 'Q  ��8    � %  TUEМ8��C �r�$JY|/�AQyA  ][�� �A�P"���T0 k� �����eA�s B1e 'Q  ��8    � %  XVEИ7��E �r�$JY|/�AQyA  ][�� �A�P"���T0 k� �����eA�s B1e 'Q  ��8    � %  XVEИ7��F �r�$JY|/�AQyA  ^[�� �A�P"���T0 k� �����eA�s B1e 'Q  ��8    � % \VEД6��H �r�$JY|/�AQyA  ^[�� �A�P"���T0 k� �����eA�s B1e 'Q  ��8    � % \WEД6��I �r $JY|/�AQyA _[�� �A�P"���T0 k� ������eA�s B1e 'Q  ��8    � % \WE��6�J �r $JY|/�AQyA _[�� �A�P"���T0 k� ������eA�s B1e 'Q  ��8    � % `WE��5�L �r $JY|/�AQyA _[�� �A�P"���T0 k� ������eA�s B1e 'Q  ��8    � % `XE��5�M �r $JY|/�AQxA `[�� �A�P"���T0 k� ������eA�s B1e 'Q  ��8    � % dXE��5�O �r $JY|/�AQxA `[�� �A�P"���T0 k� ������eA�s B1e 'Q  ��8    � % dXE��5�O �r (KY|/�AQxA `[�� �A�P3��T0 k� ������eA�s B1e 'Q  ��8    � % `YE��5�O �r (KY|/�AQxA a[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % `ZE��5�P �r (KY|/�AQxA a[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % \[E��5�Q �r (KY|/�AQxA a[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % \\E�|5�Q �r (KY|/�AQxA b[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % X\E�x5�R �r ,KY|/�AQwA b[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % X]E�x5�S �r,LY|/�AQwA b[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % X]LPt5�S �r,LY|/�AQwA c[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % T^LPp5�T �q,LY|/�AQwA c[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % T_LPp5�T �q0MY|/�AQwA c[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % T_LPl5�U �q0MY|/�AQwA c[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % T_LPl6�U �q0MY|/�AQwA d[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % T`LPh6�V �q4NY|/�AQwA d[�� �A�Q3��T0 k� ������eA�s B1e 'Q  ��8    � % P`LPd6�V �q4NY|/�AQwA d[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % PaLPd6 �V �q4NY|/�AQvA e[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % PaLP`6 �W �q4NY|/�AQvA e[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % PbLP`6 �W �q4NY|/�AQvA e[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % PbLP\6 �W �q 4NY|/�AQvA e[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % PbLP\6 �W �q 4NY|/�AQvA f[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % LcL`X6 |W �q 4NY|/�AQvA f[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % LcL`T6 |W �q 4NY|/�AQvA f[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % LcL`T6 |W �q 4NY|/�AQvA f[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % LcL`P6 |X �q �4NY|/�AQvA g[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % LcL`P6 |X �q �4NY|/�AQvA g[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % LdL`L7 |X �q �4NY|/�AQuA g[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % LdL`L7 |X �q �4NY|/�AQuA g[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % LdL`H7 |X �q �4NY|/�AQuA h[�� �A�R3��T0 k� ������eA�s B1e 'Q  ��8    � % LdL`H7 |Y �q �4NY|/�AQuA h[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % LdL`D7 |Y �q �4NY|/�AQuA h[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % LdL`D7 |Y �q�4NY|/�AQuA h[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`D7 |Y �q�4NY|/�AQuA h[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`@7 |Y �q�4NY|/�AQuA i[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`@7 |Y �q�4NY|/�AQuA i[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`<7 |Y �q�4NY|/�AQuA i[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`<7 |Y �q�4NY|/�AQuA i[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`87 |Y �q�4NY|/�AQuA j[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`87 |Y �q�4NY|/�AQtA j[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`87 |Y �q�4NY|/�AQtA j[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`47 |Y �q�4NY|/�AQtA j[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`48 |Y �q�4NY|/�AQtA j[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`08 |Y �q�4NY|/�AQtA j[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`08 |Y �q�4NY|/�AQtA k[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`08 |Y �q�4NY|/�AQtA k[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`,8 |Y �q�4NY|/�AQtA k[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`,8 |Y �q�4NY|/�AQtA k[�� �A�S3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`,8 |Y �q�4NY|/�AQtA k[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`(8 |Y �q�4NY|/�AQtA l[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`(8 |Y �q�4NY|/�AQ tA l[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`(8 |Y �q�4NY|/�AQ tA l[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`$8 |Y �q�4NY|/�AQ tA l[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`$8 |Y �q�4NY|/�AQ tA l[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`$8 |Y �q�4NY|/�AQ tA l[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL` 8 |Y �q�4NY|/�AQ sA l[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL` 8 |Y �q�4NY|/�AQ sA m[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL` 8 |Y �q�4NY|/�AQ sA m[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`8|Y �q�4NY|/�AQ sA m[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`8|Y �q�4NY|/�AQ sA m[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`9|Y �q�4NY|/�AQ sA m[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`9|Y �q�4NY|/�AQ sA m[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdL`9|Y �q�4NY|/�AQ sA n[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdLP9|Y �q�4NY|/�AQ sA n[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdLP9|Y �q�4NY|/�AQ sA n[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdLP9P|Y �q�4NY|/�AQ sA n[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdLP9P|Y �q�4NY|/�AQ$sA n[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdLP9P|Y �q�4NY|/�AQ$sA n[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdLP9P|Y �q�4NY|/�AQ$sA n[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdD�9P|Y �q�4NY|/�AQ$sA n[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdD�9P|Y �q�4NY|/�AQ$sA o[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8   � % PLdD�9P|Y �q�4NY|/�AQ$sA o[�� �A�T3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdD�:P|Y �q�4NY|/�AQ$sA o[�� �A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdD�:P|Y �q�4NY|/�AQ$sA o[�� �A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdD�:P|Y �q�4NY|/�AQ$sA o[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdD�;P|Y �q�4NY|/�AQ$sA o[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdD�;P|Y �q�4NY|/�AQ$rA o[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdD�<P|Y �q�4NY|/�AQ$rA o[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdD�=P|Y �q�4NY|/�AQ$rA o[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE�=P|Y �q�4NY|/�AQ$rA p[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE�>P|Y �q�4NY|/�AQ$rA p[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE�?P|Y �q�4NY|/�AQ$rA p[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE�@P|Y �q�4NY|/�AQ$rA p[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE�@P|Y �q�4NY|/�AQ$rA p[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE�AP|Y �q�4NY|/�AQ$rA p[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdF BP|Y �q�4NY|/�AQ$rA p[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdF CP|Y �q�4NY|/�AQ(rA p[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � %  LdF CP|Y �q�4NY|/�AQ(rA p[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � %  LdF  DP|Y �q�8NY|/�AQ(rA p[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � %  LdF  EP|Y��q�8OY|/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � %  LdD� FP|Y��q�8OY|/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � %  LdD� GP|Y��q�8OY|/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � %  LdD� GP|Y��q�<OY|/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � %  LdD� HP|Y��q�<OY|/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � %  LdD� IP|Y��q�<OY|/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � %  LdF  IP|Y��q�<OY|/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdF  IP|Y��q�<Oa�/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdF  IP|Y��q�<Pa�/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdF  JP|Y��q�@Pa�/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdF  KP|Y��q�@Pa�/�AQ(rA q[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE� LP|Y��q�@Pa�/�AQ(rA r[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE� LP|Y��q�@Pa�/�AQ(rA r[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE� MP|Y��q�@Pa�/�AQ(rA r[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE� NP|Y��q�@Pa�/�AQ(rA r[�� #�A�U3��T0 k� ������eA�s B1e 'Q  ��8    � % LdE� NP|Y��q �@Pa�/�AQ(rA r[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB� NP|Y��q �@Pa�/�AQ(rA r[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB� OP|Y��q �@Pa�/�AQ(rA r[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB� OP|Y��q �@PY|/�AQ(rA r[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB� OP|Y��q �@PY|/�AQ(rA r[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB� OP|Y��q �DPY|/�AQ(rA r[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB� OP|Y��q �DPY|/�AQ(rA r[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB� PP|Y��q �DPY|/�AQ(rA r[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB� PP|Y��q �DPY|/�AQ(rA r[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�QP|Y��q �DPY|/�AQ,rA r[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�QP|Y��q �DPY|/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�RP|Y��q �DPY|/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�RP|Y��q �DPY|/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�SP|Y��q �DPY|/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�SP|Y��q �DPa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�SP|Y��q �DPa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�TP|Y��q �DOa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�TP|Y��q �DOa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�UP|Y��q �DOa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�UP|Y��q �DOa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�VP|Y��q �DOa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�VP|Y��q �DOa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�VP|Y��q �DOa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�WP|Y��q �DOa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�WP|Y��q �DOa�/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�WP|Y��q �DOY|/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�XP|Y��q �DOY|/�AQ,qA s[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�XP|Y��q �DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�XP|Y��q �DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�XP|Y��q �DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�XP|Y��q DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q�DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q�DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q�DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q�DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q�DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q�DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q�DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q�DOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % PLdB�YP|Y��q�HOY|/�AQ,qA t[�� #�A�V3��T0 k� ������eA�s B1e 'Q  ��8    � % �Dr��R�A�)A��Y|/�IB�@�hr�;���P���c��T0 k� �#��'�eA�s B1e 'Q ��    ��� ��Dr��R�A�)A��Y|/�IB�@�hr�;���P���c��T0 k� �'��+�eA�s B1e 'Q ��    ��� ��Dr��RߒA�)A��Y|/�IB��@�hr�;���P���c��T0 k� �/��3�eA�s B1e 'Q ��    ��� ��Dr��RےA�) ��Y|/�I2��@�hq�?���P���c��T0 k� �7��;�eA�s B1e 'Q ��    ��� ��Dr��BגA�) ��Y|/�I2��CBhq�?���P���c��T0 k� �;��?�eA�s B1e 'Q ��    ��� ��Or��BϒA�) ��Y|/�I2��CBhq�G���P�w�c��T0 k� �K��O�eA�s B1e 'Q ��    ��� ��Or��B˒A�) ��Y|/�I2��CBhp�K����Pro�c��T0 k� �O��S�eA�s B1e 'Q ��    ��� ��Or��BǒA�) a��Y|/�IB��CBhp�K����Prk�c��T0 k� �W��[�eA�s B1e 'Q ��    ��� ��Or��BÒA�) a��Y|/�IB��E"ho�O����Prc�c��T0 k� �_��c�eA�s B1e 'Q ��    ��� �� Or��B�� �) a��Y|/�IB��E"ho�O����Pr_�3��T0 k� �c��g�eA�s B1e 'Q ��    ��� �� Or��B�� �) a��Y|/�IB��E"hn�O����Pr[�3��T0 k� �k��o�eA�s B1e 'Q  ��    ��� �� Or��B�� �) a��Y|/�IB��E"hm�O���IrS�3��T0 k� �p�teA�s B1e 'Q  ��    ��� ��!Or��B�� �)A��Y|/�I2��E"hm�O���IrS�3��T0 k� �t�xeA�s B1e 'Q  ��    ��� ��!Or��B�� �)A��Y|/�I2��E"ll�S���IrO�3��T0 k� �|
��
eA�s B1e 'Q  /�    ��� ��"Or��B�� a�)A��Y|/�I2��E"lk�S���IrK�3��T0 k� ����eA�s B1e 'Q  ��    ��� ��"Or��B�� a�)A��Y|/�I2��E"lk�W���IrG�3�T0 k� ����eA�s B1e 'Q  ��    ��� ��"Or��B�� a�)A��Y|/�I2��E"lj�[�"��IrC�3�T0 k� ����eA�s B1e 'Q  ��    ��� ��#Or��B�� a�)A��Y|/�IB��E"pi�[�"��I�?�3�T0 k� ����eA�s B1e 'Q  ��    ��� ��#Or��B�� a�)A��Y|/�IB��E"phB_�"��I�;��T0 k� ����eA�s B1e 'Q  ��    ��� ��$Or��B�� a�)A��Y|/�IB��E"tfB_�"��I�3��T0 k� ��'��'eA�s B1e 'Q  ��    ��� ��$Or��B�� �)A��Y|/�IB��E"xfB_�#�I�3��	T0 k� ��,��,eA�s B1e 'Q  ��    ��� �$Or��B�� �)A��Y|/�I2��E"xeB_�#�Ir/��T0 k� ��0��0eA�s B1e 'Q  �    ��� �%Or��B�� �)Q��Y|/�I2��E"|dB_�#�Ir+��T0 k� ��+��+eA�s B1e 'Q ��    ��� �%Or��B�� �)Q��Y|/�I2��E"|cB_�#�Ir+�"3�T0 k� ��'��'eA�s B1e 'Q ��    ��� �%Or��B�� �)Q��Y|/�I2��E"�bB_��Ir'�"3�T0 k� ��"��"eA�s B1e 'Q ��    ��� ��&Or��B�� �)Q��Y|/�I2��E�aB_��Ir#�"3�T0 k� ����eA�s B1e 'Q ��    ��� ��&Or��B� �)Q��Y|/�@b��E�`B_��I�#�"3�T0 k� ����eA�s B1e 'Q $�    ��� ��&Or��B� �)Q��Y|/�@b��E�_B_��I��"3�T0 k� � �eA�s B1e 'Q ��    ��� ��'Or��w� �)Q��Y|/�@b��E�]_��I��)s�T0 k� ��eA�s B1e 'Q ��    ��� #�'Or{��s� �)Q��Y|/�@b��B��\_��#�I��)s�T0 k� ��eA�s B1e 'Q ��    ��� #�(Eb{��o� �)Q��Y|/�E��B��[_��'�Ir�)s�T0 k� � �$eA�s B1e 'Q ��    ��� #�(Ebw��k� �)Q��Y|/�E��B��Z_��'�Ir�)s�T0 k� �$�(eA�s B1e 'Q ��    ��� #�)Ebw��k� �)a��Y|/�E��B��Y_��+�Ir�)s�T0 k� �(�,eA�s B1e 'Q ��    ��� #�*Ebs��c� �)a��Y|/�E��B��W_��7�Ir�)s�T0 k� �,�0eA�s B1e 'Q ��    ��� �*Ebo��_� �)a��Y|/�E��B��VR_��;�I��)s�T0 k� �0�4eA�s B1e 'Q ��    ��� �+Ebk��[� a�)a��Y|/�E��B��VR_��?�I��)s�T0 k� �0�4eA�s B1e 'Q ��    ��� �,Ebk��W� a�)���Y|/�E���B��UR_��C�I��)s�T0 k� �0�4eA�s B1e 'Q ��    ��� �,Ebg��W� a�)���Y|/�E���B��TR_��G�I��)s�T0 k� �4�8eA�s B1e 'Q ��    ��� �-Eb_�2W� a�)���Y|/�E�ïB��S�[��S�I��)s�T0 k� �4�8eA�s B1e 'Q ��    ��� �.Eb_�2S� ��)���Y|/�E�ǯB��R�[��W�Ir�)s�T0 k� �4�8eA�s B1e 'Q  ��    ��� �.Eb[�2S� ��)���Y|/�E�˯B��R�W��[�Ir�)s�T0 k� �4�8eA�s B1e 'Q  ��    ��� ��/EbW�2S� ��)���Y|/�E�ϯB��Q�W��_�Ir�)s�T0 k� �4�8eA�s B1e 'Q  .�    ��� ��/EbS�2O� ��)���Y|/�E�ӰB��Q�S��g�Ir�)s�T0 k� �4�8eA�s B1e 'Q  ��    ��� ��/EbO�"O� ��)���Y|/�ErװB��P�S��k�Ir�)s�T0 k� �4�8eA�s B1e 'Q  ��    ��� ��0EbG�"O��)���Y|/�Er߱B��P�O��s�I��)s�T0 k� �4�8eA�s B1e 'Q  ��    ��� ��0EbC�"K��)���Y|/�Er�B��O�O��w�I��)s�T0 k� �4�8eA�s B1e 'Q  ��    ��� � 0Eb?�"K��)���Y|/�Er�B��O�O���I��)s�T0 k� �4�8eA�s B1e 'Q  ��    ��� �1Eb;�"K��)���Y|/�Er�B��O�K����I��)s�T0 k� �4�8eA�s B1e 'Q  ��    ��� �1D27�K��)���Y|/�Er�B��O�K����I��)s�T0 k� �4�8eA�s B1e 'Q  ��    ��� �2D23�K�Q�)���Y|/�Er�B��O�G����AR�)s�T0 k� �4 �8 eA�s B1e 'Q  ��    ��� �2D2+�K�Q�)��Y|/�Er�B��O�C����AR�)s�T0 k� �4 �8 eA�s B1e 'Q  ��   ��� ��3D2#�O�Q�)�{�Y|/�Eb��B��N�;�×�AR�)s�T0 k� �8!�<!eA�s B1e 'Q  ��    ��� ��4D2�O�Q�)�{�Y|/�Eb��B��N�7�Û�AR�)s�T0 k� �8!�<!eA�s B1e 'Q  ��    ��� �t4D2��S��)�w�Y|/�Eb��B��N�3�ß�AR�)s�T0 k� �8!�<!eA�s B1e 'Q  ��    ��� �t 4D2��S��)�w�Y|/�Ec�B��N�+�ã�A��)s�T0 k� �8!�<!eA�s B1e 'Q  ��    ��� �t$5D2��S��)�s�Y|/�Ec�B��N'�ã�A��3�T0 k� � "�$"eA�s B1e 'Q  ��    ��� �t$5D2��W��)�s�Y|/�D3�@b�N#�ç�A��3�T0 k� �#�#eA�s B1e 'Q  ��    ��� �t,6D1���[��)�k�Y|/�D3�@b�N�ë�A��3�T0 k� �$�$eA�s B1e 'Q  ��    ��� �t06DA���_��)�k�Y|/�D3�@b�N�ï�A��3�T0 k� ��$��$eA�s B1e 'Q  ��    ��� �t06DA���c��)�g�Y|/�D3�@b�N�ï�A��s� T0 k� ��#��#eA�s B1e 'Q  ��    ��� �d47DA���c��)�c�Y|/�D3�@��N�ðA��s� T0 k� ��"��"eA�s B1e 'Q  ��    ��� �d87DA���g��)�_�Y|/�D3�@��N��ðA��s� T0 k� ��"��"eA�s B1e 'Q  ��    ��� �d<7DA���o��)�[�Y|/�D3�@��N�ӴA��s�!T0 k� ��"��"eA�s B1e 'Q  ��    ��� �d<7EQ���s��|)�W�Y|/�D3�@��N�ӴA��s�!T0 k� ��#��#eA�s B1e 'Q  ��    ��� �d@7EQ���w��x)�S�Y|/�D3�A�N�ӴBB�s�!T0 k� ��#��#eA�s B1e 'Q  ��    ��� �d@7EQ���{��t)�O�Y|/�D3�A�N߷Ӵ	BB���"T0 k� ��"��"eA�s B1e 'Q  ��    ��� �T@7EQ������p)�K�Y|/�DC�A�N׷Ӵ
BB���"T0 k� ��!��!eA�s B1e 'Q  ��    ��� �TD7EQ�����d)�C�Y|/�DC�A�N˸ӴBB���"T0 k� ��!��!eA�s B1e 'Q  ��    ��� �TD7EQ�����`)�?�Y|/�DC�C��NøӰD����#T0 k� ��!��!eA�s B1e 'Q  ��    ��� �TD7EQ����\)�;�Y|/�DC�C��N��ӰD����#T0 k� ��!��!eA�s B1e 'Q  ��    ��� �TD7EQ����X)�7�Y|/�DC�C��N��ӰD����#T0 k� ��"��"eA�s B1e 'Q  ��    ��� �TD7EQ����P)�3�Y|/�DC�C��N��ӬD����#T0 k� ��"��"eA�s B1e 'Q  ��    ��� �TD6C����D)�'�Y|/�DC�C��Nћ��D����$T0 k� ��"��"eA�s B1e 'Q  ��    ��� ��@6C�|	³�@)�#�Y|/�DC�C��Nѓ��D����$T0 k� ��$��$eA�s B1e 'Q �    ��� ��@6C�x
»�8)��Y|/�DC�C��Nы��D��s�$T0 k� ��%��%eA�s B1e 'Q ��    ��� ��@6C�p�ê4)��Y|/�DS�C��Nу��D��s�%T0 k� �|'��'eA�s B1e 'Q ��    ��� ��<6C�`�ϫ$)��Y|/�DR��C��N�w��D��s�%T0 k� �d*�h*eA�s B1e 'Q ��    ��� ��86C�X׫ )��Y|/�DR��C��N�o��D��s�&T0 k� �X+�\+eA�s B1e 'Q ��    �   ��86C�P߫)��Y|/�DR��C�N�g��D��s�&T0 k� �L-�P-eA�s B1e 'Q ��    �  ��46C�L�)���Y|/�DR��C�N�_��D�#�s�'T0 k� �@.�D.eA�s B1e 'Q ��    �  ��06C�D�)���Y|/�DR��C�N�W��D�'���'T0 k� �40�80eA�s B1e 'Q ��    �  ��,6C�4���)���Y|/�DR��C�N�G��D�+���(T0 k� �3� 3eA�s B1e 'Q ��    �  ��(6I�,�	��)���Y|/�DR��C�N�?��D�/���(T0 k� �4�4eA�s B1e 'Q ��    �  ��$6I�$�	��)���Y|/�DR��C�N�7��Er3���)T0 k� �6�6eA�s B1e 'Q ��    �  �� 6I� �	��)���Y|/�Db��C�N�/��|Er3���)T0 k� ��8� 8eA�s B1e 'Q ��    �  ��6I��	��)���Y|/�Db��C�N�'��xEr7���*T0 k� ��9��9eA�s B1e 'Q ��    �  ��5I��/�	��)��Y|/�Db��C�N���tEr?���*T0 k� ��<��<eA�s B1e 'Q ��    � 	 |T5I��7�	��)�Y|/�Db��D�N���pEr?�s�+T0 k� ��>��>eA�s B1e 'Q ��    � 
 wT5I� �C�	��)�Y|/�Db��D�N���lErC�s�+T0 k� ��?��?eA�s B1e 'Q  ��    �  r                                                                                                                                                                            � � �  �  �  c A�  �J����  �      6 \���� ]�%d%d � 
�� dz.     	    � ��     dz. ��                   4		 Z           ��     ���   0			           Y��  * *	    � �_     YlC H=    P�              Z �         � �      ���   (
            Y�S     
	    Z�     Y�S Z�                     	 Z �        	     ���   8�          qP   � �
     ����     qP����                     9  Z            �  �  ���   (
	          OT.   � �	   . N�     Ou� &�    �`              S	 Z            �     ���   P
B          ��d �      B�r�    ��d�r�                             ���"              �  ���    8		 1              q��         V K�     q�� K��    �� V               	  3��                ��@   0	
           t��        j t     t�  q     � -               
   � �                ��@   0	          ��;   |	      ~���    ��;���8       S             S  ��          L�     ��J   8

          ���o   `       ��t    ���o�                         �         	  ��     ��@   0
          V�v  H	      � ��q     V� ���     :                   A �         
 P     ��@   8	
'           ���J ��     � ��]    ���J ��]                            ���u             ^  ��@    		 5                  ��      �                                                                           �                               ��        ���          ��                                                                 �                         �܂�  ��        ���"   ���܂����  ��   S                   x                j  �       �                         ��    ��        ���      ��  ��           "                                                 �                            �� � K �� � ������� 	  
              
   �   �A� ���J       �$ `c@ �� @d  �d  d� �� �e� �� f� �� 0f� �D  g@ �� g� ߤ \� ��  \� � 0Ȁ �� 0�  �H 0ǀ �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0� ���� ����� ����� � 
�< V� 
�� V� 
�\ W ���� � � �j� � k� �� 0o� �$ `p  �� p� � q  �$  q  � �t� �  u� �d 0r@ �� 0r� �$ s  �D  s  ��  s`  � �^@ � _@���� � <� p� <� p� <�  p� AD �[� BD  \� B� ]  ;� ``� <� a� <� a� <�  a� $ `t� � u�  u� 
�< W� 
�< W� 
�| W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����   %����  ������  
�fD
��L���"����D" � j  "  B   J jF�"    B�j l � 
����
��"     
�j,� B �
� �  �  
� ��    ��     ���       q��  ��     ���      ��    ��     ���          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �?      ��LT ��        � �T ��        �        ��        �        ��        �     ��    ��gl���        ��                         �$ (   �                                     �                ����            ���� ���%��   % �� F �            14/27 (51%) amnov y    5:30                                                                        3  3     �C
2�?C
� �;	CAKC C3C$C �J�+ J�; � J�; �	kjG 
kr7 �C.! � C61 �C71 �C:1 � C<$ �B�7 � B�? �C, � C4 �kVD � k^Dc"�<c "�NS"�<S*�K ~*8{ � *G{N  *P{ ~*8{ � *G{N  *P{N  *J{N  *P{ �"*P �  )�`N  *P{X  *P{ �&�- � 
�< � 
�@ � 
�B$**� �+"�9 � ,"�K �-�5 � 
�D r  "Q t ~  "K } u "V  2!� � � 3" � 4*@ �  *NX � 6*@ �  *NX �  *NX �  *Ne �:*4h �;"h � <"K p  ="B p(  "J p@  "F v                                                                                                                                                                                                                         p� P @       $   @ 
            ^ P E d  ���� M               �������������������������������������� ���������	�
��������                                                                                          ��    �N~�|� ��������������������������������������������������������   �4, :  * �� #� Q�� ���� � �=��                                                                                                                                                                                                                                                                                                                                @�                                                                                                                                                                                                                                             	          7 !   ��  L�J      M  	                           ������������������������������������������������������                                                                                                                                           �    ��                        ��                 	 	 ������� ����������������� ����������� ����������� ���� ������������������������������� � ����� ���������� �� ��� �� ������ � �������������   �������������� ������������� � ��������������� ����������� �� ���������������������                                   J             K
�J                                     ������������������������������������������������������                                                                      	                                                	                   �  �                  ��      ��              	 	 
  	 
 
 �������������� �   ����  �������������������������� ���������  ���������� ������� �����   � �� ����� ���������������� ����������� �������� ����  ���������� �������������������� �� ������������������������               x                                                                                                                                                                                                                                                          
                                                 �             


           �   }�         wwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwww , J >                                 � ��!Y �\                                                                                                                                                                                                                                                                                       YY	n  	�        m            m            l      m                                                                                                                                                                                                                                                                                                                                                                                                                     � <� �  � <��  �  ��  � (��  � 0��  � Z��  ���������������������o���������������������         <   t�E :! D          �   & AG� �  �              U��                                                                                                                                                                                                                                                                                                                                    p I F   �                       !��                                                                                                                                                                                                                            Y    �� �~ ��      �� 4      ������� ����������������� ����������� ����������� ���� ������������������������������� � ����� ���������� �� ��� �� ������ � �������������   �������������� ������������� � ��������������� ����������� �� ��������������������� �������������� �   ����  �������������������������� ���������  ���������� ������� �����   � �� ����� ���������������� ����������� �������� ����  ���������� �������������������� �� ������������������������        �     $�����������������������������������������������U���U���f��i����f��������U�ffU�ff|fff�vff�h�ffYff��������f�i�fffff��fffffffffffff������������f���fj��ff��ffi�lfk�ʪ���������������������������������������������������������������k�j�ff˖ff��ff��fffffffffff�ff��fff��fhvffgfffffffflf�ffffffffffff�f�f�f��|f�uUfffUffl�fffffffffff�fffk�fff��kf���f�fffffffffff��������ȩ��i���j���f���k���f������f���ƪ��f���f���f���f���f����fffffffffffff�fflfffffffffffƩfffffffff�k��f�fff�fk��k�Ʃ���Z���fffff�̼ffffʗW��UUUff�U�ɘUfl�Wfffl�fffff�f�̵vUx�Ux�̅x��U��XYf���j���l���f���ɩ������j���i������ƫ��ƚ�����������������������g�gVi�U�f��Z��evV��ƅ�U�e�U�fVVƋ��kkxWxh�uUȘuUȗ�Uȇ�u�x�����w�fgu��wuUww�UU�uUU�uUY�Uuy��Wy���f�Z�f�Vy�x�xWX�xUXUXuZ�XuY��U[�ɩ����������[���|���\���Y���U��������������������ʺ�������������fWVf�U��kU��i�v��jV�Y�Vx�e\��fUf�������W����ʇww˧��̹�w�j��Yl��ux��y�����XU����z���UX���x�h�UUy�U����������u�x��W��UY�uU{�Xu�����������U���w���X������������������ʛ��k�������ƪ��������ɪ�����yfeX�fku��liffh�flgff�e|���U�iXw��l��[f�Xu�f�x|�lu�l��W�u��Wuu�u�w�x��xwl����f�����gl��u�f�UUUUWx�YʌeV��U��e[��U���Z˛�����ʚ��������������������������������x����    B   &   .   � ��                       4     �  �����J����      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ��� ��� �    � �$ ^$    ��_�  �F  �   )   �   �    >�����������J������   p���� ��   p���� �$ ^h  ��     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h     `d ��     `d �$ ^$ �@       �      �     ��    `d �  `b���������� � �X�LX  ��L X         ��   "���� � ��� �� � ��� �$ ^$         �� 7 %      "       ���B��            �����  ��  yf  y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                           �            �  �� ��U�U]�U���U�� ��������UUUUU��������������������� ����UUU^U�����U]������������    �   ��  ^�  �^� UU���]����Վ                         �  �      �   �  �  �  ��  �U  �U  �U����U���]U��\�\�U��UU]�UUU]�UUU��������������]��]]��U]��UUUUUUUU�������������U�U��UU��U]]��U]�UU��U^��UU�����]]�U]�UU��U\�UU�UUU�   �   ^�  ^�  X�  U�  U�  U�    �U  �U  �U  �U  �  �   �   �UUU\UUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU]\�UUU��UU]�UUU\�UU]�UU��UX�U��U�UU��U\�UU��U��UU��UU��UUU݅U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUXU�  U�  U�  X�  Y�  ^�  �   �                                 �UUU�U^�� ��  ��  �        ���U�u�UU�UU��UUUUUU�UUU���� ���U^~�U^W�UU�UUU��UUUUUUU^������ UUU^�UU�~����� X�  ��          �                              wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                          t� O� ���O���O�������tG�O2$�""�3#"""4"23344w                                �   �   �   "   #   7   w   w   w   w                 wp C7 ttC4��O�����fw��fV~vefevff www  ��                        p   @   N   �p  v`  V`  g   w   p   @                 ww {�G J����� t�G ��Ow�K�w����{�K���{���{���t���wpw�0  w@      ~�  �  {�  {�  w�  K�  ��  �   �   w   w   w   w   �        t@	DD@G�@t��w�pwE�ptf^� fTG Vf  V  g  D                                       w�  v�  f`  g   w   w   w                ww wvU fe vf w }����}���}�� �� �� }�   �                p   p   f   @   �   p   p   �   @                              w  v  U   f  O  �� �� |� �~ }� �� ��  ��  ww  �@    p   g   Up  fp  �p  �~  ~� w� ��� ��� ��  ��  �w  ww   w         v  U  f   O������s��� ��� �� �� ��  ��  ww  �@    `   U   fp  �p  �p  �p�4p���}���}���� ��  �w  �w  ww   w       � ���w��w���y��p	�~� 	w �w�	�������H��D� wwp  C3  G     �  ��������	��p �~� 	w �w 	�� � p                           wp �w ��� ��# ��� ��� ~w� w�        p   p   p                 w� �  y�����	��	��wy����   �   �   �   w   w   �   w     w� �  y�����y��y��wy����   �   �   �   w   w   �   w   N _�^^gw�n�fvgvUgwffgwww ��        `   `   p   p                 w  �                     ��y �w������y���DD��p  ~@      	y��	t�	tI�ww  30  Dp   @          w  �   w                >�  .�  3p  wp  wp  wp  wp      w� �  w                        �   � ��� G�� �p  �p  wp  	p      ~� n� Vp Gp  p               wD �DD t�G��w�wt^�Feg    eW vfWpff`w�p��p~�w��p                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "  "!    " ""  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                              "! "   "      ""  !"""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �                      "  "!    " ""  !"!" "                ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  �   �   �   �   �       �     �"  "  �   "                                    �   �   �            �� �� �� g} �� vw                  � �� ��  ��    �     �                                                                                                                                                                                                          
   �   �  ��  �� ������-�� "��  �  
�  �C 
UU US �UD TE0 �� 
�� ʐ �  ̻  "�  "   " �� ����   �  �˰ ̻� �ݰ �w� ��� ����������˹�̹���ڙ��ٻ��ݰ̻� ˘  ��  3D  TD� 340 340 3D0 30 
��  ��  "/  "/  �� ���� �    ��                  "      �           �  �   �   ��  �            ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                      "  .���"    �     �                                                                                                                                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    ""  ""       @   H   H   D   D   L   �   �   �   ��� .���" ��"   /�  �  �              � ��         �� �� �� g} �� vw                     ��  ��  ���   ���� �                                                                                                                                                                                                            "  "(��ȩ�ܚ��ۊ����� ��  �   �   �   �   �� ��� ̻� ˽� ��� �w� �������������������������� �̻ ���         �   �       �   �   "" �+� Ȼ� ɫ� ɨ� ��                �� �I��3 ��D 
UD 
UD TD  T�  ˸  ��  �� ̰ �+ ��"/ �"/  ����  �D� 3E@ 4EJ 4ED ET DT �@ �� ��  �� ̰��+ "/ �"/���� ��  ��  �                            �   �    �   �       �   �   �                .          ܰ  ˻  ��  �w  ׶  vv        +  "  "     �  �                        �   ���                            �   �                                                                                                    w 
�� ɚ� ���
�˻Ɋ�����������-� �"+ ". "$ "$ �U  Z�  Z�  J�  J�  �D  ��  ��  ɘ ˰ "  �"/�"" "  �  �            g���z��ȩ�����ة�� ���  ̰  ̰  ˰  ��  �  N�� T4�CD  CD0 C40 C30 3;� ܰ �� �� �  �  "  �""�"" �"/���  � �  �      �     �   �   ��  �"" �""  ""   "                 �   ��   �                            � ����                 �  ��  �               �                                           � ��                  �  �˰ ��� �wp ���                                                                                                                                                                 UDD UU �D �;3 �ˈʙ�˫����""- ""+ �"����  �           J� �D�M�D���4���ˠ ��� ̽� ��� ��ٰ�۰"˰""+�""!��"�  �                        �� �ɪ�ܙ������ ��� ��� ��� ��� ��� H��        �� ��� ۻ� }݉ ��� ��� ��� �˼ ��� �ٚ��ک��М��J� "                           � � �  (�  .   .   )�  )�  �   �    �     �   �   �   �   �   �      �  �  �  �  �  �   �                                    �     �                                      � ����ݼ� ����                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����          �   �   �   �  �  �  �  �                                                                                                                                                                                                                 �  �� 	�� �� ̻  ̻  "+ "" "" �" �N  �D  �C �C �3 
�3 33 ���̈ ,� ""  """ ""�� ���                    � ��˰���Ъ�wp���й�vz˸w�������ܻ��ػ��������C;���;���;��"� "  "  
"� � , �"" """"" � ��� ����               �          �  �� ��� ��   �                    �   �   �             � ����  �                                 ��  ��  �          ���� ��� ����          �   �   �   �  �  �  �  �                          ����                               ���                          ����                  �   �� �       �  �  ��  �   �   �   �                                    �����̬̽��̽��̽���ת
wz� ��� ��� ˙� �) "+ .# 32� 33� �3> �3> �� � "  " "" "   "/� �  �                            �   ˰  ��  �̰ ��� �̻���ː�۹������̅�̙U�����
�ŀ���̵�̵K�D��"L�"  ""  "" ��.����������     �  ��  �   ��  ��            "   "   "   "   ��   ��  �  �   �    �               �   � � �  ��� ��  �                    �                        ���� ��� ����                            ��  ��  ���  �  �  �   �   ��  �                            �   ���                            �   �                                                                                                   �  ��� ��� }�� wݪ �� 	�� �� �ͼ ��� ��� ̘� �ͻ +���"�8"8  8� �� �U��EU��3 ̻�"̰""�" ��" �"                             �   ��� �˹��˚���ڍ�̽���ͽ��ͽ���ݼ��л�� ��D �UT EUT UU0 C3  2"  ""  -�  ��  ��  �   � ��"/ �" � ���    �        �   ��  ��  ��  ���        �                         ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ��� ���                                                   ����     �   �  �  �  ��  �   �                           ��   ��                  �  �  �� � ���    �  �                         ̰ �� ̻ {�����vz� w��  ��  ��  ̘  	�  
� "��,̻�"�� "#3  34  D  
�  �  " "" """ ! ��  ��                               ˹� �ɩ ��� �͋ ��� ��� ��̀��Ȑ���лܹнȝ0ݙ�@43�PCD�@@E�@ E�@ U�� H�  K�  �   ��    �� "�" ���                          �  �   ��  �  ��                �   �   �   "   "   "  !�    ��                              �                        ���� ��� ����                      �  �� ��  �    � ���                                                                                                                                                                                                 ̘����	�������͹���۸�����̌�+���(����ی��ی�N=��NC��U �� 	�� �� ��  ��  ��  ��  �� �� �� ��"� �    �            ��  ��  ̽� �݋ �ݨ�����)*������˚���ɛ���̽ݩ��ݚ���ɚ،̴X��E���E������������������������ ��� ��� �����������" � � �      �   �   �   �   �   �   �                   �   �   �   �   �   �   �   �   �  ��  �     ��     �   �  ��  ��  �   �            �   �   �   �    �                             �          �                        �         �  �� �  �� ��                                                                                                                                                   �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������  �  �  �   �   �            �   ��  ��  �  ɠ �  ��  ��        �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""������������������������""""�������DA�A�A""""�������H�H�DH�HH�""""������D""""������HADD���H""""��������D��""""�������H��H�H�H�""""�������A�D�HH�H""""������������������������"""$���4���4���4���4���4���4UUUUUUUUUUUUUUUUUU333DDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUEAUEQUUUTDDUUUU3333DDDDEQQQDUEUTDUUUU3333DDDDDDEUEUEUDTEUUUUU3333DDDDQDEQUUQUUQUUUDUUUUUU3333DDDDADAEQEQTEUDUUUU3333DDDDEUEUQUTDDUUUUU3333DDDDEUEQEEDUTDEUUUUU3333DDDDUUUUUUUUUUUUUUUUUUUUUUUU3333DDDDUUU4UUU4UUU4UUU4UUU4UUU43334DDDD"""������������������""""���������������������""""������II������""""������IIII""""������DI�I�""""������DI�I�""""�����IIDIIIA""""��������DD""""������IADD�A��""""��������I���I�������I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� = l � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����((�l(=����������������    � �aa � � � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����((�(( ���������������� x X � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����(-(5(Xx���������������� w w � �aa �	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	�� � ��ww����������������  � � �aa � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���� i���(���������������� �  � �aa � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � ��� u u��((����������������� ` m � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��m(`���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a��(M���������������� � � � �aa � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �a�� 
(����������������� � � u!a �  � � � �� � �� � � � � � �		 � � � �� � �� � � � � � ��� �)��(-(����������������� � � � � � � �  � � � � � �� � �� � �			 � � � �� � �� � � � ����(6(5���������������� u � � � � � � � � � � � �� � �� � � � � � � �		 � � �� � �� �� u u��(�x����������������  � �!!! � � � � � � � �� � ��"# �A�A�A�A�A�A� �	#	" � �� � �� �$% ���&&��ww����������������'( �))) �*++++,-.,-./0 �A�A�A�A�A�A� �	0	/,-.,-.+1++	*�&2���(+����������������34 �5 u u �*+++++6++6+/7 �A�A�A�A�A�A� �8/+6++6++1++*�&2��(W(�����������������9:  �AA � � � � � � � �� � ��"# �A�A�A�A�A�A� �#" � �� � �� �$% ���))�(a(����������������� U;'(AA � � � � � � � �� � �� � � � � � � � � � �� � �� �� u u��(����������������� =<34AA � � � � � ��� ��� � � �	 � ��� ��� � � � � ��� �A��l(=����������������    � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(( ���������������� x X � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �A��(Xx���������������� w w � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� �=�:	9ww����������������  � � �AA � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�>�; 
�(���������������� �  � �AA � � � � � � � � �� � � � � � � � � � � � � � � � � �� � � � � � ���	3?	<(+((����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+���������������� � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(����������������� � a � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����l(�(a(����������������� �  � �aa � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �����y(�(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqC
2�?C
� �;	CAKC C3C$C �J�+ J�; � J�; �	kjG 
kr7 �C.! � C61 �C71 �C:1 � C<$ �B�7 � B�? �C, � C4 �kVD � k^Dc"�<c "�NS"�<S*�K ~*8{ � *G{N  *P{ ~*8{ � *G{N  *P{N  *J{N  *P{ �"*P �  )�`N  *P{X  *P{ �&�- � 
�< � 
�@ � 
�B$**� �+"�9 � ,"�K �-�5 � 
�D r  "Q t ~  "K } u "V  2!� � � 3" � 4*@ �  *NX � 6*@ �  *NX �  *NX �  *Ne �:*4h �;"h � <"K p  ="B p(  "J p@  "F v3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������#�$��+�R�K�^�T�J�K�X��7�U�M�O�R�T�_� � � � �,�>�0�������������������������������������������.�G�R�K��2�G�]�K�X�I�N�[�Q� � � � � � �,�>�0�������������������������������������������+�R�K�^�K�O��C�N�G�S�T�U�\� � � � � � �@�9�1�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������@�9�1� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������,�>�0� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                