GST@�                                                           Zq     Z�                                               n	                        � h� 2���J���<a�����    ����        Ā      #    ����                                d8<n    �  ?    0�����  �
fD�
�L���"����D"� j   " B   J  jF�"     �j B  
���
��
�"    "�j��,  " ��
                                                                                  ����������������������������������      ��    a= Qb0 4 141 c  cc  cc  	     
     	   
        gG� �� 	(� (�                 -nn 21	         :8�����������������������������������������������������������������������������������������������������������������������������  bb    11                                                             �F  )          == �����������������������������������������������������������������������������                                �h  h   �  ��   @  #   �   �                                                                                'w w 2-1n	n  �)F    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E h �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    Er���.�H
!��|/�   $F@�4.�� � `�  T0 k� �C�#4� %�@2 ��A$0 � ��   �  Er��� .�P
!��|/�   (F@�4/�� � a�  T0 k� �C�#4� %�@2 ��A$0 � ��   �  Er����.�X
!��|/�   ,F@�8/�� � a�  T0 k� �C�#4� %�@2 ��A$0 � ��   �  Er����.�`
!��|/�   ,G@�</�� � b�  T0 k� �C�#D� %�@2 ��A$0 � ��   �  D����.�h
!��|/�   0G@�</�� � b�  T0 k� �C�#D� %�@2 ��A$0 � ��   �  D����.�p
!��|/�   4G@�@/�� � b�  T0 k� �C�#D� %�@2 ��A$0 � ��   �  D����.�|
���|/�   8G@�@/�� � c�  T0 k� �C�#D� %�@2 ��A$0 � ��   �  D����.��
���|/�   8H@�D0�� � c�  T0 k� �C�#D� %�@2 ��A$0 � ��   �  D����.��
���|/�   <H@�H0�� � c�
  T0 k� �C�#T� %�@2 ��A$0 � ��   �  D����.��
���|/�   @H@�H0�� � d�
  T0 k� �C�#T� %�@2 ��A$0 � ��   �  D�'���/��
���|/�   @I@�L0�� � d�
  T0 k� �C�#T� %�@2 ��A$0 � ��   �  D�+���/��
���|/�   DI@�L0�� � d,#�
  T0 k� �C�#T� %�@2 ��A$0 � ��   �  D�/�Ӵ/��
���|/�   HI@�P0�� � e,#�
  T0 k� �C�#T� %�@2 ��A$0 � ��   �  D�3�Ө/��
��|/�   HI@�T0�� � e,#�	  T0 k� �C�#t� %�@2 ��A$0 � ��   �  D�;�Ӡ/��
��|/�   LJ@�T1�� � e,#�	  T0 k� �C�#t� %�@2 ��A$0 � ��   �  D�?�Ӕ/��
��|/�   PJ@�T1�� � f,#�	  T0 k� �C�#t� %�@2 ��A$0 � ��   �  D�C�S�/����|/�   PJ@�P1�� � f,$ 	  T0 k� �C�#t� %�@2 ��A$0 � ��   �  D�G�S�/����|/�   TJ@�H1�� � f,4 	  T0 k� �C�#t� %�@2 ��A$0 � ��   �  D�K�S�/���#�|/�   XK@�D2�� � g,4   T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�O�S�/���+�|/�   XK@�@2�� � g,4  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�W�S�/���/�|/�   \K@�<2�� � g,4  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�[�S|.���7�|/�   \K@�83�� � g,4  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�_�Sx.� �;�|/�   `L@�43�� � h,4  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�g�Sp.��G�|/�   dL@�03�� � h,D  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�k�Sl.�K�|/�   hL@�,4�� �i,D  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�o�Sh.$�S�|/�   hL@�(4�� �i,D  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�s�Sd.,�W�|/�   lM@�$4�� �i,D  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�w�S`.4�_�|/�   lM@� 4�� �i,D  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�{�S\.<�c�|/�   pM@�5�� �j,D	  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D��SX.D�g�|/�   pM@�5�� �j,D	  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D���ST.L�o�|/�   tM@�5�� �j,D	  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D���SP-T�s�|/�   tN@�5�� �j,D	  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D���SL-\�w�|/�   xN@�6�� �k,D
  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D���SH-d�{�|/�   xN@�6�� �k,T
  T0 k� �C�#İ %�@2 ��A$0 � ��   �  D���SD-l�|/�   |N@�6�� �k,T
  T0 k� �C�#İ %�@2 ��A$0 � ��   �  D���SD-t�|/�   |N@�6�� �k,T
  T0 k� �C�#İ %�@2 ��A$0 � ��   �  D���S@-|�|/�   �O@� 7�� �l,T  T0 k� �C�#İ %�@2 ��A$0 � ��   �  D��S<-��|/�   �O@� 7�� �l,T  T0 k� �C�#İ %�@2 ��A$0 � ��   �  D��S8-��|/�   �O@��7�� �l,T  T0 k� �C�#԰ %�@2 ��A$0 � ��   �  E�����\m@�o��,  �,,B�4�L3�   T0 k� ��m��m%�@2 ��A$0 �  ��   � !��E�����^m8�o��,  �,,B�8�T3�   T0 k� ��n��n%�@2 ��A$0 �  ��   � "��E�����`m0�k��,  �(,B�<�\3�   T0 k� ��o��o%�@2 ��A$0 �  �� 
  � #��E����b},�k��,  �(-B�@#�`3�   T0 k� ��p��p%�@2 ��A$0 �  �� 
  � $��E����d}$�g��,  �$-B�D+�h3�   T0 k� ��r��r%�@2 ��A$0 �  �� 
  � %��E����f}�c��,  �$-B�H3�p3�   T0 k� ��t��t%�@2 ��A$0 �  �� 
  � &��E����i}�_��,  � -B�L;�x3�   T0 k� ��w��w%�@2 ��A$0 �  �� 
  � '��E����k}�_��,  �-B�TC��3�   T0 k� ��y��y%�@2 ��A$0 �  �� 
  � (��E����m��[��,	  �,B�XK��3�   T0 k� ��{��{%�@2 ��A$0 �  �� 
  � )��E����o��	}[��,	  �,B�\S��3�   T0 k� ��}��}%�@2 ��A$0 �  �� 
  � *��E����q�� 	}W��,	  �,E�`"[��3�   T0 k� ��{��{%�@2 ��A$0 �  �� 
  � +��E����s�� 	}S��,	  o,E�h "c��3�   T0 k� ��z��z%�@2 ��A$0 �  �� 
  � ,��E����u��!	}S��,
  o,E�l!"k��3�   T0 k� ��y��y%�@2 ��A$0 �  �� 
  � -��E����w��!	}S��,
  o+E�p""s��3�   T0 k� ��y��y%�@2 ��A$0 �  �� 
  � .��E����y��"	�O��,
  o+E�x""{��3�   T0 k� ��z��z%�@2 ��A$0 �  �� 
  � /��E�#���{��"	�O��,
  o+E�|#R�"�3�   T0 k� ��{��{%�@2 ��A$0 �  �� 	  � 0��E�#���}��#	�O��,
  _ +E��$R��"� 3�   T0 k� ��|��|%�@2 ��A$0 �  �� 	  � 1��E�#�����#	�K��,  ^�*E��%R��"�!3�   T0 k� ��}��}%�@2 ��A$0 �  �� 	  � 2��E�#������$	�K��,  ^�*E��&R��"�"3�   T0 k� ����%�@2 ��A$0 �  �� 	  � 3��E�#�޼���$	}K��,  ^�*E��'R��"�#3�   T0 k� ��~��~%�@2 ��A$0 �  �� 	  � 4��E�#���%	}K��,  ^�*E��(R��"�$3�   T0 k� ��y��y%�@2 ��A$0 �  �� 	  � 5��E�#����&	}K�",  ^�)E��)R��"�%"��   T0 k� ��t��t%�@2 ��A$0 �  �� 	  � 6��E�#����&	}K�",  N�)E��*R��"�&"��   T0 k� ��q��q%�@2 ��A$0 �  �� 	  � 7��E�#��~��'	}K�",  N�)E��+R��"�'"��   T0 k� ��n��n%�@2 ��A$0 �  �� 	  � 8��C�#��}��'	�K�",  N�)E�,B��"�("��   T0 k� ��l��l%�@2 ��A$0 �  �� 	  � 9��C�#���}��(	�K�",  N�)E�-B��"�)"��   T0 k� �|l��l%�@2 ��A$0 �  �� 	  � :��C����|��)	�K�",  N�)E�.B��*"��   T0 k� �tl�xl%�@2 ��A$0 �  �� 	  � ;��C����{��*	�K�",  N�)E�/B��+"��   T0 k� �ll�pl%�@2 ��A$0 �  �� 	  � <��C����{��+	�K�",  N�)E�0B��-"��   T0 k� �dk�hk%�@2 ��A$0 �  �� 	  � <��C����z��+	}K�",  N�)E�2���."��   T0 k� �`j�dj%�@2 ��A$0 �  �� 	  � <��C����y��,	}K�",  N�)E�3��� /"��   T0 k� �Xi�\i%�@2 ��A$0 �  �� 	  � <��C����xL�-	}K�",  N�)E�4���S$0"��   T0 k� �Ph�Th%�@2 ��A$0 �  �� 	  � <��C���|wL�.	}K��,  >�*E�6���S,13�   T0 k� �Lg�Pg%�@2 ��A$0 �  �� 	  � <��C���tvL�/	}K��,  >�*E�7���S023�   T0 k� �Dg�Hg%�@2 ��A$0 �  �� 	  � <��C���puL�/K��,  >�*E�8���S833�   T0 k� �@f�Df%�@2 ��A$0 �  �� 	  � <��C���htL�0K��,  >�+E�:���S<43�   T0 k� �8e�<e%�@2 ��A$0 �  �� 	  � <��C���dsL�0K��,  >�+E�;���S@53�   T0 k� �4d�8d%�@2 ��A$0 �  ��   � <��C���\rL�1K��,  >�+E�=���SH63�   T0 k� �,c�0c%�@2 ��A$0 �  ��   � <��C���XqL�1K��,  >�,Eo�>���SL73�   T0 k� �(b�,b%�@2 ��A$0 �  ��   � <��C����Pp\�2K��,  >�-E` @���SP83�   T0 k� � a�$a%�@2 ��A$0 �  ��   � <��C����Lo\�2K��,  >�-E`A���ST93�   T0 k� �_� _%�@2 ��A$0 �  ��   � <��C����Dn\�3K��,  >�.E`C����T:3�   T0 k� �^�^%�@2 ��A$0 �  ��   � <��C���@m\�3K��,  .�.E`D����X:3�   T0 k� �[�[%�@2 ��A$0 �  ��   � <��C���8l\�3 �K�!�,  .�/E`F����\;"s�   T0 k� �Y�Y%�@2 ��A$0 �  ��   � <��C���4k\�3 �K�!�,  .|0E`H����`<"s�   T0 k� �W�W%�@2 ��A$0 �  ��   � <��C���,j\�4 �K�!�,  .|1E`I����`="s�   T0 k� �U�U%�@2 ��A$0 �  ��   � <��C���$h\�4 �K�!�,  .x2E`K����d>"s�   T0 k� � R�R%�@2 ��A$0 �  ��   � <��D ߉� g\�4 �K�!�,  .t2E`L����d?"s�   T0 k� ��Q� Q%�@2 ��A$0 �  ��   � <��D ۉ�f\�4 �K�!�,  .p3E`N����h@"s�   T0 k� ��R��R%�@2 ��A$0 �  ��   � <��D Ӊ�e\�4 �K�!�,  .l4EP P����h@"s�   T0 k� ��R��R%�@2 ��A$0 �  ��   � <��D ω�cl�4 �K�!�,  .l5EP Q����hA"s�   T0 k� ��R��R%�@2 ��A$0 �  ��   � <��D ˉ�bl�4 �K�!�,  h6EP$S����lB"s�   T0 k� ��R��R%�@2 ��A$0 �  ��   � <��D Ê��al�4 �K�!�,  h7EP$T����lC"s�   T0 k� ��Q��Q%�@2 ��A$0 �  ��   � <��D ����_l�4 �K�!�,  d8EP$V����lC"s�   T0 k� ��P��P%�@2 ��A$0 �  ��   � <��D ����^l�4 �K��,  d8EP$W����lD3�   T0 k� ��O��O%�@2 ��A$0 �  ��   � <��D ����]L�4 �K��,  d9EP(Y����lE3�   T0 k� ��K��K%�@2 ��A$0 �  ��   � <��D ����[L�4 �K��,  `:EP(Z����lF3�   T0 k� ��H��H%�@2 ��A$0 �  ��   � <��D ����ZL�4 �K��,  `;EP(\����lF3�   T0 k� ��F��F%�@2 ��A$0 �  ��   � <��D����XL�4 �K��,  `<EP(]����lG3�   T0 k� ��C��C%�@2 ��A$0 �  ��   � <��D����WL�5 �K��,  `=E@(^���lH3�   T0 k� ��A��A%�@2 ��A$0 �  ��   � <��D����VL�5 �K��,  �`=E@(`���hH3�   T0 k� ��?��?%�@2 ��A$0 �  ��   � <��D����TL�5 �K��,  �`>E@(a���hI3�   T0 k� ��>��>%�@2 ��A$0 �  ��   � <��D����SL�6 �K��,  �`?E@(b���hJ3�   T0 k� ��<��<%�@2 ��A$0 �  ��   � <��D���QL�6 �K��,  �`@E@(c� �dJ3�   T0 k� ��;��;%�@2 ��A$0 �  ��   � <��D{���PL�6 �K��,  �`@E@(d� dK3�   T0 k� ��9��9%�@2 ��A$0 �  ��   � <��Ds���NL�7 �K��,  dAE@$e� dL3�   T0 k� ��8��8%�@2 ��A$0 �  ��   � <��Dk���LL�7 �K��,  dBE@$f�`L3�   T0 k� ��6��6%�@2 ��A$0 �  ��   � <��Dc���K,�8K��,  dBE@$g�\M3�   T0 k� ��4��4%�@2 ��A$0 �  ��   � <��E�_���I,�9K��,  hCE0$h�\N3�   T0 k� ��3��3%�@2 ��A$0 �  ��   � <��E�W���G,�9K��,  hDE0 i�XN3�   T0 k� ��1��1%�@2 ��A$0 �  ��   � <��E�O���F,�:K��,  �lDE0 i�TO3�   T0 k� ��/��/%�@2 ��A$0 �  ��   � <��E�G���D,�:K��,  �lEE0 j�TO3�   T0 k� ��.��.%�@2 ��A$0 �  ��   � <�E�?���B,�;K��,  �pFE0j�PP3�   T0 k� ��,��,%�@2 ��A$0 �  ��   � <�~E�7��xA�<]K��,  �pFE0k�LP3�   T0 k� ��*��*%�@2 ��A$0 �  ��   � <�}E�/�t?�<]K��,  �tFE k|HQ3�   T0 k� ��*��*%�@2 ��A$0 �  ��   � <�|E�'�p=�=]K��,  �tGE lxDQ3�   T0 k� ��)��)%�@2 ��A$0 �  ��   � <�{E��l;�>]K��,  ~xGE lp@R3�   T0 k� ��)��)%�@2 ��A$0 �  ��   � <�zE��h9�>]K��,  ~|GE ml<S3�   T0 k� ��(��(%�@2 ��A$0 �  ��   � <�yE��d8��?�K�|,  ~|HE mh8S3�   T0 k� ��'��'%�@2 ��A$0 �  ��   � <�xE��`6��?�K�|,  ~�HE m`4T3�   T0 k� ��%��%%�@2 ��A$0 �  ��   � <�wE���\4��@�K�|,  ~�HB�m\0T3�   T0 k� ��#��#%�@2 ��A$0 �  ��   � <�wE���X2��@�K�|,  ~�HB�m�T,U3�   T0 k� ��!��!%�@2 ��A$0 �  ��   � <�wE��T0��A�K�|,  ~�HB�n�P(U3�   T0 k� ����%�@2 ��A$0 �  ��   � <�wE��P.��A�K�|,  ~�HB�n�H V3�   T0 k� �|��%�@2 ��A$0 �  ��   � <�wE�ߐP,��B�K�|,  ��HB�n�@V3�   T0 k� �|��%�@2 ��A$0 �  ��   � <�wE�אL+��B�K�|,  ��GB�n�<V3�   T0 k� �x�|%�@2 ��A$0 �  ��   � <�wE�Ӑ�H)��B�K�|,  ��GB� n�4�W3�   T0 k� �p�t%�@2 ��A$0 �  ��   � <�wE�ˑ�H'��B�K�|,
  ��GB� n�,�W3�   T0 k� �l�p%�@2 ��A$0 �  ��   � <�wD?Ñ�D%��C�K�|,
  ��GB� n�(	�X3�   T0 k� �d�h%�@2 ��A$0 �  ��   � <�wD?���D#��C�K�|,
  ��FB� m� 	� X3�   T0 k� �`�d%�@2 ��A$0 �  ��   � <�wD?���D!��C�K�|,	  ��FB�$m�	��Y3�   T0 k� �`�d%�@2 ��A$0 �  ��   � <�wD?���@ ��C�K�|,	  ��EB�$m�
��Y3�   T0 k� �\�`%�@2 ��A$0 �  ��   � <�wD?���@��C�K�|,  ��EC (m�
��Y3�   T0 k� �\�`%�@2 ��A$0 �  ��   � <�wD?���@��C�K�|,  ��DC (m�
��Z3�   T0 k� �\�`%�@2 ��A$0 �  ��   � <�wD?���@ �C�K�|,  ��CC ,l��
��Z3�   T0 k� �\�`%�@2 ��A$0 �  ��   � <�wD?���@ �C�K�|,  ��CC ,l����[3�   T0 k� �\�`%�@2 ��A$0 �  ��   � <�xD?�� -@ �C�K�|,  ��BC 0l����[3�   T0 k� �l�p%�@2 ��A$0 �  ��   � <�yD?{� -@ �C�K�|,  ��AC 0k����[3�   T0 k� �x�|%�@2 ��A$0 �  ��   � <�zD?s� -@ �C�K�|,  ��@C 4k����\3�   T0 k� ����%�@2 ��A$0 �  ��   � <�{D?o� -D �C�K�|,  ��@C 4j����\3�   T0 k� ����%�@2 ��A$0 �  ��   � ;�|DOg� -D �C�K�|,  ��?C 8j���]3�   T0 k� ����%�@2 ��A$0 �  ��   � :�}DO_� -D �C�K�|,  ~�>C <i���]3�   T0 k� ����%�@2 ��A$0 �  ��   � 9�~DOW� -H �C�K�|,  ~�=C @i��]3�   T0 k� ����%�@2 ��A$0 �  ��   � 8�DOO� -HL�CmK�|,  ~�<C@h��^3�   T0 k� ����%�@2 ��A$0 �  ��   � 7��DOG� -LL�CmK�|,  ~�;CDg��^3�   T0 k� ��	��	%�@2 ��A$0 �  ��   � 6��E�?� -L
L�CmK�|,  ~�:CHg��^3�   T0 k� ����%�@2 ��A$0 �  ��   � 5��E�;� -P	L�CmK�|,  n�9CLf��_3�   T0 k� ����%�@2 ��A$0 �  ��   � 4��E�3� -PL�CmG�|,  n�7CLf��_3�   T0 k� ����%�@2 ��A$0 �  ��   � 3��E�+� =TL�CmG�|,  n�6CPe��_3�   T0 k� ����%�@2 ��A$0 �  �� 	  � 2��E�#� =XL�CmG�|,  n�5CTd�x`3�   T0 k� ����%�@2 ��A$0 �  �� 	  � 1��E�� =\L�CmG�|,  n�4CXcxp`3�   T0 k� ����%�@2 ��A$0 �  �� 	  � 0��E�� =`L�CmC�|,  >�3C\bph`3�   T0 k� �� �� %�@2 ��A$0 �  �� 	  � /��E�� =`L�CmC�|,  >�2C`bh`a3�   T0 k� ������%�@2 ��A$0 �  �� 	  � .��E�� =d L�C=C�|,  >�0Cda`Xa3�   T0 k� ������%�@2 ��A$0 �  �� 	  � -��E��� =k�L�C=?�|,  >�/C h`XPa3�   T0 k� ������%�@2 ��A$0 �  �� 	  � ,��E��� =o�L�C=?�|,  >�.C l_P�Ha3�   T0 k� ������%�@2 ��A$0 �  �� 	  � +��E�� =s�L�C=;�|,  >�,C p^H�@b3�   T0 k� ������%�@2 ��A$0 �  �� 	  � *��E�� =w�L�C=;�|,  >�+C t]@�8b3�   T0 k� ������%�@2 ��A$0 �  �� 	  � )��E�� =�L�Cm7�|,  n�*C x\4�0b3�   T0 k� ������%�@2 ��A$0 �  �� 	  � (��E�ߦ M����Cm7�|,  n�(C |[,�(b3�   T0 k� ������%�@2 ��A$0 �  �� 	  � '��E�ק M����Cm3�|,  n�'C �Z$� b3�   T0 k� ������%�@2 ��A$0 �  �� 	  � &��E�Ϩ M����Cm/�|,  n�&C �Y�b3�   T0 k� ������%�@2 ��A$0 �  �� 	  � %��E�˩ M����Cm/�|,  n�$C �X	��b3�   T0 k� ������%�@2 ��A$0 �  �� 	  � $��E�ê M����Bm+�|,  n�#C �W	��b3�   T0 k� ������%�@2 ��A$0 �  �� 	  � #��E��� M����B]'�|,  n�!C �V	�� b3�   T0 k� �����%�@2 ��A$0 �  �� 	  � "��E��� M����B]#�|,  n� B�U	����b3�   T0 k� ����%�@2 ��A$0 �  �� 	  � !��F�� M����B]#�|,  n�B�T	����b3�   T0 k� ����%�@2 ��A$0 �  �� 	  �  ��F�� M����A]�|,  ^�B�S	����a3�   T0 k� ����%�@2 ��A$0 �  �� 	  � ��F�� M����A]�|,  ^�B�R	����a3�   T0 k� ����%�@2 ��A$0 �  �� 	  � ��F�� M����@m�|,  ^�B�P	����a3�   T0 k� ����%�@2 ��A$0 �  �� 	  � ��F�� ]����@m�|,  ^�B�O	����a3�   T0 k� �#��'�%�@2 ��A$0 �  �� 	  � ��F�� ]����?m�|,  ^�B�N	����`3�   T0 k� �+��/�%�@2 ��A$0 �  �� 	  � ��F�� ]����?m�|,  �B�M	����`3�   T0 k� �/��3�%�@2 ��A$0 �  �� 	  � ��F�� ]����>m�|,  �B��K	���_3�   T0 k� �7��;�%�@2 ��A$0 �  �� 
  � ��F�� ]����>}�|,  �B��J	���_3�   T0 k� �?��C�%�@2 ��A$0 �  �� 
  � ��F�������=}�|,   �B��I	���^3�   T0 k� �/��3�%�@2 ��A$0 �  �� 
  � ��F�������<}�|,   �B��H	���]3�   T0 k� �'��+�%�@2 ��A$0 �  �� 
  � ��F�������;}�|,   �C �F	���]3�   T0 k� �#��'�%�@2 ��A$0 �  �� 
  � ��E�������;}�|,   �C �Eд�\3�   T0 k� �#��'�%�@2 ��A$0 �  �� 
  � ��E�������:���|/�  �C �DЬ�[3�   T0 k� �#��'�%�@2 ��A$0 �  �� 
  � ��E�{�����9���|/�  �|	C �BШ�[3�   T0 k� �'��+�%�@2 ��A$0 �  �� 
  � ��E�w�^���8���|/�  �|C �AФ�Z3�   T0 k� �+��/�%�@2 ��A$0 �  �� 
  � ��E�w�^���7���|/�  �xC �?М�Y3�   T0 k� �/��3�%�@2 ��A$0 �  �� 
  � ��E�s�^���6���|/�  �tC �>И�X3�   T0 k� �3��7�%�@2 ��A$0 �  �� 
  � ��E�s�^���5���|/�  �pC=АxW3�   T0 k� �;��?�%�@2 ��A$0 �  �� 
  � ��E�s�^'���4��|/�  �lC;���tW3�   T0 k� �C��G�%�@2 ��A$0 �  �� 
  � ��E�s�^/���3��|/�  ~k�C:���pV3�   T0 k� �K��O�%�@2 ��A$0 �  ��   � ��E�o�^7���2��|/�  ~k�E�9���lU3�   T0 k� �S��W�%�@2 ��A$0 �  ��   � ��E�o�^?���1��|/�  ~g�E�7�x�hT3�   T0 k� �[��_�%�@2 ��A$0 �  ��   � 
��E�o�^?���0��|/�  ~c�E� 6�t�dS3�   T0 k� �[��_�%�@2 ��A$0 �  ��   � 	��E�s�^C���.
��|/�  ~_�E�$4�l�`R3�   T0 k� �_��c�%�@2 ��A$0 �  ��   � ��E�w��G���-
��|/�  ~_�E�,3�d`Q3�   T0 k� �c��g�%�@2 ��A$0 �  ��   � ��E�{��G���,
��|/�  ~[�E�01�`\P3�   T0 k� �c��g�%�@2 ��A$0 �  ��   � ��E��K���+
��|/�  ~[�E�40�XXO3�   T0 k� �g��k�%�@2 ��A$0 �  �   � ��E���O���)
��|/�  ~[�E�8.�TXN3�   T0 k� �g��k�%�@2 ��A$0 �  ��   � ��E���O���(
��|/�  ~[�E�@-�LTM3�   T0 k� �k��o�%�@2 ��A$0 �  ��   � ��E���O���'
��|/�  ~W�E�D+�DPK3�   T0 k� �k��o�%�@2 ��A$0 �  ��   � ��E���O���%
��|/�  ~W�CAH)�@PJ3�   T0 k� �k��o�%�@2 ��A$0 �  ��   � ��E���S���$
��|/�  ~W�CAL(�8LI3�   T0 k� �o��s�%�@2 ��A$0 �  ��   �  ��E���S���#
��|/�  ~S�CAT&�4LH3�   T0 k� �o��s�%�@2 ��A$0 �  ��   �����E����W���!
,��|/�  ~S�CAX%�,�LG3�   T0 k� �s��w�%�@2 ��A$0 �  ��   �����E����[��� 
,��|/�  ~S�CA\#�(�HF3�   T0 k� �w��{�%�@2 ��A$0 �  ��   �����E����_���
,��|/�  ~S�CA`!� �HE3�   T0 k� �{���%�@2 ��A$0 �  ��   �����E����_�	ܠ
,��|/�  ~O�CAd �
�HC3�   T0 k� �{���%�@2 ��A$0 �  ��   �����E��� ~c�	ܠ
,��|/�  ~O�CAh�	�HB3�   T0 k� �����%�@2 ��A$0 �  ��   �����E��� ~g�	ܠ
,��|/�  ~O�CAp�	�HA3�   T0 k� ������%�@2 ��A$0 �  ��   �����E��� ~k�	ܠ
,��|/�  ~O�CAt��H@3�   T0 k� ������%�@2 ��A$0 �  ��   �����E��� ~o�	ܠ
,��|/�  ~K�CAx �H?3�   T0 k� ������%�@2 ��A$0 �  ��   �����E��� ~s�	ܠ
,��|/�  ~K�CA|  �H>3�   T0 k� ������%�@2 ��A$0 �  ��   �����E��� ~w�	�
,��|/�  ~K�CQ���H=3�   T0 k� ������%�@2 ��A$0 �  ��   �����E��� ~{�	�
,��|/�  ~K�CQ���H<3�   T0 k� ������%�@2 ��A$0 �  ��   �����E��� ~�	�
��|/�  ~G�CQ���L;3�   T0 k� ������%�@2 ��A$0 �  ��   �����E��� ~��	�
��|/�  ~G�CQ���L:3�   T0 k� ������%�@2 ��A$0 �  ��   �����E��� ���	�
��|/�  ~G�CQ���L93�   T0 k� ������%�@2 ��A$0 �  ��   �����E��� ���	ܠ
��|/�  ~G�IQ�� �P83�   T0 k� ������%�@2 ��A$0 �  ��   �����E��� ���	ܠ
��|/�  ~G�IQ����P83�   T0 k� ������%�@2 ��A$0 �  ��   �����E�� ���	ܠ
��|/�  ~C�IQ����T73�   T0 k� ������%�@2 ��A$0 �  ��   �����E�� ���	ܠ
��|/�  ~C�IQ�	���T63�   T0 k� ������%�@2 ��A$0 �  ��   �����E�� ���	ܠ
��|/�  ~C�IQ����!T53�   T0 k� ������%�@2 ��A$0 �  ��   �����E�� ���	�
��|/�  ~C�Ia����!X43�   T0 k� ������%�@2 ��A$0 �  ��   �����E���	�
��|/�  �C�Ia����!X33�   T0 k� ������%�@2 ��A$0 �  ��   �����E'���	�
��|/�  �?�Ia����!\23�   T0 k� ������%�@2 ��A$0 �  ��   �����E/���	�
��|/�  �?�Ia����!\13�   T0 k� ������%�@2 ��A$0 �  ��   �����E7���	�
��|/�  �?�Ia����!\03�   T0 k� ������%�@2 ��A$0 �  ��   �����E?���	ܠ
��|/�  �?�IQ����!\/3�   T0 k� ������%�@2 ��A$0 �  ��   �����EG����	ܠ
��|/�  ?�IQ� ���1\.3�   T0 k� ������%�@2 ��A$0 �  ��   �����B�O����	ܠ

��|/�  ?�IQ�����1`-3�   T0 k� ������%�@2 ��A$0 �  ��   �����B�W����	ܠ

��|/�  ?�IQ�����1`,3�   T0 k� ������%�@2 ��A$0 �  ��   �����B�_����	ܠ

��|/�  ;�IQ�����1`*3�   T0 k� ������%�@2 ��A$0 �  ��   �����B�g����	�

��|/�  ?�Ia�����1`)3�   T0 k� ������%�@2 ��A$0 �  ��   �����B�o����	�

��|/�  ?�Ia�����1`(3�   T0 k� ������%�@2 ��A$0 �  ��   �����B�w����	�

��|/�  ?�Ia�����1`'3�   T0 k� ������%�@2 ��A$0 �  ��   �����B�����	�

��|/�  ?�Ia�����1d%3�   T0 k� ����%�@2 ��A$0 �  ��   �����B������	�

��|/�  ?�Ia�����1d$3�   T0 k� ����%�@2 ��A$0 �  ��   �����B��������

��|/�  �?�CA�����1d"3�   T0 k� ����%�@2 ��A$0 �  ��   �����B��������

��|/�  �?�CA�����Ad!3�   T0 k� ����%�@2 ��A$0 �  ��   �����B��������

��|/�  �C�CA�����Ad 3�   T0 k� ����%�@2 ��A$0 �  ��   �����B�������

��|/�  �C�CA�����Ah3�   T0 k� ����%�@2 ��A$0 �  ��   �����B�������

��|/�  �G�CA�����Ah3�   T0 k� ����%�@2 ��A$0 �  ��   �����B�����L�
���|/�  �G�E������Ah3�   T0 k� ����%�@2 ��A$0 �  ��   �����B�����L�
���|/�  �K�E������Al3�   T0 k� ����%�@2 ��A$0 �  ��   �����B�����L�
���|/�  �K�E������Al3�   T0 k� ����%�@2 ��A$0 �  ��   �����B��� �#�L�
���|/�  �O�E������Al3�   T0 k� ����%�@2 ��A$0 �  ��   �����E��� �'�L�
���|/�  �S�E������Ap3�   T0 k� ����%�@2 ��A$0 �  ��   �����E��� �/� �
���|/�  �S�E������Ap3�   T0 k� ���#�%�@2 ��A$0 �  ��   ���  E��� �3� �
���|/�  �W�E������Qt3�   T0 k� �'��+�%�@2 ��A$0 �  ��   ��� E��� �7� �
���|/�  �[�E������Qt3�   T0 k� �+��/�%�@2 ��A$0 �  ��   ��� E��� �?� �
���|/�  �[�E������Qx3�   T0 k� �3��7�%�@2 ��A$0 �  ��   ��� E��� �C� �
���|/�  �_�E������Q|3�   T0 k� �7��;�%�@2 ��A$0 �  ��   ��� E��/G���
���|/�  �c�E������Q|3�   T0 k� �C��G�%�@2 ��A$0 �  ��   ��� B��/O���
���|/�  �g�E������
р3�   T0 k� �K��O�%�@2 ��A$0 �  ��   ��� B��/S���
���|/�  �k�E������
ф	3�   T0 k� �W��[�%�@2 ��A$0 �  ��   ��� B��/W���
���|/�  �o�E������
ш3�   T0 k� �_��c�%�@2 ��A$0 �  ��   ��� B�#�/_���
���|/�  �s�E������
ь3�   T0 k� �g��k�%�@2 ��A$0 �  ��   ��� 	B�+�/c���
���|/�  �w�E�����
ѐ3�   T0 k� �k��o�%�@2 ��A$0 �  ��   ��� E�3�/g���
���|/�  �{�E���
@�Q�3�   T0 k� �o��s�%�@2 ��A$0 �  ��   ��� E�;�/o���
���|/�  ��E���
@�Q�3�   T0 k� �w��{�%�@2 ��A$0 �  ��   ��� E�C�/s���
���|/�  ���E���
@�Q�3�   T0 k� �{���%�@2 ��A$0 �  ��   ��� E�K�/w���
���|/�  ���E���
@�Q�3�   T0 k� �����%�@2 ��A$0 �  ��   ��� E�S�/���
���|/�  ���E���
@�Q� 3�   T0 k� ������%�@2 ��A$0 �  ��   ��� E�W�/����
���|/�  ���E��� �Q��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� E�_�/����
���|/�  ���Eѿ� �Q��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� E�g�/����
���|/�  ��Eѿ� #�Q��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� E�o�/����
���|/�  ��Eѻ� '�Q��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� E�w�/����
���|/�  ��Eѻ� '�Q��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� E��/����
���|/�  ��Eѷ�0+�Q��3�   T0 k� ������%�@2 ��A$0 �  ��   ���  C@��/����
���|/�  ��E᷿0/�A��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� "C@��/����
���|/�  ��E᳾0/�A��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� $C@��/����
��|/�  ��E᯽03�A��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� &C@��/����
��|/�  ��E᯻07�A��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� (C@��/����
��|/�  ��E᫺07�A��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� *C@������
��|/�  ǩE᧹@;�A��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� ,C@������
��|/�  �ϪE᣸@;�1��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� .C@������
�#�|/�  �׬E៷@7�1��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� 0CP������
�'�|/�  ��E៶@7�1��3�   T0 k� ������%�@2 ��A$0 �  ��   ��� 2CP������
�+�!�/�  ��Eᛵ@3�1��"s�   T0 k� ������%�@2 ��A$0 �  ��   ��� 4CP������
�3�!�/�  ��Eᗴ�3�1��"s�   T0 k� ������%�@2 ��A$0 �  ��   ��� 6CP������
�7�!�/�  ���E��/�A��"s�   T0 k� ������%�@2 ��A$0 �  ��   ��� 8CPϿ��� 
�;�!�/�  ��E��/�A��"s�   T0 k� ����%�@2 ��A$0 �  ��   ��� :CPӽ���
�C�!�/�  ��E��/�A��"s�   T0 k� ����%�@2 ��A$0 �  ��   ��� <CPۼ��
�G�!�/�  ��E��+�A��"s�   T0 k� ����%�@2 ��A$0 �  ��   ��� >CP߻��
�K�!�/�  �#�E��+�A��"s�   T0 k� ����%�@2 ��A$0 �  ��   ��� @CP�� �
�O�!�/�  �+�E��'� a��"s�   T0 k� �#��'�%�@2 ��A$0 �  ��   ��� BCP���
�W�!�/�  �3�E���'� a��"s�   T0 k� �+��/�%�@2 ��A$0 �  ��   ��� DCP�� �
�[�!�/�  �;�E�{��'� a��"s�   T0 k� �3��7�%�@2 ��A$0 �  ��   ��� FC`��(�
�_�!�/�  �C�D�w��#� a��"s�   T0 k� �;��?�%�@2 ��A$0 �  ��   ��� HC`���0�
�c�|/�  �K�D�w��#� a��3�   T0 k� �C��G�%�@2 ��A$0 �  ��   ��� JC`���8� 
�g�|/�  �S�D�s��#���3�   T0 k� �K��O�%�@2 ��A$0 �  ��   ��� LCa��<�$
�k�|/�  �[�D�o�����3�   T0 k� �S��W�%�@2 ��A$0 �  ��   ��� NCa��D�(
�o�|/�  �_�D�k�����3�   T0 k� �X �\ %�@2 ��A$0 �  ��   ��� PE���L
�,
�w�|/�  �g�D�k�����3�   T0 k� �`�d%�@2 ��A$0 �  ��   ��� RE���T�0
�{�|/�  �o�D�g�����3�   T0 k� �h�l%�@2 ��A$0 �  ��   ��� TE���\�4
��|/�  �w�D�c���1��3�   T0 k� �p�t%�@2 ��A$0 �  ��   ��� VE���d�4
݃�|/�  ��D�c���1��3�   T0 k� �x
�|
%�@2 ��A$0 �  ��   ��� XE���l�8
݇�|/�  ��D�_���1��3�   T0 k� ����%�@2 ��A$0 �  ��   ��� ZE�#��t�<
݋�|/�  ��D�[���1��3�   T0 k� ����%�@2 ��A$0 �  ��   ��� \E�'��|�@
ݏ�|/�  ��D�[���1��3�   T0 k� ����%�@2 ��A$0 �  ��   ��� ^E�+����D
ݓ�!�/�  ��D�W���A��"��   T0 k� ����%�@2 ��A$0 �  ��   ��� `E�/����D
ݗ�!�/�  ���D�S�@�A��"��   T0 k� ����%�@2 ��A$0 �  ��   ��� bE�3����H
ݛ�!�/�  ���D�S�@�A��"��   T0 k� ����%�@2 ��A$0 �  ��   ��� dE�7����L
ݛ�!�/�  ���D�O�@�A��"��  T0 k� �� �� %�@2 ��A$0 �  ��   ��� fE�;����P
ݟ�!�/�  ���D�K�@�A��"��  T0 k� ��!��!%�@2 ��A$0 �  ��   ��� hE�?� ��P
ݣ�!�/�  ���D�K�@�Q��"��  T0 k� ��"��"%�@2 ��A$0 �  ��   ��� jE�C� ��T
ݧ�!�/�  ���D�G�0�Q��"��  T0 k� ��#��#%�@2 ��A$0 �  ��   ��� lE�C� ��X
ݫ�!�/�  ���D�G�0�Q��"��  T0 k� ��$��$%�@2 ��A$0 �  ��   ��� nE�G� ��X
ݯ�!�/�  ���D�C�0�Q��"��  T0 k� ��%��%%�@2 ��A$0 �  ��   ��� pE�K� ��\
ݳ�!�/�  ���D�C�0�Q��"��  T0 k� ��&��&%�@2 ��A$0 �  ��   ��� rE�K���`
ݷ�!�/�  ���D�?�0�a��"��  T0 k� ��"��"%�@2 ��A$0 �  ��   ��� tE�O���`
ݷ�|/�  ���D�?� �a��3�  T0 k� ����%�@2 ��A$0 �  ��   ��� vE�O���d
ݻ�|/�  ���D�;� �a��3�  T0 k� ����%�@2 ��A$0 �  ��   ��� xE�O���h
ݿ�|/�  ���D�7� �a��3�  T0 k� ��� %�@2 ��A$0 �  ��   ��� zE�S���h
���|/�  ���D�7� �a��3�  T0 k� ��%�@2 ��A$0 �  ��   ��� |E�S�� �l
���|/�  ��D�3� #�a��3�  T0 k� ��%�@2 ��A$0 �  ��   ��� ~E�S� !�l
���|/�  ��D�3� '�a��3�  T0 k� ��%�@2 ��A$0 �  ��   ��� �E�S�"�p
���|/�  ��D�/�'�a��3�  T0 k� �� %�@2 ��A$0 �  ��   ��� �E�S��#�t
���|/�  ��D�/�+�a��3�  T0 k� �$�(%�@2 ��A$0 �  ��   ��� �E�S��#�t
���|/�  ��D�/�/���3�  T0 k� �,�0%�@2 ��A$0 �  ��   ��� �E�S� $�x
���|/�  ��D�+�3���3�  T0 k� �4�8%�@2 ��A$0 �  ��   ��� �E�S��(%�x
���|/�  �#�D�+�7���3�  T0 k� �<�@%�@2 ��A$0 �  ��   ��� �E�S��0%�|
���|/�  �'�Ea'��;���3�  T0 k� �D�H%�@2 ��A$0 �  ��   ��� �E�S��8&�|
���|/�  �/�Ea'��?��3�  T0 k� �L�P%�@2 ��A$0 �  ��   ��� �E�S��@'݀
���|/�  �3�Ea#��G��3�  T0 k� �X�\%�@2 ��A$0 �  ��   ��� �E�S��H'݀
���|/�  �7�Ea��K��3�  T0 k� �`�d%�@2 ��A$0 �  ��   ��� �E�O��P(݄
���|/�  �;�Ea��O��3�  T0 k� �h"�l"%�@2 ��A$0 �  ��   �   �E�O��X(݄
���|/�  �?�Ea��S��3�  T0 k� �p#�t#%�@2 ��A$0 �  ��   �   �EQO��`)݈
���|/�  �C�Ea��W��3�  T0 k� �x%�|%%�@2 ��A$0 �  ��   �  �EQK��l*݈
���|/�  �K�Ea��_��3�  T0 k� ��'��'%�@2 ��A$0 �  ��   �  �EQK��t*��
���|/�  O�Ea��`#�3�  T0 k� ��(��(%�@2 ��A$0 �  ��   �  �EQG��|+��
���|/�  W�Ea��d+�3�  T0 k� ��)��)%�@2 ��A$0 �  ��   �  �EQG���+��
���|/�  c�D1��l/�3�  T0 k� ��)��)%�@2 ��A$0 �  ��   �  �EQC���,��
���|/�  o�D1��p3�3�  T0 k� ��*��*%�@2 ��A$0 �  ��   �  �EQ?���,��
���|/�  w�D1��x7�3�  T0 k� ��*��*%�@2 ��A$0 �  ��   �  �EQ?���-��
���|/�  ���D1��|?�3�  T0 k� ��+��+%�@2 ��A$0 �  ��   �  �EQ;���-��
���|/�  ���D1���C�3�  T0 k� ��+��+%�@2 ��A$0 �  ��   �  �C�7���.��
��|/�  ���E�����	G�3�  T0 k� ��,��,%�@2 ��A$0 �  ��   �  �C�3���.��
��|/�  ���E�����
O�3�  T0 k� ��,��,%�@2 ��A$0 �  ��   �  �C�3���/��
��|/�  ���E�����S�3�  T0 k� ��-��-%�@2 ��A$0 �  ��   �  �C�/���/��
��|/�  ���E�����[�3�  T0 k� ��-��-%�@2 ��A$0 �  ��   �  �C�+���0��
��|/�  ���E�����_�3�  T0 k� ��.��.%�@2 ��A$0 �  �� 
  �  �C�+���0��
��|/�  ���E�����c�3�  T0 k� ��.��.%�@2 ��A$0 �  �� 
  �  �C�'��1��
��|/�  ���E�����h 3�  T0 k� ��.��.%�@2 ��A$0 �  �� 
  � 	 �C�'��1��
�#�|/�  ���F ����l3�  T0 k� ��-� -%�@2 ��A$0 �  �� 
  � 	 �C�#��1��
�'�|/�  ���F ����t3�  T0 k� �-�-%�@2 ��A$0 �  �� 
  � 	 �C�#��2��
�+�|/�  ���F���x3�  T0 k� �,�,%�@2 ��A$0 �  �� 
  � 
 �C��2��
�/�|/�  ���F����3�  T0 k� �,�,%�@2 ��A$0 �  �� 
  � 
 �C��3��
�7�|/�  ���F����3�  T0 k� �,� ,%�@2 ��A$0 �  �� 
  �  �C��3��
�;�|/�  ���F����3�  T0 k� �$,�(,%�@2 ��A$0 �  �� 
  �  �C��4��
�C�|/�  ���F����3�  T0 k� �0-�4-%�@2 ��A$0 �  �� 
  �  �C��$4��
�G�|/�  ���F����3�  T0 k� �8-�<-%�@2 ��A$0 �  �� 
  �  �C��04��
�K�|/�  ���F����	3�  T0 k� �@.�D.%�@2 ��A$0 �  �� 
  �  �C���85��
�S�|/�  ���F���R�
3�  T0 k� �H*�L*%�@2 ��A$0 �  �� 
  �  �C���@5��
�W�|/�  ���D��� R�3�  T0 k� �P'�T'%�@2 ��A$0 �  �� 	  �  �C���H5��
�_�|/�  ���D���R�3�  T0 k� �\%�`%%�@2 ��A$0 �  �� 	  �  �C���P5��
�g�|/�  ���D�#��R�3�  T0 k� �d$�h$%�@2 ��A$0 �  �� 	  �  �C���\6��
�k�|/�  ���D�'��R�3�  T0 k� �l#�p#%�@2 ��A$0 �  �� 	  �  �A���d6� 
�s�|/�  ���D�+�� R�3�  T0 k� �t"�x"%�@2 ��A$0 �  �� 	  �  �A���l6�
�w�|/�  ���D�/��(R�3�  T0 k� ��!��!%�@2 ��A$0 �  �� 	  �  �A���t6�
��|/�  ���D�3��0R�3�  T0 k� �� �� %�@2 ��A$0 �  �� 	  �  �A���|6�
·�|/�  ��D�7��8 R�3�  T0 k� �� �� %�@2 ��A$0 �  �� 	  �  �A����6�
Ώ�|/�  ��D�;��@ R�3�  T0 k� �� �� %�@2 ��A$0 �  �� 	  �  �A��R�6�
Γ�|/�  ��D�?��H!��3�  T0 k� ��!��!%�@2 ��A$0 �  �� 	  �  �A��R�6�$
Λ�|/�  � D�C��P"��3�  T0 k� ��"��"%�@2 ��A$0 �  �� 	  �  �A��R�6�,
ޣ�|/�  �D�G��X#��3�  T0 k� ��#��#%�@2 ��A$0 �  �� 	  �  �A��R�6�0
ޫ�|/�  D�K��`#��3�  T0 k� ��$��$%�@2 ��A$0 �  �� 	  �  �A��R�5�8
޳�|/�  D�O��h$��3�	  T0 k� ��$��$%�@2 ��A$0 �  �� 	  �  �BA���5�@
޻�|/�  D�S��p%R�3�	  T0 k� ��"��"%�@2 ��A$0 �  �� 	  �  �BA���5�D
޿�|/�  $D�[��x%R��	  T0 k� �� �� %�@2 ��A$0 �  �� 	  �  �BA���5�L
���|/�  (D�_���&R��	  T0 k� ����%�@2 ��A$0 �  �� 	  �  �BA���5�T
���|/�  ,	Fc���'R��	  T0 k� ����%�@2 ��A$0 �  � 	  �  �BA���4�X
���|/�  0
Fg���'R��	  T0 k� ����%�@2 ��A$0 �  �� 	  �  �B����4�`
���|/�  8Fk���(B��	  T0 k� ����%�@2 ��A$0 �  �� 	  �  �B����4�h
���|/�  <Fs���)B��
  T0 k� ��� %�@2 ��A$0 �  �� 	  �  �B����3�p
���|/�  @Ft ��)B��
  T0 k� ��%�@2 ��A$0 �  ��   �  �B��� 3�x
���|/�  �HFx��*B��
  T0 k� ��%�@2 ��A$0 �  ��   �  �B���3��
��|/�  �LF���+B��  T0 k� ��%�@2 ��A$0 �  ��   �  �B�#��3��
��|/�  �TF���+� �  T0 k� �� %�@2 ��A$0 �  ��   �  �B�#��2��
��|/�  �XE����,�!�  T0 k� �$�(%�@2 ��A$0 �  ��   �  �B�'��2��
��|/�  �`E����,�"�  T0 k� �,�0%�@2 ��A$0 �  ��   �  �B�'��$2��
�#�|/�  �dE��	��-�#�  T0 k� �0�4%�@2 ��A$0 �  ��   �  �B�+��,2��
�+�|/�  �dE��
��.�$�  T0 k� �8�<%�@2 ��A$0 �  ��   �  �B�+��41��
�3�|/�  �hE���.B�$�  T0 k� �D�H%�@2 ��A$0 �  �   �  �B�/��<1��
�;�|/�  �pE���/B�%�  T0 k� �P�T%�@2 ��A$0 � ��   �  �B�3��@1��
�C�|/�  �tE���/B�&�  T0 k� �\�`%�@2 ��A$0 � ��   �  �B�7��H1��
�K�|/�  �|E�� 0B�'�  T0 k� �h�l%�@2 ��A$0 � ��   �  �B�7��P1��
�S�|/�  �|E��0B�(3�  T0 k� �p�t%�@2 ��A$0 � ��   �  �E�;��T0��
�[�|/�  ��E��12�*3�  T0 k� �|��%�@2 ��A$0 � ��   �  �E�?�	\0��
�c�|/�  ��E���12�+3�  T0 k� ����%�@2 ��A$0 � ��   �  �E�C�	d0��
�k�|/�  ��E���$22�,3�  T0 k� ����%�@2 ��A$0 � ��   �  �E�G�	h0��
�s�|/�  ��E���,22�-3�  T0 k� ��	��	%�@2 ��A$0 � ��   �  �E�K�	p0��
�{�|/�  ��E���422�.3�  T0 k� ����%�@2 ��A$0 � ��   �  �E�O�	t/� 
���|/�  �E���<3R�/��  T0 k� ����%�@2 ��A$0 � ��   �  �E�O�	|/�
���|/�  � E���D3R�1��  T0 k� ����%�@2 ��A$0 � ��   �  FS�	�/�
���|/�  �!E���L3R�2��  T0 k� �� �� %�@2 ��A$0 � �   �  FW�	�/�
���|/�  �!E���T3R�3��  T0 k� ������%�@2 ��A$0 � ��   �  F_�	�/� 
���|/�  �"E� �\3R�4��  T0 k� ������%�@2 ��A$0 � ��   �  Fc�	�.�(
���|/�  �#E��d4b�5��  T0 k� ������%�@2 ��A$0 � ��   �  Fg�	�.�0
Ϸ�|/�  �$E��l4b�6��  T0 k� ������%�@2 ��A$0 � ��   �  E�k�	�.�8
Ͽ�|/�  ��%E��x4b�7��  T0 k� ����%�@2 ��A$0 � ��   �  E�o�	�.�D
���|/�  ��&E�Ҁ4b�8��  T0 k� ����%�@2 ��A$0 � ��   �  E�s�	�.�L
���|/�  ��'E�$҈4b�9��  T0 k� �C��G�%�@2 ��A$0 �   �   �  E�{�	�.�T
���|/�  ��(E�,Ґ3b�:��  T0 k� �C��G�%�@2 ��A$0 � �   �  E��	�-�\
���|/�  ��(E�0��3b�;��  T0 k� �C��G�%�@2 ��A$0 � ��   �  E���	�-�d
���|/�  � )E�8��3b�<��  T0 k� �C�#4� %�@2 ��A$0 ���   �  E���	�-�l
���|/�  �*E�@��3b�=��  T0 k� �C�#4� %�@2 ��A$0 ���   �  E���	�-�t
���|/�  �+E�D��3R�>��  T0 k� �C�#4� %�@2 ��A$0 ���   �  E���	�-�|
���|/�  �+E�L��3R�?��  T0 k� �C�#4� %�@2 ��A$0 ���   �  E���	�-��
��|/�  � ,E�P ��2R�@��  T0 k� �C�#4� %�@2 ��A$0 ���   �  E���s�,��
��|/�  �$-E�X ��2R�A��  T0 k� �C�#D� %�@2 ��A$0 ���   �  E���s�,��
��|/�  �,-E�\ r�2R�B��  T0 k� �C�#D� %�@2 ��A$0 ���   �  E���s�,��
��|/�   4.@�d!r�1 ��B��  T0 k� �C�#D� %�@2 ��A$0 ���   �  E���s�+��
�'�|/�   </@�h!r�1 ��C��  T0 k� �C�#D� %�@2 ��A$0 ���   �  Dѷ�s�+��
�/�|/�   @/@�p"r�1 ��D��  T0 k� �C�#D� %�@2 ��A$0 ���   �  Dѻ�s�*��
�7�|/�   H0@�t"r�0 ��E��  T0 k� �C�#d� %�@2 ��A$0 ���   �  D�Ôs�*��
�?�|/�   P1@�|"r�0 ��F��  T0 k� �C�#d� %�@2 ��A$0 ���   �  D�˕s�)��
�G�|/�   T1@��#s / ��G��  T0 k� �C�#d� %�@2 ��A$0 ���   �  D�ϖs�)��
�O�|/�   \2@��#s. ��G��  T0 k� �C�#d� %�@2 ��A$0 ���   �  D�חs�(��
�W�|/�   `3@��#s. ��H��  T0 k� �C�#d� %�@2 ��A$0 ���   �  D�ۗ��'��
�_�|/�   h3@��$s- ��I��  T0 k� �C�#t� %�@2 ��A$0 ���   �  D��� '��
�g�|/�   l4@��$c , ��J��  T0 k� �C�#t� %�@2 ��A$0 ���   �  D���&��
�s�|/�   t4@��$c$+ ��J��  T0 k� �C�#t� %�@2 ��A$0 ���   �  D���%��
�{�|/�   x5@��%c,+ ��K��  T0 k� �C�#t� %�@2 ��A$0 ���   �  D����$�
���|/�   �6@��%c0* ��L��  T0 k� �C�#t� %�@2 ��A$0 ���   �  D����$�
���|/�   �6@��%c8) ��M��  T0 k� �C�#�� %�@2 ��A$0 ���   �  D���%�
��|/�   �7@��&c<( ��M��  T0 k� �C�#�� %�@2 ��A$0 ���   �  D���%� 
��|/�   �7@��&cD' ��N3�  T0 k� �C�#�� %�@2 ��A$0 ���   �  D���&�(
��|/�   �8@��&cH& ��O3�  T0 k� �C�#�� %�@2 ��A$0 ���   �  D���&�0
��|/�   �8@��'cL% ��O3�  T0 k� �C�#�� %�@2 ��A$0 ���   �  D���'�8
��|/�   �9@��'�P$ ��P3�  T0 k� �C�#�� %�@2 ��A$0 ���   �  D�#��'�@
��|/�   �9@��'�X$ ��Q3�  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�+��'�H
���|/�   �:@��(�\# ��Q3�  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�3��(�P
���|/�   �:@��(�`" ��R3�  T0 k� �C�#�� %�@2 ��A$0 � .�   �  D�7��(�X
���|/�   �;@��(�d! ��R3�  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�?��)�d
 ��|/�   �;@��(�h  ��S3�  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�G��)�l
 ��|/�   �<@��)�l ��T3�  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�K��)�t
 ��|/�   �<@��)�t ��T�  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�S��*�|
 ��|/�   �=@��)�x ��U�  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�[�� *��
 ��|/�   �=@��)�| ��U�  T0 k� �C�#�� %�@2 ��A$0 � ��   �  D�_�� *��
 ��|/�   �=@��*�� ��V�  T0 k� �C�#İ %�@2 ��A$0 � ��   �  D�g�d +��
�|/�   �>@��*�� ��W�  T0 k� �C�#İ %�@2 ��A$0 � ��   �  D�k�d +��
�|/�   �>@��*�� ��W�  T0 k� �C�#İ %�@2 ��A$0 � ��   �  D�s�d +��
�|/�   �?@��*�� ��X�  T0 k� �C�#İ %�@2 ��A$0 � ��   �  D�{�d +��
�|/�   �?@��+�� ��X�  T0 k� �C�#İ %�@2 ��A$0 � ��   �  D��d ,��
'�|/�   �@@��+�� ��Y�  T0 k� �C�#԰ %�@2 ��A$0 � ��   �  D�T ,��
/�|/�   �@@� +�� ��Y�  T0 k� �C�#԰ %�@2 ��A$0 � ��   �  D�T ,��
7�|/�   �@@�+�� ��Z�  T0 k� �C�#԰ %�@2 ��A$0 � ��   �  E��T ,��
?�|/�   �A@�,�� ��Z�  T0 k� �C�#԰ %�@2 ��A$0 � ��   �  E��T ,��
G�|/�   �A@�,�� ��[�  T0 k� �C�#԰ %�@2 ��A$0 � ��  �  E��T ,��
K�|/�   �B@�,�� ��[�  T0 k� �C�#� %�@2 ��A$0 � ��   �  E��T,��
S�|/�    B@�,�� ��\�  T0 k� �C�#� %�@2 ��A$0 � ��   �  E��T,��
[�|/�    B@�,�� ��\�  T0 k� �C�#� %�@2 ��A$0 � ��   �  E���T-��
c�|/�   C@�-�� ��]�  T0 k� �C�#� %�@2 ��A$0 � ��   �  E����-�
k�|/�   C@�-�� ��]�  T0 k� �C�#� %�@2 ��A$0 � ��   �  E�ü�-�
s�|/�   C@�-�� ��]�  T0 k� �C�$� %�@2 ��A$0 � ��   �  E�ǽ�-�
{�|/�   D@� -�� � ^�  T0 k� �C�$� %�@2 ��A$0 � ��   �  E�Ͼ�-�
!��|/�   D@�$-�� � ^�  T0 k� �C�$� %�@2 ��A$0 � ��   �  E�ӿ�-�$
!��|/�   D@�(.�� � _�  T0 k� �C�$� %�@2 ��A$0 � ��   �  E����-�,
!��|/�   E@�(.�� � _�  T0 k� �C�$� %�@2 ��A$0 � ��   �  E����-�8
!��|/�   E@�,.�� � `�  T0 k� �C�#4� %�@2 ��A$0 � ��   �  Er���.�@
!��|/�    E@�0.�� � `�  T0 k� �C�#4� %�@2 ��A$0 � ��   �                                                                                                                                                                              � � �  �  �  c A�  �J����  �     6 \��� ]�	n	n � �  <  K K      � �p�     PR �p    �	           	 Z           P�    ���   0
% 
           -p�   � �     � α�     -�� �~    ����    � �        Z          ���     ���   0
           ��   1 1     ��3     � ���    
T�   	            	 Z           @�    ���  P
	         ���   � �
	    ���    ��4� ��    	�I   	            # Z           @�    ���   P	         ����  ��	      .�r�    �����r�                               ���               1  ���    P             �      �         B        �                      ��                                       ���   �                          Oh0          V ��[     O:� �s�    ��              
 
   ��         �  �  ��@   (
          7�~        j �@�     7W �C    R��    � �        
    ��        �  �  ��@   	@

           ��          ~ �6�      �    ��                  �          �@     ��H   H	$
          l��         � �cf     lU� �]    ] _                
  � �         	  �  �  ��B   H
	!          �� ��	     �7     Q��    r��                       ���        
       �  ��@      0            �     �         �        �                      ��                                       ��@   �                               ��      �                                                                           �                               ��        ���          ��                                                                 �                         ���T  ��        �=Z    ���T=Z         "                   x                j  �   �   �                               ==       �,   ��    ,   (�    ��                                      . (        �                           - ����� O 7  l �    ��            
  	     
  #   {	� �}�D       �  }` �D  }� � a� 	_� �t� 	`� u� 	a u� ��  }` �� }� ��  }` פ v` J n� J$ n� H� n� L�  s@ 
� V� 
�\ W  
�< W� 
� W� 
�\ W� �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ � }`���� � 
�| V ���� � 
�� V� 
�\ W  
�< W� 
�� W� 
�| W����� � <� d  <�  d@ �d �`� �� a� ��  a� �� b  �D �[� �D \� �d  \� ɤ  ]  �� ]` )� `e� *D f����� � 
�| W  
�< W� 
� W� 
�\ W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����          ������  
�fD
��L���"����D" � j  "  B   J jF�"     �j  B
 ��
��
��"    "�j�� , " �
� �  �  
�  1��  ��     � �  �    -��  ��     � �           ��     � �          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  �$      �� � �  ���        � �T ���        �        ��        �        ��        �    ��     ��� h��        ��                         �$ ( 	�� ��                                     �                ����          
   2 ����%��     2               85 Sanderson    sh     0:04                                                                       5   0      �bS �BS �"$ � �" � �"" �" �*$8 �*4P � "P
kj1 krc�[/ c�kB� B�( B�# �cV: J� � � J� � �J� � �c~ � � c� � �c� � � c� � c� � � � � �	� � �	� � �� � �� �� � � � �-!"�- ""�!#"�$*�%"� � &"� �'� � �(
� � �)"$ � �*" � �+"" � �,"
 �-*$* �.*4B �/"B � 0*Or �1*(z �  *Hr �3"' �4*$G � * _ � *G �7"' � *G � * _X :"K �X  "K �<!� |8 ="I �H >"P �P  "O �                                                                                                                                                                                                                         $ �             @ 
     &�      Q P E a  ��                   	 �������������������������������������� ���������	�
��������                                                                                          ��  �4� >  ������������� �!�"�#�j�k�&�'�(�)�*�l�m�n�.�/�0�1�o�p�q�5�6�0�1�M�r�N�:�;�0�1�<�`�>�1�?�@�A�B�s�D�A�E  �~�, -  * Z�� �@,@r�@� �&��;��                                                                                                                                                                                                                                                                                                                                 ��@��A                                                                                                                                                                                                                                      �  	  #    ��  D�J    	 �                             ����������������������������������������  ����������(�                                                                                                                                       �      � 8    ]        �        � ��          	  
 	 
 	 	 ���� ����������������� ����������� ����������� ���� ������������������������������� � ����� ���������� �� ��� �� ������ � �������������   �������������� ������������� � ��������������� ����������� �� ��������������������� ��           1                   �         	� �	  H�J      �  	                           ���������������������������� �����������������������                                                                                                                                              �        �      �        !    ��             
 	  
	 
 	 	 ����������� �   ����  �������������������������� ���������  ���������� ������� �����   � �� ����� ���������������� ����������� �������� ����  ���������� �������������������� �� ������������������������  ���               x                                                                                                                                                                                                                                                             
                                                 �             


             �   }�         �#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�"" , J >               	                  � h3�� �\                                                                                                                                                                                                                                                                                    2-1n	n  �)F                      e            m   D             c                                                                                                                                                                                                                                                                                                                                                                                                                 � q� �  � ��  �  ��  � #��  � #��  � ��  ����������(����������������u�����������g����|�                ��              	 	 �   & AG� �  �   
              �                                                                                                                                                                                                                                                                                                                                      p B C    �          &             !��                                                                                                                                                                                                                            Y   �� �~ ���      �� B 	     ���� ����������������� ����������� ����������� ���� ������������������������������� � ����� ���������� �� ��� �� ������ � �������������   �������������� ������������� � ��������������� ����������� �� ��������������������� ������������� �   ����  �������������������������� ���������  ���������� ������� �����   � �� ����� ���������������� ����������� �������� ����  ���������� �������������������� �� ������������������������  ���             $�����������������������������������������������f���f���f��ff��ff��UX����fffffffffffff�ffffffffff����ffl�fff�ffffffffffffffffflff������������ʪ��l���fl��f�h�f�k�������������������������������������������������������������������k���gW��ey�k���fkf�fff�fff�fffj��wUUUU�w��lffjfffffff�ffffffl�u�˦U��[�fj��ff�fff�ffffffff��Ƽfjk��fk��ff�̶fjf�fjfffkfffjfffj�����������������������������������������������������������������ff˩fi��jz˜ev��Ŧ���[W�gW��hW���w������w�w�xw������ʗyƜ�Z���X��wW�������������l���l���l����xw�ff�U�f��\fjj[fj�[fi�[fhy\fiz|�������������������������������������������������������������������k�u���U�U�UgU�Ue[�U���U���U���U��uUx�UwUUW�UUXwUW��UW��Uuz�UUX���wUx�uUxx��wxx��wxw�wwwU�w�U�Uw{ʨy��U�y�UkYz�ky���yuUzy��zZ�U�������������������������������������������������������������������iu�vj��Uz��uU����ɚ�U���u{���YuUx�U���U���Wuy�ww���wx���w�ɇX��wU���ww��UXuxwY��x��w���w������yl[��j[��j[��jU��i���h�U�g�w��x��������������������������������������������������������y��f�ffff���w������������x�����wXgUUxkUX�f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff��$�&    0          � ��                      B     �   ����������      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$     `d  �@    �f ��    �f �$ ^$ �@      �       �     �  h 
� � v                  x          �            �������2     �   ��     �   �$ ^$   a      �      � ��     � �$ ^$  	n   x x        �  �              ���             }PS   yL  ��������������������������������GvdDGw6wGwcfGwsfGwv6Gww6GwwcGwwcDDDDwwwwffffffffffffffffUUUUttttDDDDwwwwffffffffffffffffUUUUtttwN���t���wN��wt��wwN�wwt�wwwNwwwtGwweGwwU�tvf�wff�Fff�Fff��df��ffwwwwUUUUffffftDDft33gt5egt6Vgt5gwwwwUUUUffffDDDD3333eeeeVVVVwwwwwwwwUUUUffffDDFF35FfefDDVVFUufGfwwwwGwwwGwwwUUUUffffDDDDUUUUffffwwwwwwwuwwwuUUUUffffDDDDUUUUffffwwwwUUUUffffddDDfd33DD6VUd5eft6WwwwwUUUUffffDDGf35GfVVGvefGv6VGvwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwN�Fft�FfwN�dwt�fwwNGwwtGwwwDwwwtwt6Wwt5gwt6Wwt5gwt6Wwt5gtt6Wwt5gDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD6VGd5fGd6VGd5fGd6VGd5fGd6VGd5fGdFt5gFt6WFt5gFt6WFt5gFt6WFt5gFt6W5fGw6VGw5fGw6VGw5fGw6VGw5fGG6VGwgwwwvwwwwgwwwvwwwwgwwwvwwwwgwwwvGt6WGt5gDt6WDt5gND6WNt5gNt6WNt5g6VGd5fGf6VGw5fDD6VGU5fGf6VGf5fGfDDDDffffwwwwDDDDUUUUffffffffffffFt5gft6Wwt5gDD6WUt5gft6Wft5gft6W5fGt6VGt5fGD6VGD5fD�6VG�5fG�6VG�GwwwDwww�Gww�Dww~�Gww�Dww�DGw~�DNt6SNt5fNt6VNteeNwFVNwteNwwFfffd3333ffffVVVVeeeeVVVVeeeeffffDDDD333DffcDVVSDeecDVVSDeecDfVSDFecDUUUUDDDDDDDDDDDDDDDDDDDDDDDDDDDDD333D6ffD6VVD5fdD6VDD5fDD6VDD5fD3333ffffVVVVDDDD33335UUU5Vff5VDD3333ffffVVVVDDDD3333UUUUffffDDDD6VGfefGfVVGwDDDD3333UUUUffffDDDDffffffffwwwwDDDD3333UUUUffffDDDDft5cft6Vwt5eDDDD3333UUUUffffDDDD3333ffffeeeeDDDD3333UUUVffeVDD5V333DffcDeecDF6SDD5cDD6SDD5cDD6SDD333D6ffD5eeD6VVD5eeD6VVD5ffD6Vd5fG�fVG�efG�VVG�edw�VGw�dww�Ffffffffwwwwwwww����DDDDNNDD��������gwwwwwwwwwww��wwDDGwDDDw��DG���Dwwwwwwwwwwwww~��wwn�wwvwwwwgwwwvFfffFfffCeeeCVVVCeeeCVVVCeeeCVVVfDDDfDDDfDDDVDDDfDDDVDDDfDDDVDDDDfSDD5cDD6SDD5cDD6SDD5cDD6SDD5cDD6VDD5fDD6VDD5fDD6VDD5fDD6VDD5fD5VDD5VDD5VDD5VDD5VDD5VDD5VDD5VDDDDDDDDDADDDADDDDDDDDDDDADDDADDDDDDDDDDDDDDwDDDDDDDDDDDDDwDDDDD5VDD5VDD5VDD5VDD5VDD5VDD5VDD5VD5cDD6SDD5cDD6SDD5cDD6SDD5cDD6SDDDDfDDDfDDD5DDD6DDD5DDD6DDD5DDD6fffdfffdeeedVVVdeeedVVVdeeedVVVdCeeeCVVVCeeeCVVVCeeeCVVVCeeeCVVVfDDDVDDDfDDDVDDDfDDDVDDDfDDDVDDDD6SDD5c3D6VfD5eeD6VVDVffDDDDDDDDDDDD3333ffffeeeeVVVVffffDDDDDDDDD6VD35fDffVDeefDVVVDfffDDDDDDDDD5VDD5VDD5V335UUU5UUU5UUUVfffDDDDDDDDDDDD3333UUUUUUUUUUUUffffDDDDDD5VDD5V335VUUUVUUUVUUUVffffDDDDD5cDD6S3D5ffD6VVD5eeD6ffDDDDDDDDD5fD36VDfefDVVVDeefDfffDDDDDDDDDDDD5DDD6DDD5DDD6DDD5DDD6DDD5DDD6eeedVVVdeeedVVVdeeedVVVdeeedVVVdwwww�twwww~ww�w�wtwwtwwww~w�wwwwDDDDDDDDDADDDDDADDDDDDDDDDDtDD4DDqt4DDDD4DDsDDDDDDDDDDDD7AtCADADDADADDDDDDDADDDADDADqDADqDDDDDADDDADDDAADAADqADDAGADDDDwwwywww�www�www�www�www�www�www�������������������������www�www�www�www�www�www�www�www����������������������!�����!�-����������!-�����������!�����wwwwwwwtwwwOwww�wwt�ww�wwOGww�D��������������-��������������������������!����������-������NNNNNNNNNNNNN���FfwfDDDDDDDDDDDDNNNDNNNDNNND����gvftDDDDDDDDDDDDwts"wwB2ww22ws#Cws#4ww2twws�www�www�www�www�www�www�www�wwwywwww��������wwww������!��������wwwwww��w��w2��w���w��t���(�wy���������y���w�����y��Gwwwwt33Dt343CeeeCVVVEeeetVVVvEee�DVVzDFf�DDDfDDDVDDDe333VfffeeeeVVVVffffDDDDDDDDDDDD3333ffffeeeeVVVVffffDDDDDDD5DDD6333efffVeeeeVVVVffffDDDDeeedVVVdeeedVVVGeedgVVDzfdD�DDD�Df��NvDGN�DNN�DND~DGD��NDNt�DDDN#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFw"GC42wsDCwt�Cwt��ws�DGt�T7DfEGt{�Gwz��w���wt�Gw��wt�Gw�wtw�{�Gww��w��w2��w���w��w���x�wy����wwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wt3Gwt4wCGGttwG4�twO�wGt�GwE��wTfNw~D�����������������DD��ww�N��D�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wfuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGy�wwy�wtw�wOw�w�w�D�w2?�wCOGww�Dwwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGww23ws""wr22w244w#tD�t3~�}�ww}O3#�w""7w##'wCC#wDG2w3G~������wwwwVtwwUvwwenwwvWwwv�wwtwwtGww�3#�w""7w##'wCC#wDG2w3G~��7���wwww}�ww}�ww}�www�www}www}wwwwwwwr��ww��ww���w4��w��ww��www}ww'r'ww"GCw2wswCwtwCwtw�wswDGtwB'tww"w#w�2w�3w�3wG4wtGDwww"wr!r'wrwuUUG4wwD4wwCtwwCtww7tww7twwGtww8�3�3�3�8�3�3�33333"2#333"33UUUUwwwtwwwtwwwtwwwtwwwtwwwtwwwt��33�?33�?33�?333333#23323#3UUUUwwwwwwwwwwwwwfgvwwwwwwwwwwwwUUUUwwwtwwwtwwwtfwfdwwwtwwwtwwwtUUUUwwwwwwwwwwwwwwwwwwuwwwWwwwwwUUUUwwwWwwwWwwwWwwuwwwuwwUuwwwUwC�38C838C�38C833C332C"33C2#3UUUUwww~www~www~www~www~www~www~UUUUwfwnwvw~wfw~wvw~www~wfw~wgw~UUUUuwwwuwwwuwwwwWwwwWwwwWuwWUwwUUUUwwwwwwwwwwwwwwwwWwwwwwwwwwwwUUUUwwwdwwwdwwwdwwwdwwwdwwwdwwwdUUUUwwwwwwwwwwwwwwwwwwwwwwwwwwwwUUUVwwwvwwwvwwwvwwwvwwwvwwwvwwwvGtwwGtwwGtwwGtwwGtwwGtwwGtwwGtwwwwwtwwwtwwwtwwwtwwwtwwwtwwwtwwwtww�www�www�www�www�www�www�www�w�www�www�www�www�www�www�www�wwwwwwdwwwdwwwdwwwdwwwdwwwdwwwdwwwdwwwvwwwvwwwvwwwvwwwvwwwvwwwvwwwvGtUUGTffGTffEdffEdffFdffFdffFdffUUUUfffffffffffffffffffffffff���UUUUffffffffffffffffffffffff����UU�Uff�eff�Vff�Vff�fff�fff�fʦ�f�UUU�fff�fff�fff�fff�fff�fff�fffUUUUffffffffffffffffffffffffffffwwwdwwwdd333d333d333d333d333dwwwwwwww33333333333333333333wwwvwwwv33363336333633363336FdffFdffAC333C333C333C333C333��������33333333333333333333�f�f�fFf�33�333�333�333�333�3�fff�fff33333333333333333333ffffffff33333333333333333333333d333d333d333d333d3333����wwww333333333333333333333333����wwww333633363336333633363333����wwwwC333C333C333C333C3333333����wwww33�333�333�333�333�33333����wwww�����<��5UUU5UUSU553SS2#33"532 5�����<��5UUU5UUUU555SSSS33333��������UUUUUUUU5555SSSS3333��������UUU�UU_�55=�SS]�33;������l���eUUUUUUSU552SS2#S3"3S2 0�����<��5UUU5UUSU552SS2#33"332 0����ȩ��S�UUU��US:�U59��38��009������<��UUUUUUUU5555SSSS33333������ÓUUX�UUS�SSX�553�338�003�����3���UUUU5UUUU555SSSS33333�����̚�Ue�5UX�U5Y�5X��S9��3����������UUUUUUUSU5523S2#"302 0�����<��5UUU5UUSU552SS2#33"302 0�����<��5UUV5UUUU555SSSU33353��������UUUUUUUUU5553SSS33330����l���eUUSUUU3SSS%U3"5S2#3S" "#  %                     200            "          "                         0;�  ��  �� ��  ۰  ۰  ��  ��                          #                         P"R                         "#                       "#  "                    0"                                                    �  9                     �#�� ��� ��� ��  �       02(�" �  � ��0(�������� �����   �                    "                         205            "         R 20R                                                                                    ��  ��  �� �� �  �  �  �   �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��  �S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����      �� �� �� ܈ ܈ ��  �   �  �����݈�<̈�������             ������݈��͈���     �       �������݈�8���        ��������8���������   �  ��  �� 3� ������ ���  �� �� �� � ܙ ܙ�ܙ ܙ����؈���؈���؈���Ù��ݙ��ݙ��݈��������������������̈��܈����̈����������������������͈������݈����������͈���������ܙ��	�������� ��� ��� ��� ��� ��� ��� ���  ܙ ܙ ܙ ܙ ܙ ܙ ܹ �ə��ݙ��ݙ��ݙ��ݙ��ݙ��ݙ��̙������������ܙ��ܙ��ܙ��ܙ��̙�����������ݙ��ݙ��ݙ��ݙ��ݙ��̙����ə��ə��ə��ə��ə��ə��	��������� ��� ��� ��� ��� ��� ��� ��  ��  �  �  �                ����	���ܹ����	������      �����������͙��������      ���������ə��ܙ���� �      �����������͙���̼����      � ��  �                     wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "! ""! " ""  "!  "       " ""                       ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                                               "! ""! " ""  "!  "       " ""                 ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �        "!  "" "  """     " ""   "" !"""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                       �  �  ��� �                     �  �˰ ˻� w�� k}� gw� z�� ��� ��� ��� ��� ��  �� ���"�ȍ�̽�"��4  4H H� D�� X�D X� Ą  ��" 
��  "  "" ""  ��    �   ��  ��  ��  ��  ��  ̐  ��  �0  �0  �0  T   C   3   �   ��  +�  ""  ""� /�� / �    ��                 �   �                           �   �  "������"    /   �  �   ��                             �                        ���� ��� ����                                                                                                                                                                                                                                              �   �  �  �� ",� ."� "�  �3  >3  �4 
�� �� "�""�"�(�"�   ��� ��� ��� �g} ��װ�vz��gz�8ʪ�C���T8��U]��,ʌ�"ȩ "ː �    �   �   "  "  "  �" ��  ��ɜ�ʨ�����,���/���������     �        �   �   �   �   ��  ��  ��        �       �    �             �  ��  �  �  ��     ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����            �����                                                                                                                                                                                                                                  �  �   ��  �   �  �  �  ��  ��  ��  I�  T:  UJ  T   T  T  J  T�  �� 
�� � �  �˰ ��� ��p���p��� ��� ˹� ̻� �̙ ̼� ˼� �ܘ �٪�؋�Ѓ=�Ш3� �C  �0  ��  ;"� "/ �� ��  ��� ,� ""/ """  ���     �      �                           �  ��  �  ��  �                           �   �   �   "   "   "  !�    ��                                                               �               �  �  ��  �   �   �                                                                                                                                                                                                       "  �� �� �������ɪ �̙ ��  ��  �  �  �  �  �  	�  �  D  D  3   3   3   �   �   �   �  � ��+  �"     �        ��  ��  ��  ��  �� 	�p ����ə��������̻��˻ ̻� ̻  ˻  ��  ��  D�@ D�T UZ� 4U�@3D�@�DJ��K�� ̻�(̰�*������,�"�""!�"! �� �                      "   "  "                  �  �      �   �   �             �   �  "  "  "  �"  ̰  ˰  ��  ��  �               �   �                             ��� ���� ��                                                                                                                                                                                                       �  �  �  �  w  
�  ��̙̊��̉��̌ݼ̌ݼ̘ͼ� ��� �� ��� �8��33�33�H�U���M����٘лڭл,���,���"� �     �    �   �   �   �   }   ��  ��  ɘ� ��� �ܚ��٩�̽��̽�˹��.��""�3�"33��33� C�: �D3��C�Ћݸ�ؙ��ݪ���̲�򻲿�"/�����   �    	   	   	   	                                         �     �     �   �   �   �   �   �   ��  ���  �  � �                     ��� ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �  �� ̽ �� �w 
�� ���������̸��̽���ݼ����� ��� ���
8�ȣ3���333�333�C0TUT0�C� �ݰ ��� 
�� ,�  ,�  �"� �  ��           �   �   �   �   ��  ��� ������̚�˚��ک���ۻ�ݻ���� �ݰ �"  3:  3:  33  33� DC0 T=� �ۀ ��� 
�� ,�  +�  �"� � ����   �       �   �   @   �   �   �   �   �   �"  ""  !� �� ��  �               �   ������  ��                      �   �                      �������  ���    �        � ��                    ���� �                                  �  � �                       � �� �                 ��� "   "   "   "        ��   �  �  �� �  ��  �             �  �                                       �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                 �� �̽���ݪ۽w�}�֪�vv���p��� ��� 
�" ��" �""/�"" �����                     �   �                      �������  ���    �                    ��  ��  ���  ��  �  �  �   �                                                                                                                                                                              �� ��� ��� ww� ��� vv� w�  �  �  �  �   �   �  3� ;� <� "� "# "�."��! ���� �� ��� �   �                           �   �   ��  ��  ��� ��� ��� ������̰�ۻ���8��3�@38� 3�@ 8�P H�  8�  ��  ��  �� �"  ""  "! � ����                              � �� ��� ��    ̹� ˘P ��@ �U@ UT@ T30 33  30       �  ��  ��  ww  ��  vv  w                �                        ���� ��� ����                  �  ������� ��                                                                                                                                                                                                                     �  �� 
�� �������˚��̻ۈ�˽��+T��(T�""U�2"EJ�"T�3 EJ� Z� Z� �3 "�� ,�� ʡ "��"""""" ��  �        �  ��� ܽЪ��p��}`�wg`�pw ��  ً  ��  ��� ۽� ۈ�  ��  �� �۰ >�� >"  0�  0"   "  �� " �  ��  �   /��  �   ��          �   ��� �� ����                   �                    � �               �   �                �   �       ��  � �                    ��  ��  ��                                                                                                                                                                                                                                        �   �  �  ��  ̽  ��  �w 
������ə����̹��̻+�̉������ �� ��� H�� DH� 3ES 33 �35 ݘ� �ۿ������ʸ��˽����"�����            �   �   ��  ��  ������鈙����ܻ��ۙ��٪��͉��ͻ���۸��  ��  �:� 3:� 34� �D� Ӆ]��EͰ�ۘ��� ڭ ,°�+� ��/ �  �  �   �   �   �   �   ��       �                   �   �          �                           �                                        ��  ��   �   �   �               �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                               DN 䤤�J��@J��@J��@J��ND��N����    
�   ̜ ����� �Q�    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                         "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""�������������������""""���������D""""������D�J�""""��������D�""""������JDADJ�J�""""������DA�D�JJ�""""��������AA�A""""��������AA�A�""""��������������J��J��"""$���4���4���4���4���4���4������������������333DDD���������������D����3333DDDDA�D�H�H�D�H����3333DDDDAAA�H�H�D�H����3333DDDDH��������D������3333DDDDH�DH��H��H��H�D�����3333DDDDHH����������D����3333DDDDAAA�D��H�D�����3333DDDDD��H�����HDD����3333DDDDH��H��H��D���H�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""��������������������""""����DDD�III""""������A�I�I""""����������IAIA""""�������DI���""""������DI�I�""""�����I�DA�I��I�""""�������DI���""""������DI�I�"""$���4���4���4���4���4���4������������������333DDD���������������������3333DDDDDLL��LDD�D����3333DDDD�LLDLLLD��L����3333DDDDLALALLLL�L�L����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD�L��L��L��L���L�����3333DDDD���D�L�DD�����3333DDDDL�L�L�L��L�D����3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H��                                 ((((( 
	(((( """"��������AA�A                	 
  (%($(#("(! (((ADA�LL��L�D����3333DDDD   ������� ������� �� ������������  (((((2	10/(.(-(,(+LL����������D����3333DDDD   ��	�
��������    ��������������������  (!()(%($ :198(((7(6(5""""����������A������        ����     ! " # # $! % &  ����  ' ((B(A(@?>108(=((( (<""""�������I�I������ ) * + , - .  �Ӥ�  / 0 � 1 2�� 3 4  ��� / 5 6+*) S S SRQPO(( (N(,(+(M(.L""""�������I��D���I�������     7 8 9 : : : : : ; < = = = = = = > ?::::: @ A B     ^]\[Z SY(X(W(V(U(5(N((7�D�M�D���M������3333DDDD C CC 7 8 DD  E F G H         DD  E F G H A B CCC ihgfedcb(a(((V((`D�M�A�����MD�����3333DDDD    7 8�#� ���%��        ��!���%�� A B    utsrqponbml((+(k(M 
""""�����AMAD������   Q 7 8                       A B(Q   �� � �|{znby(6(5(Mxw""""������������������ V W X 7 8                       A B(XWV � � � � � �����b(� 
xwwfFfFDfFFfFffdFffff3333DDDD V W \ 7 8                       A B(\WV � � � � � ����� ��ww�(+DDFFDfFFfdFffff3333DDDD V W ] ^ _ ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` ` a b(]WV � � � � ������ ���((W(�""""wwwwwwwGGD V W c d e f g h i j V W  k h i d e f l V W(j m(h(g(f(e(dcWV� � � �� �������l(�(a(�""""wwwwwwqwAqwAwA V W n o p q ] r s t V Wn ] r u o p q v V W(t(s(r(](q(p(onWV � � � � � � ������y(�(�""""wwwwqwqAwAqAqAq V W w f g h i d e f V W x i d e f k h y V W(f(e(d(i(h(g(f(QWV ��� � � � ������((�l(=A�A�A�A��LD�����3333DDDD V W z { ] r u o p q V W | u o p q ] r u V W(q(p(o(u(r(](q }WV����� � � �����((�(( �A�LDL�L�D�L�����3333DDDD V W ~  � � � � � � � � � � � � � � � ���(��(��(�(�((~WV � � � ��� � �����(-(5(Xx""""wwwwwwDGAD � � � � � � �  �   �  � �� �� �  � �� � � � �� � � � � ��� �����(�xww""""wwwwqqDAAq �     � � � � � � � � � � � �����������    � �� � � ��� �����ww�(""""wwwwwwwGGwGGwGwGw � � � � � � � � � � � � � � � � ����������� � � � ���� � � ��� ������(+((�UQUUQUUQUUQUUUDUUUUU3333DDDD � � � � � � � � � � � � � � � � � �� � � � � � ��� � � � �� � � � � ��� �����(W(�m(`DEQQUUDUTEUUUU3333DDDD � � � ��� � � � � ��� � � �� � ���� � � � � ���� � � � � � ��� � �� ���(a((M""""������������������������ � � � � � � � � � � � � � � � ��� � � � � � � � � � �� � � �� ���� � � � � ���(-(� 
(�""""�������DAADAI � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � ���� � � � � � ����(( (-(��A�AM�M�DM��M334CDDDD � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � � �� � � � � � � � ���(X((6(5DD����M��DM�����3333DDDD � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �� � �� � � � � � ���l((�x""""wwwwwwDGqGq � � � � � � � � � � � � � � � �� � � � � � � � � � � �� � � �� � �� � � � � � ���yxww""""wwwwwwwGwwDGwwwwwwww + � � � i � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����ww�(+ADAH�DJ�H�H�����3333DDDD � W � � u u �  � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � ������((W(��H��J�AD�DH�D����3333DDDD333333333333333333333333333333333333333333333333333333333333����  
�fD
��L���"���""""�������DD������D" � j  "  B   J jF� ����
��� �����
���� ����
��� �����
��� 0 q""""������DH���""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqqbS �BS �"$ � �" � �"" �" �*$8 �*4P � "P
kj1 krc�[/ c�kB� B�( B�# �cV: J� � � J� � �J� � �c~ � � c� � �c� � � c� � c� � � � � �	� � �	� � �� � �� �� � � � �-!"�- ""�!#"�$*�%"� � &"� �'� � �(
� � �)"$ � �*" � �+"" � �,"
 �-*$* �.*4B �/"B � 0*Or �1*(z �  *Hr �3"' �4*$G � * _ � *G �7"' � *G � * _X :"K �X  "K �<!� |8 ="I �H >"P �P  "O �3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD������������������������������������������������������������������������������������������� �!����� � � �m�n�|�}�c�d�v�w��� � � � � ��������������������������������������"�#�j�k�&�'�(����� � � ������������������ � � � � ��������������������������������������)�*�l�m�n�.�/������#��<�G�T�J�K�X�Y�U�T��a� �b� ��������������������������������������0�1�o�p�q�5�6����������������������������������������������������������0�1�M�r�N�:�;����������������������������������������������������������0�1�<�`�>�1�?����������������������������������������������������������@�A�B�s�D�A�E���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������/�.�7� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������2�0�.� ��"������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������;�K�Y�[�S�K��1�G�S�K����������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                