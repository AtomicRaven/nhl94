GST@�                                                            \     �                                                ���� Q   @��             dT 2�������J���vr�����    ����        6     #    ����                                d8<n    �  ?     ������  �
fD�
�L���"����D"� j   " B   J  jF�"    
 �j, 
���
��
�"  ""B�j��" 
 ��
  �                                                                               ����������������������������������      ��    bb= QQ0 4 111 44            		 

                     ��� �   � �                 nn ))
         88�����������������������������������������������������������������������������������������������������������������������������oo    go      +      '           ��                     	  7  V  	                  �            8: �����������������������������������������������������������������������������                                $`  �   ;  ��   @  #   �   �                                                                                'w w  )n)n
  �    6�   �1��F!} "� �! @�� ~ ��6 +�� ~ ��6��� ~ ��6 "�� ~ ��6�!# �!& �f�n|�~ 2� Ø �6 *^��g 2@y� O  �Z�} |��g>ͪ <2� 7?Õ 7?2 `2 `2 `2 `2 `2 `2 `2 `2 `����: �?0�� ~ ��6 (�� ~ ��s� ��: �?04��[̀�0W�� ~ ��r N#�� ~ ��qx� z�W��! @� ��: �?0<�! {�'�òƤ�� ~ ��w V�� ~ ��r��� ~ ��w #V�� ~ ��r�! @� ��: �?���[}�o|� g~��8�8�8! {�ò�L�� ~ ��w V�� ~ ��r(B��� ~ ��w �� ~ ��r(+��� ~ ��w �� ~ ��r(��� ~ ��w �� ~ ��r�! @��: �w(�� ~ ��6 +�� ~ ��6 �?0�� ~ ��6 (�� ~ ��s� �:� =2� !} "� ��Ø ! {�o~o�%��%��%��%��%�H�	>ê {���#�#��� �E � �                                                                                                             ddeeeefffffgggghhhhhiiiijjjjjkkkklllllmmmmnnnnnoooopppppqqqqrrrrrsssstttttuuuuvvvvvwwwwxxxxxyyyyzzzzz{{{{|||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ cddddeeeefffffgggghhhhhiiiijjjjkkkkkllllmmmmnnnnnoooopppppqqqqrrrrsssssttttuuuuvvvvvwwwwxxxxxyyyyzzzz{{{{{||||}}}}~~~~~������������������������������������������������������������������������������������������������������������������������������������ ccccdddddeeeeffffgggghhhhhiiiijjjjkkkklllllmmmmnnnnoooopppppqqqqrrrrsssstttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{|||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ bbbbccccddddeeeeffffgggghhhhhiiiijjjjkkkkllllmmmmnnnnoooopppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxxyyyyzzzz{{{{||||}}}}~~~~������������������������������������������������������������������������������������������������������������������������������������ aaaabbbbccccddddeeeeffffgggghhhhiiiijjjjkkkkllllmmmmnnnnooooppppqqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ````aaabbbbccccddddeeeeffffgggghhhhiiijjjjkkkkllllmmmmnnnnooooppppqqqrrrrssssttttuuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ____````aaabbbbccccddddeeeffffgggghhhhiiijjjjkkkkllllmmmnnnnooooppppqqqrrrrssssttttuuuvvvvwwwwxxxxyyyzzzz{{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� ]^^^____````aaabbbbcccddddeeeefffgggghhhhiiijjjjkkkllllmmmmnnnooooppppqqqrrrrsssttttuuuuvvvwwwwxxxxyyyzzzz{{{||||}}}}~~~����������������������������������������������������������������������������������������������������������������������������������� \\]]]^^^^___````aaabbbbcccddddeeeffffggghhhhiiijjjjkkkllllmmmnnnnoooppppqqqrrrrsssttttuuuvvvvwwwxxxxyyyzzzz{{{||||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� [[[\\\]]]^^^^___````aaabbbccccdddeeeffffggghhhhiiijjjkkkklllmmmnnnnoooppppqqqrrrsssstttuuuvvvvwwwxxxxyyyzzz{{{{|||}}}~~~~����������������������������������������������������������������������������������������������������������������������������������� YZZZ[[[\\\\]]]^^^___````aaabbbcccddddeeefffggghhhhiiijjjkkkllllmmmnnnoooppppqqqrrrsssttttuuuvvvwwwxxxxyyyzzz{{{||||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� XXXYYYZZZ[[[\\\]]]^^^___````aaabbbcccdddeeefffggghhhhiiijjjkkklllmmmnnnoooppppqqqrrrssstttuuuvvvwwwxxxxyyyzzz{{{|||}}}~~~����������������������������������������������������������������������������������������������������������������������������������� VVWWWXXXYYYZZZ[[[\\\]]]^^^___```aaabbbcccdddeeefffggghhhiiijjjkkklllmmmnnnooopppqqqrrrssstttuuuvvvwwwxxxyyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� TUUUVVVWWWXXXYYZZZ[[[\\\]]]^^^___```aabbbcccdddeeefffggghhhiijjjkkklllmmmnnnooopppqqrrrssstttuuuvvvwwwxxxyyzzz{{{|||}}}~~~���������������������������������������������������������������������������������������������������������������������������������� RSSSTTTUUVVVWWWXXXYYZZZ[[[\\\]]^^^___```aabbbcccdddeefffggghhhiijjjkkklllmmnnnooopppqqrrrssstttuuvvvwwwxxxyyzzz{{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� PPQQRRRSSTTTUUUVVWWWXXXYYZZZ[[\\\]]]^^___```aabbbccdddeeeffggghhhiijjjkklllmmmnnooopppqqrrrsstttuuuvvwwwxxxyyzzz{{|||}}}~~���������������������������������������������������������������������������������������������������������������������������������� NNNOOPPPQQRRRSSTTTUUVVVWWXXXYYZZZ[[\\\]]^^^__```aabbbccdddeefffgghhhiijjjkklllmmnnnoopppqqrrrsstttuuvvvwwxxxyyzzz{{|||}}~~~���������������������������������������������������������������������������������������������������������������������������������� KKLLMMNNNOOPPPQQRRSSSTTUUVVVWWXXXYYZZ[[[\\]]^^^__```aabbcccddeefffgghhhiijjkkkllmmnnnoopppqqrrsssttuuvvvwwxxxyyzz{{{||}}~~~���������������������������������������������������������������������������������������������������������������������������������� HHIIJJKKLLLMMNNOOPPPQQRRSSTTTUUVVWWXXXYYZZ[[\\\]]^^__```aabbccdddeeffgghhhiijjkklllmmnnoopppqqrrsstttuuvvwwxxxyyzz{{|||}}~~���������������������������������������������������������������������������������������������������������������������������������� EEFFGGHHHIIJJKKLLMMNNOOPPPQQRRSSTTUUVVWWXXXYYZZ[[\\]]^^__```aabbccddeeffgghhhiijjkkllmmnnoopppqqrrssttuuvvwwxxxyyzz{{||}}~~���������������������������������������������������������������������������������������������������������������������������������� AABBCCDDEEFFGGHHIIJJKKLLMMNNOOPPQQRRSSTTUUVVWWXXYYZZ[[\\]]^^__``aabbccddeeffgghhiijjkkllmmnnooppqqrrssttuuvvwwxxyyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� ==>>??@@ABBCCDDEEFFGGHHIJJKKLLMMNNOOPPQRRSSTTUUVVWWXXYZZ[[\\]]^^__``abbccddeeffgghhijjkkllmmnnooppqrrssttuuvvwwxxyzz{{||}}~~��������������������������������������������������������������������������������������������������������������������������������� 889::;;<<=>>??@@ABBCCDDEFFGGHHIJJKKLLMNNOOPPQRRSSTTUVVWWXXYZZ[[\\]^^__``abbccddeffgghhijjkkllmnnooppqrrssttuvvwwxxyzz{{||}~~��������������������������������������������������������������������������������������������������������������������������������� 234455677889::;<<==>??@@ABBCDDEEFGGHHIJJKLLMMNOOPPQRRSTTUUVWWXXYZZ[\\]]^__``abbcddeefgghhijjkllmmnooppqrrsttuuvwwxxyzz{||}}~��������������������������������������������������������������������������������������������������������������������������������� ,,-../001223445667889::;<<=>>?@@ABBCDDEFFGHHIJJKLLMNNOPPQRRSTTUVVWXXYZZ[\\]^^_``abbcddeffghhijjkllmnnoppqrrsttuvvwxxyzz{||}~~��������������������������������������������������������������������������������������������������������������������������������� $%&&'(()*++,-../00123345667889:;;<=>>?@@ABCCDEFFGHHIJKKLMNNOPPQRSSTUVVWXXYZ[[\]^^_``abccdeffghhijkklmnnoppqrsstuvvwxxyz{{|}~~���������������������������������������������������������������������������������������������������������������������������������   !"#$$%&'(()*+,,-./0012344567889:;<<=>?@@ABCDDEFGHHIJKLLMNOPPQRSTTUVWXXYZ[\\]^_``abcddefghhijkllmnoppqrsttuvwxxyz{||}~���������������������������������������������������������������������������������������������������������������������������������   !"#$%&'(()*+,-./001234567889:;<=>?@@ABCDEFGHHIJKLMNOPPQRSTUVWXXYZ[\]^_``abcdefghhijklmnoppqrstuvwxxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������    Rr�!dS�Eb����CCᗵ|,��C�@E P(G�3s�>3�T0 k� �H�L14 'Q�1G�"H1 ��/    � 6 -Rr�!dW�Eb����DCᗵ|,��C�8E L(G�4s�>3�T0 k� �<�@14 'Q�1G�"H1 ��/    � 6 (Rr�!T[�Eb����ECᓵ|,��C�0E H'G�5s�=3�T0 k� �0�414 'Q�1G�"H1 ��/    � 6 #Rr�"T_�Eb����FCᓵ|,��C�(E D'G�6s�<3�T0 k� �$�(14 'Q�1G�"H1 ��/    � 6 Rr�"T_�Eb��	P�GCᓵ|,��C� E @&G�7s�<3�T0 k� ��14 'Q�1G�"H1 ��/    � 6 Rr�"Tc�Eb��	P�HCᏵ|,��C�E <&G�8c�;3�T0 k� ��14 'Q�1G�"H1 ��/    � 6 Rr�"Tg�Eb��	P�ICᏵ|,���C�E 8%G�8c�:3�T0 k� ��� 14 'Q�1G�"H1 ��/    � 6 Rr�"Tg�Eb��	P�JCድ|,���C�E 4$G�9c�:"s�T0 k� ����14 'Q�1G�"H1 ��/    � 6 
Rr�"�k�Eb��	P�KCድ|,���C� E 0$G�:c�9"s�T0 k� ����14 'Q�1G�"H1 ��/    � 6 Rr�#�k�Eb��	`�LCᇵ|,���C��E ,#G�;c�8"s�T0 k� ����14 'Q�1G�"H1 ��/    � 6 Rr�#�o�ER��	`�LC�|,��C��E (#G�;S�7"s�T0 k� ����14 'Q�1G�"H1 ��/    � 6��Rr�#�o�ER��	`�MC�|,��C��E $"G�<S�6"s�T0 k� ����14 'Q�1G�"H1 ��/    � 6��Rr�#�o�ER��	`�MC��|,��C��E  "G�=S�6"s�T0 k� ����14 'Q�1G�"H1 ��/    � 6��Rr�#�o�ER��	`�NC�{�|,��C��E !G�>S�5"s�T0 k� ����14 'Q�1G�"H1 ��/    � 6��Rr�#�o�ER����OC�w�|,�߉C��E !G�>S�4"s�T0 k� ����14 'Q�1G�"H1 ��/    � 6��Rr�$�o�ER����OE�s�|,�ۉC��E  G�?S�3"s�T0 k� ����14 'Q�1G�"H1  ��/    � 6��Rr�$�o�ER����PE�o�|,�׉C�E  G�@C�3"s�T0 k� ����14 'Q�1G�"H1  ��/    � 6��Rr�$�o�C�����QE�k�|,�ӉC�E G�@C�2"s�T0 k� �p�t14 'Q�1G�"H1  .�/    � 6��Rr�$�o�C�����RE�g�|,�ˊC�E G�AC�23�T0 k� �d�h14 'Q�1G�"H1  ��/    � 6��R��$�o�C�����RE�c�|,�ǊC�E C�BC�13�T0 k� �X�\14 'Q�1G�"H1  ��/    � 6��R��$�k�C�����SE�_�!�,�C�E C�BC�13�T0 k� �L�P14 'Q�1G�"H1  ��/    � 6��R��$�k�C�����TE�[�!�,�C�E  C�C��03�T0 k� �@�D14 'Q�1G�"H1  ��/    � 6��R��$�k�C�����UE�W�!�,�C�E/�C� D��03�T0 k� �(�,14 'Q�1G�"H1  ��(    � 6��R��%�g�C�����UE�S�!�,�D�E��C� D��/3�T0 k� �
�
14 'Q�1G�"H1  ��(    � 6��R��%�g�C�����VE�O�!�,�Dx E��C� E��/3�T0 k� ��14 'Q�1G�"H1  ��(    � 6��R��%�c�C�� ��WD1K�!�,�Dp E��EQ�E��/3�T0 k� ����14 'Q�1G�"H1  ��(    � 6��R��%�c�AR���WD1G�!�,�Dd!E��EQ�F��/3�T0 k� ����14 'Q�1G�"H1  ��(    � 6��R��%�_�AR���XD1C�!�,�D\!E��EQ�GC�/3�T0 k� ����14 'Q�1G�"H1  ��(    � 6��Ub�%�[�AR���YD1;�!�,��DT"E��EQ�GC�.3�T0 k� ����14 'Q�1G�"H1  ��(    � 6��Ub�%�W�AR���YD17�!�,��DL"E��EQ�HC�."��T0 k� ����14 'Q�1G�"H1  ��(    � 6��Ub�%�W�AR���ZD13�!�,��DD#E��EA�HC�."��T0 k� ����14 'Q�1G�"H1  ��(    � 6��Ub�&S�AR���[D1/�|,{�D<#E��EA�IC�."��T0 k� ����14 'Q�1G�"H1  ��(    � 6��Ub�&O�AR���[EQ'�|,s�D0$E��EA�I3�."��T0 k� ����14 'Q�1G�"H1  ��(    � 6��Ub�&K�AR���\EQ#�|,o�D($E��EA�I3�/"��T0 k� ����14 'Q�1G�"H1  ��(    � 6��Ub�&G�AR���]EQ�|,g�D %E��EA�J3�/"��T0 k� ����14 'Q�1G�"H1  ��(    � 6��Ub�&C�AR�	��]EQ�|,_�D%E��EA�J3�/"��T0 k� ����14 'Q�1G�"H1  ��(    � 6��Ub�&?�AR�
��^EQ�|,W�D%E��EA�J3�/"��T0 k� �� �� 14 'Q�1G�"H1  ��(    � 6��Ub�&;�AR���^EQ�|,O�D&E��E1�KC�0"��T0 k� ������14 'Q�1G�"H1  ��(    � 6��AR�&3�AR���_EQ�|,G�D�&E��E1�KC�0"��T0 k� ������14 'Q�1G�"H1  ��(    � 6��AR�&/�AR��`EP��|,?�D�'E��E1�KC�1"��T0 k� ������14 'Q�1G�"H1  ��(    � 6��AR�&+�AR��`EP��|,7�D�'EϼE1�KC�13�T0 k� ������14 'Q�1G�"H1  ��(    � 5��AR�''�AR��aEP�|,/�D�'E߸E1�KC�13�T0 k� ������14 'Q�1G�"H1  ��(    � 4��AR�'�AR��aC��!�,'�D�(Eߴ
E1�KC�13�T0 k� ����14 'Q�1G�"H1  ��(    � 3��C�'�AR��bC��!�,�E��(E߰	E1�JC�23�T0 k� ����14 'Q�1G�"H1  ��(    � 2��C�'�AR��bC�߿!�,�E��)E߬E!�JC�23�T0 k� ����14 'Q�1G�"H1  ��(    � 1��C�'�AR��cC�׿!�,�E��)EߤE!�JC|23�T0 k� ����14 'Q�1G�"H1  ��(    � 0��C�'�AR��cC���!�,�E�*EߠE!�JC|23�T0 k� ����14 'Q�1G�"H1  ��(    � /��C�'�AR� �dC���!�,��E�*EߜE!�JC|23�T0 k� �|��14 'Q�1G�"H1  ��(    � .��C�'��AR� �dC���!�,��E�+EߔE!�JC|23�T0 k� �x�|14 'Q�1G�"H1  ��(    � -��C�'��AR� �eC��!�,�E��+EߐE!�ISx23�T0 k� �p�t14 'Q�1G�"H1  ��(    � ,��C�'�AR� �eC��!�,��E��,E߈E!�ISx33�T0 k� �l�p14 'Q�1G�"H1  ��(    � +��C�'�AR� |fC��!�,�ۑE��,E߄E!�ISx33�T0 k� �d �h 14 'Q�1G�"H1  ��(    � *��C�(ߠAR� xfC��!�,�ӑE��-E�| E!�ISt33�T0 k� �`�d14 'Q�1G�"H1  ��(    � )��C�(�۠AR� pgC���|,�ˑD0|.E�{�E!�ISt33�T0 k� �X�\14 'Q�1G�"H1  ��(    � (��C�(�ӟAR� lgC��|,ῑD0t.E�s�E!�ISt33�T0 k� �P
�T
14 'Q�1G�"H1  ��(    � '��C�(�˟AR� dhC���|,᷒D0l/E�o�E!�ISt33�T0 k� �L�P14 'Q�1G�"H1  ��(    � &��C�|(�ßAR� \hC���|,ᯒD0d0E�g�E!�HSp33�T0 k� �D�H14 'Q�1G�"H1  ��(    � %��C�x(㻞AR� XhC��|,᧒D0\0A�c�E!�HSp43�T0 k� �<�@14 'Q�1G�"H1  ��(    � $��C�t(㳞AR�PiC�w�|,្D0P1A�[�E!�HSp43�T0 k� �0	�4	14 'Q�1G�"H1  ��( 
   � $��C�p(㫞AR�HiC�o�|,ᓒD0H2A�S�E!�HSp43�T0 k� �$�(14 'Q�1G�"H1  ��( 
   � #��C�l(㣝AR�DjC�g�|,ዒD0@3A�O�E!�Hcl43�T0 k� � �$14 'Q�1G�"H1  ��( 
   � #��C�d(㛝AR�<jC�_�|,გD083A�G�E!�Hcl43�T0 k� ��14 'Q�1G�"H1  ��( 
   � "��D`(㓝AR�4kC�W�|,�{�D004A�?�E!�Hcl43�T0 k� ��14 'Q�1G�"H1  ��( 
   � "��D\(㋜AR�,kC�O�|,�o�D0(5A�;�E!�Gcl43�T0 k� ��14 'Q�1G�"H1  ��( 
   � !��DX(ボAR�$kC�G�|,�g�D0 6A�3�E!�Gcl43�T0 k� ��14 'Q�1G�"H1  ��( 
   � !��DP)�{�AR�lD C�|,�_�D@7A�+�E!�Gch53�T0 k� ����14 'Q�1G�"H1  ��( 
   � !��DL)�s�AR�lD ;�|,�W�D@7A�'�E!�Gch53�T0 k� ����14 'Q�1G�"H1  ��( 
   � !��DH)�k�AR�lD 3�|,�O�D@8A��E!�Gch53�T0 k� ����14 'Q�1G�"H1  ��( 
   �  ��D@)�c�AR�mD +�|,�C�D@ 9A��E!�Gch53�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �D<)�[�AR�� mD #�|,�;�DO�:A��E!�Gch53�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �}D4)�S�AR���mD �|,�3�DO�;A��E!�Gcd53�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �{D0)�K�AR���nD �|,�+�DO�<A��E!�Fsd53�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �yD()�C�AR���nD �|,�#�DO�=A���E!�Fsd53�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �wD$)�;�AR���oD �|,�DO�>A���E!�Fsd53�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �uD)�3�AR���oD��|,�DO�?A���E!�Fsd63�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �sD)�+�AR���oD��|,�DO�@A���E!|Fs`63�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �qD)#�AR���pD��|, ��D_�AA���E!|Fs`63�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �oD)�A����pD��|, �D_�AA���E!|Fs`63�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �mD )�A���pD��|, �D_�BA���E!xFs`63�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �kD�)�A��߰pD��|, �D_�CA���E!xFs`63�T0 k� ����14 'Q�1G�"H1  ��( 
   �  �iD�)�A��ߨqD��|, ەD_�DA޿�E!tEs\63�T0 k� ��	��	14 'Q�1G�"H1  ��( 
   �  �gD�*��A��ߠqD��|, ӕI��EA޷�E!tEs\63�T0 k� �x	�|	14 'Q�1G�"H1  ��( 
   �  �eD�*�A�ߘqD��|, ǕI��FAޯ�E!tE\63�T0 k� �p	�t	14 'Q�1G�"H1  ��( 
   �  �cD�*�A�ߐrD��|, ��I��GAާ�E!pE\73�T0 k� �h
�l
14 'Q�1G�"H1  ��X 	   �  �aC��*�A�߈rD��|,��I��GAޟ�E!pE\73�T0 k� �`
�d
14 'Q�1G�"H1  �X 	   �  �_C��*ۖA�߀rD��|,��I�|HAޗ�E!lDX73�T0 k� �X�\14 'Q�1G�"H1  ��X 	   �  �]C��*ӖA��xrD��|0��I�xIAޏ�E�lDX73�T0 k� �P�T14 'Q�1G�"H1  ��X 	   �  �[C�*˖A��psC��|0��I�tIA��E�lD�X83�T0 k� �H�L14 'Q�1G�"H1  ��X 	   �  �YC�*ÖA��hsC��|0��I�lJA��E�hC�T83�T0 k� �@�D14 'Q�1G�"H1  ��X 	   �  �WC�*��A���`sC��|4��I�hJA�w�E�hC�T83�T0 k� �8�<14 'Q�1G�"H1  ��X 	   �  �UC�*��A���XsC��|8��I�dJA�l E�dB�P83�T0 k� �0�414 'Q�1G�"H1  ��X 	   �  �SC�*��A���PsC�{�|8w�E_\KA�d E�dB�L93�T0 k� �(�,14 'Q�1G�"H1  ��X 	   �  �QC�*��A���HtC�s�|<o�E_XKA�\E�`A�L93�T0 k� � �$14 'Q�1G�"H1  ��X 	   �  �OC�*��A��?DtC�k�|@g�E_TLA�TE�`A�H93�T0 k� ��14 'Q�1G�"H1  ��X 	   �  �MC�*��A��?<tC�c�|D_�E_LLA�LE�\@�D93�T0 k� ��14 'Q�1G�"H1  ��X 	   �  �KC�x*��AR�?4tC�[�|H�W�E_HLA�DE�\?�@:3�T0 k� ��14 'Q�1G�"H1  ��X 	   �  �IC�p*��AR�?,tC�S�|L�K�E_@MA�<C�X?�@:3�T0 k� � �14 'Q�1G�"H1  ��X 	   �  �GC�h*�AR�?$tC�K�|P�C�E_<MA�4C�T>�<:3�T0 k� ����14 'Q�1G�"H1  ��X 	   �  �FC�\*�w�AR�?tC�C� |T�;�E_4MA�,C�T=�8:3�T0 k� ����14 'Q�1G�"H1  ��X 	   �  �EC�T*�o�AR�?sC�;� |X�3�E_0NA�(C�P=�4;3�T0 k� ����14 'Q�1G�"H1  ��X 	   �  �DC�L*�g�C�?sC�3� |\�'�E_(NA� C�L<�0;3�T0 k� ����14 'Q�1G�"H1  ��X 	   �  �CC�D+�_�C�OsC�+� |`��C� OA�C�H;�,;3�T0 k� ����14 'Q�1G�"H1  ��X 	   �  �BC�<+�W�C�N�sC�#� |d��C�OA�C�H;�$;3�T0 k� ����14 'Q�1G�"H1  ��X 	   �  �AC�(*�G�C�N�rC�� |l��C�PA� 
C�@:�<3�T0 k� ����14 'Q�1G�"H1  ��X    �  �@C� *�?�C�N�rC�� |p���C�PA��C�<:�<3�T0 k� ����14 'Q�1G�"H1  ��X    �  �?C�*�7�C�N�rC�� |t��C��PE]�C�89�<3�T0 k� ����14 'Q�1G�"H1  ��X    �  �>D)�/�C�N�rC��� |x��C��PE]�C�48�<3�T0 k� ����14 'Q�1G�"H1  ��X    �  �=D)�'�C�N�qC��� �|��C��QE]�C�08�=3�T0 k� ����14 'Q�1G�"H1  ��X    �  �<D )��C�N�qC��� ���ۗC��QE]�C�,7� =3�T0 k� ����14 'Q�1G�"H1  ��X    �  �;D �)��C�N�qD�� ���ϘC��QE]�C�(6��=3�T0 k� ��	��	14 'Q�1G�"H1  ��X    �  �:D �(��C�N�pD�� ���ǘC��RE]�C�$5��=3�T0 k� ��	��	14 'Q�1G�"H1  ��X    �  �9D �(��C�^�pD�� �����C��RE]�C� 5��=3�T0 k� ��	��	14 'Q�1G�"H1  ��X    �  �8D �(���C�^�pD�� �����C��RE]�C�4��>3�T0 k� ��	��	14 'Q�1G�"H1  ��X    �  �8D �(���C�|^�oD�� �����C��SE]�C�3��>3�T0 k� ����14 'Q�1G�"H1  ��X    �  �8D �(��C�x^�oE�� �����C��SE]�C�2��>3�T0 k� ��	��	14 'Q�1G�"H1  ��X    �  �8D �'��C�t^�nE�� �����C��SE]�C�1��>3�T0 k� ��
��
14 'Q�1G�"H1  ��X    �  �8D �'�ߑC�p^�nE�� �����C��SE]�C�0��>3�T0 k� �x
�|
14 'Q�1G�"H1  �X    �  �8D�'QϑC�d^xmE�� ��_�A^�TE]�C��/R�?3�T0 k� �h�l14 'Q�1G�"H1  �X    �  �8D�'QǑD`^plE�� ��_w�A^�TE]�C��.R�?3�T0 k� �`�d14 'Q�1G�"H1  ��X    �  �8D�&Q��DX^hlE�� ��_o�A^|TE]|A �-R�?3�T0 k� �X�\14 'Q�1G�"H1  ��X    �  �8D�&Q��DT^`kE�� ��_g�A^tUE]tA �,R�?3�T0 k� �P�T14 'Q�1G�"H1  ��X    �  �8D�&Q��DP^XkE�� ��__�A^lUEMlA �+R�?3�T0 k� �H�L14 'Q�1G�"H1  ��X    �  �8D�&Q��DH^PjE�{� ��_W�A^dUEMdA �*R�@3�T0 k� �@
�D
14 'Q�1G�"H1  ��X    �  �8Dx&Q��D@^HjD>s� ��_O�A^\UEM\A �*R�@3�T0 k� �8	�<	14 'Q�1G�"H1  ��X    �  �8Dl%Q��M<^@iD>k� ��_G�A^TVEMTA �)R�@3�T0 k� �0�414 'Q�1G�"H1  ��X    �  �8Dd%Q��M4^8iD>c� ��_?�A^LVEMLA �(R�@3�T0 k� �(�,14 'Q�1G�"H1  ��X    �  �8D\%Q��M0^0iD>[� ��_7�A^DVEMDA �'R�@3�T0 k� � �$14 'Q�1G�"H1  ��X   �  �8C�T%A�M(�(hD>W� ��_3�A^@VEM<A �&R�@3�T0 k� ��14 'Q�1G�"H1  ��X    �  �8C�L%Aw�M$�$hD>O� ��_+�A^8WEM4A �&R�A3�T0 k� ��14 'Q�1G�"H1  ��X    �  �8C�D%Ao�M �gD>G� ��_#�A^0WEM,A �%RxA3�T0 k� ��14 'Q�1G�"H1  ��X    �  �8C�<$Ag�M�gD>?� ��_�A^(WEM$A �$RtA3�T0 k� � �14 'Q�1G�"H1  ��X    �  �8C�0$A_�M�fD>7� ��_�A^(WEMA �$RpA3�T0 k� ����14 'Q�1G�"H1  $�X    �  �8C�($AW�M�fD>/� ��_�A^$WEMA �#RhA3�T0 k� <�	� 	14 'Q�1G�"H1  ��_    �  �8C� $AO�M��fD>'� ��_�A^WE�A �"RdA3�T0 k� = 	�	14 'Q�1G�"H1  ��_    �  �8C�$AG�M"��fD>� ��^��A^WE� A �!R`A3�T0 k� =	�	14 'Q�1G�"H1  ��_    �  �8C�$A?�M" ��fL>� ��^��A^WE��A �!R\B3�T0 k� =
�
14 'Q�1G�"H1  ��_    �  �8C�#A7�M!���fL>� ��^�A^WE��A � RTB3�T0 k� =
�
14 'Q�1G�"H1  ��_    �  �8C� #�/�M!���fL>� ��^�A^WE��A �RPB3�T0 k� ��14 'Q�1G�"H1  ��_    �  �8C��#�'�M!���eL>� ��^�A]�WE��A �RLB3�T0 k� ��14 'Q�1G�"H1  ��_    �  �8C��#��M!���eL=�� ��^ߙA]�WE��A �RHB3�T0 k� ��14 'Q�1G�"H1  ��_    �  �8C��#��M!���eL=�� ��^ۙA]�WE��A �RDB3�T0 k� ��14 'Q�1G�"H1  ��_    �  �8C��#��M!���eL=�� ��^әA]�WE��A �R<B3�T0 k� ��14 'Q�1G�"H1  ��_    �  �8C��#��M!���eL=�� ��^ϚA]�WE��A �R8C3�T0 k� �� 14 'Q�1G�"H1  ��_   �  �8C��"���M���eL=�� ��^˚A]�WEܸA �R4C3�T0 k� � �$14 'Q�1G�"H1  ��_    �  �8C��"���M���eL=�� ��^ÚA]�WEܰA �R0C3�T0 k� �$�(14 'Q�1G�"H1  ��_    �  �8C��"��M���dL=�� ��^��A]�WEܤA �R,C3�T0 k� �(�,14 'Q�1G�"H1  ��_    �  �8L�"��M���dL=�� ��^��A]�WEܜA �R(C3�T0 k� �(�,14 'Q�1G�"H1  ��_    �  �8L�"�ߔM���dL=�� ��^��A]�WEܔA �R$C3�T0 k� �,�014 'Q�1G�"H1  ��_    �  �8L�"�הM���dL=�� ��^��A]�WC܈A �R C3�T0 k� �0�414 'Q�1G�"H1  ��_    �  �8L�"�ϕM��|dLM�� ��^��A]�WC�xA �RC3�T0 k� �4�814 'Q�1G�"H1  ��_    �  �8L�"�ǕM�tdLM�� ��^��A]�WC�hA �RC3�T0 k� �4�814 'Q�1G�"H1  ��_    �  �8L�"���M�ldLM�� ��^��A]�WC�\A �RD3�T0 k� �8�<14 'Q�1G�"H1  ��_    �  �8L�!���C�ddLM�� ��^��A]�WC�PA �RD3�T0 k� �<�@14 'Q�1G�"H1  ��_    �  �8Lx!���C�`dLM�� ��^��A]�WC�@A |RD3�T0 k� �@�D14 'Q�1G�"H1  ��_    �  �8Lp!���C�XdLM�� ��^��A]�WC�4A xRD3�T0 k� �D�H14 'Q�1G�"H1  ��_    �  �8Ll!���C�	�PdLM�� |�^��A]�VC�(A xRD3�T0 k� �D�H14 'Q�1G�"H1  ��_    �  �8Ld!�C�	�HdLM�� |�^��A]�VC�A tR D3�T0 k� �H�L14 'Q�1G�"H1  ��_    �  �8L\!�C�	�DdLM�� } ^��A]�VC�A tQ�D3�T0 k� �L�P14 'Q�1G�"H1  ��_    �  �8LT!���C�	�<dLM�� } ^{�A]�VC�A pQ�D3�T0 k� �P�T14 'Q�1G�"H1  ��_    �  �8LL!���C�	�8dLM�� } ^w�A]�VC��A lQ�D3�T0 k� �P�T14 'Q�1G�"H1  ��_   �  �8L/H!�{�C�	�4dLM�� }^s�A]�VC��A lQ�D3�T0 k� �T�X14 'Q�1G�"H1  ��_    �  �8L/@ �s�C�	�,dLM� }^o�A]�VC��A hQ�E3�T0 k� �X�\14 'Q�1G�"H1  ��_    �  �8L/8 �o�C�|	�(dLM{� }^k�A]�VC��A hQ�E3�T0 k� �\�`14 'Q�1G�"H1  ��_    �  �8L/4 �g�C�x	�$dLMw� }^g�A]�VC��A dQ�E3�T0 k� �\�`14 'Q�1G�"H1  ��_    �  �8L/, �_�C�p	� dLMo� }^c�A]�VC��A `Q�E3�T0 k� �`�d14 'Q�1G�"H1  ��_    �  �8L/( �[�C�l	�dLMk�}^_�A]|VCۼA `Q�E3�T0 k� �d�h14 'Q�1G�"H1  ��_    �  �8L/  �S�C�d	�dLMg�}^[�A]xVC۰A \Q�E3�T0 k� �h�l14 'Q�1G�"H1  ��_    �  �8L/ �K�C�\	�dLMc�}^W�A]tVCۨA \Q�E3�T0 k� �h�l14 'Q�1G�"H1  ��_    �  �8L/ �G�C�X	�dLM_�}^S�A]pVCۜ A XQ�E3�T0 k� �l�p14 'Q�1G�"H1  ��_    �  �8L/ �?�C�P	�dLM[�}^O�A]lVC۔!A XQ�E3�T0 k� �p�t14 'Q�1G�"H1  ��_    �  �8L/  ;�C�H	�dLMW�}^K�A]hVCی!A TQ�E3�T0 k� �t�x14 'Q�1G�"H1  ��_    �  �8L/  3�C�@	�dLMS�}^G�A]dVCی"A TQ�E3�T0 k� �x�|14 'Q�1G�"H1  ��_    �  �8L.�  /�C�8	� dLMO�}^C�A]`VCې#A PQ�F3�T0 k� �x�|14 'Q�1G�"H1  ��_    �  �8L.� '�C�0	� dLMK�}^?�A]\VCې$A PQ�F3�T0 k� �|��14 'Q�1G�"H1  ��_    �  �8L.� #�C�,	��dLMG�}^?�A]\VA[�$A LQ�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.� �D$�dLMC�}^;�A]XVA[�%A LQ�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.� �D�dLM?�}^7�A]TVA[�&A HQ�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.� �D�dLM;�}^3�A]PVA[�&A HQ�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.� �D�dLM7�}^/�A]LVA[�'A DQ�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.� �D �dLM3�}^+�A]LVA[�(A DQ�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.� �D ��dLM/�}^+�A]HVA[�(A DQ�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.���D ��dLM+�}^'�A]DVA[�)A @Q�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.���D ��dLM+�}^#�A]@VA[�)A @Q�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.��D ��dLM'�}^�A]@VA[�*A <Q�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.��D ��dLM#�}^�A]<VA[�+A <
Q�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.��D ��dLM�}^�A]8VA[�+A 8
Q�F3�T0 k� ����14 'Q�1G�"H1  ��_    �  �8L.��D��dLM�}^�A]4VA[�,A 8
Q�G3�T0 k� �� �� 14 'Q�1G�"H1  ��_    �  �8L.�ߧD��dLM�}^�A]4VA[�,A 8	Q�G3�T0 k� �� �� 14 'Q�1G�"H1  ��_    �  �8L.�ۧD�,�dLM�}^�A]0VA[�-A 4	Q�G3�T0 k� �� �� 14 'Q�1G�"H1  ��_    �  �8L.�רD�,�dLM�}^�A],VA[�-A 4	Q�G3�T0 k� ��!��!14 'Q�1G�"H1  ��_    �  �8L.�ӨD�,�dL=�}^�A],VA[�.A 4Q�G3�T0 k� ��!��!14 'Q�1G�"H1  ��_    �  �8L.�ϨD�,�dL=�}^�A](VA[�.A 0Q�G3�T0 k� ��"��"14 'Q�1G�"H1  ��_    �  �8L.�˩D�,�dL=�}^�A]$VA[�/A 0Q�G3�T0 k� ��"��"14 'Q�1G�"H1  ��_    �  �8L.�éD�,�dL=�}^�A]$VA[�/A 0Q�G3�T0 k� ��#��#14 'Q�1G�"H1  ��_    �  �8L.���Dx,�dL=�}^�A] VA[�0A ,Q�G3�T0 k� ��#��#14 'Q�1G�"H1  ��_    �  �8L.���Dl,�dL<��}]��A] VA[�0A ,Q�G3�T0 k� ��#��#14 'Q�1G�"H1  ��_    �  �8L.���Dd,�dD<��}]��A]VA[�1A (Q�G3�T0 k� ��$��$14 'Q�1G�"H1  ��_    �  �8L.���C�X,�dD<��}]��A]VA[�1A (Q�G3�T0 k� ��$��$14 'Q�1G�"H1  ��_    �  �8L.���C�P,�dD<��}]��A]VA[�2A (Q�G3�T0 k� ��%��%14 'Q�1G�"H1  ��_    �  �8L.���C�H,�dD<��}]��A]VA[�2A $Q�G3�T0 k� ��%��%14 'Q�1G�"H1  ��_    �  �8L.���C�<,�dD<��}]�A]VA[�3A $Q�G3�T0 k� ��%��%14 'Q�1G�"H1  ��_    �  �8L|��C�4,�dE���}]�A]VA[�3A $Q�G3�T0 k� ��&��&14 'Q�1G�"H1  ��_    �  �8Lx��C�(,�dE���}]�A]VA[�4A $Q�G3�T0 k� ��&��&14 'Q�1G�"H1  ��_    �  �8Lt��C� ,�dE���}]�A]VA[�4A  Q�H3�T0 k� ��'��'14 'Q�1G�"H1  ��_   �  �8Lp��C�,�dE���}]�A]VA[�4A  Q�H3�T0 k� ��'��'14 'Q�1G�"H1  ��_    �  �8Ll��C�,�dE���}]�A]VA[�5A  Q�H3�T0 k� ��'��'14 'Q�1G�"H1  ��_    �  �8Ll��C�,�dE���}]�A]VA[�5A Q�H3�T0 k� ��(��(14 'Q�1G�"H1  ��_    �  �8C�h��M�,�dE���}]�A]VA[�6A Q�H3�T0 k� ��(��(14 'Q�1G�"H1  ��_    �  �8C�d��M�,�dE���}]�A]VA[�6A Q�H3�T0 k� ��(��(14 'Q�1G�"H1  ��_    �  �8C�`��M�,�dE���}]ߜA] VA[�6A Q�H3�T0 k� ��)��)14 'Q�1G�"H1  ��_    �  �8C�\��M�,�dE���}]ߜA] VA[�7A Q�H3�T0 k� ��)��)14 'Q�1G�"H1  ��_    �  �8C�X���M�,�dE���}]ۜA\�VA[�7A Q�H3�T0 k� ��*��*14 'Q�1G�"H1  ��_    �  �8C�T��M�,�dE���}]ۜA\�VA[�8A Q|H3�T0 k� ��*��*14 'Q�1G�"H1  ��_    �  �8E�P�{�M�,�dD���}]לA\�VA[�8A Q|H3�T0 k� ��*��*14 'Q�1G�"H1  ��_    �  �8E�H�{�M�,�dD���}]לA\�VA[�8A Q|H3�T0 k� ��+��+14 'Q�1G�"H1  ��_    �  �8E�D�w�M�,�dD���}]ӜA\�VA[�9A QxH3�T0 k� ��+��+14 'Q�1G�"H1  ��_    �  �8E�@�s�M�,�dD���}]ӜA\�VA[�9A QxH3�T0 k� ��,��,14 'Q�1G�"H1  ��_    �  �8E�<�o�M/�,�dD���}]ϜA\�VA[�9A QtH3�T0 k� ��,� ,14 'Q�1G�"H1  ��_    �  �8E�8�o�M/�,�dD���}]ϜA\�VA[�:A QtH3�T0 k� �.�.14 'Q�1G�"H1  ��     �  �8E�0�k�M/�,�dD����]˜A\�VA[�:A QtH3�T0 k� �0�014 'Q�1G�"H1  ��     �  �8E�,�g�M/�,�dD���]˜A\�VA[�:A QtH3�T0 k� �1�114 'Q�1G�"H1  ��     �  �8E�(�c�M/�,�dD���]˜A\�VA[�;A QpH3�T0 k� �1�114 'Q�1G�"H1  ��     �  �8E�$�_�M/x,�dD���]ǜA\�VA[�;A QpH3�T0 k� � 2�214 'Q�1G�"H1  ��     �  �8A� �[�M/p,�dD���]ǜA\�VA[�;A QpH3�T0 k� ��/� /14 'Q�1G�"H1  ��     �  �8A��W�M/l,�dD��}]ÜA\�VA[�<A QlH3�T0 k� ��-��-14 'Q�1G�"H1  ��     �  �8A��S�M/d,�dD��}]ÜA\�VA[�<A QlI3�T0 k� ��+��+14 'Q�1G�"H1  ��     �  �8A��O�M\,�dD��}]ÜA\�VA[�<A QlI3�T0 k� ��*��*14 'Q�1G�"H1  ��    �  �8A� �K�MT,�dD��
} ]��A\�VA[�=A QhI3�T0 k� ��)��)14 'Q�1G�"H1  ��     �  �8A� �G�ML,�dD��} ]��A\�VA[�=A QhI3�T0 k� ��(��(14 'Q�1G�"H1  ��     �  �8A� �C�MH�dD��|�]��A\�VA[�=A QhI3�T0 k� ��(��(14 'Q�1G�"H1  ��     �  �8A�  �?�M@�dD��|�]��A\�VA[�>A  QhI3�T0 k� ��(��(14 'Q�1G�"H1  ��     �  �8A�� �;�M8�dD����]��A\�VA[�>A  QdI3�T0 k� ��(��(14 'Q�1G�"H1  ��     �  �8A�� �3�M4�dD����]��A\�VA[�>A  QdI3�T0 k� ��(��(14 'Q�1G�"H1  ��     �  �8A��!�/�M,�dD�|��]��A\�VA[�>A  QdI3�T0 k� ��(��(14 'Q�1G�"H1  ��     �  �8A��!�+�M(�dD�|��]��A\�VA[�?A  Q`I3�T0 k� ��(��(14 'Q�1G�"H1  ��     �  �8A��!�'�C� �dD�x��]��A\�VA[�?A  Q`I3�T0 k� ��(��(14 'Q�1G�"H1  ��     �  �8A��!��C��dD�t��]��A\�VA[�?A  Q`I3�T0 k� ��)��)14 'Q�1G�"H1  ��     �  �8A��!��C��dD�t��]��A\�VA[�?A   Q`I3�T0 k� ��)��)14 'Q�1G�"H1  ��     �  �8A��!��C��dD�p��]��A\�VA[�@A �Q`I3�T0 k� ��)��)14 'Q�1G�"H1  ��     �  �8A��"��C��dE�p��]��A\�VA[�@A �Q\I3�T0 k� ��)��)14 'Q�1G�"H1  ��     �  �8A��"��C���dE�l��]��A\�VA[�@A �Q\I3�T0 k� ��)��)14 'Q�1G�"H1  ��     �  �8A��"��C���dE�h!��]��A\�VA[�@A �Q\I3�T0 k� ��)��)14 'Q�1G�"H1  ��     �  �8A��"���C����dE�h#��]��A\�VA[�AA �Q\I3�T0 k� ��*��*14 'Q�1G�"H1  ��     �  �8A��"���C����dE�d%��]��A\�VA[�AA��QXI3�T0 k� ��*��*14 'Q�1G�"H1  ��     �  �8A��"���E����dE�d&��]��A\�VA[�AA��QXI3�T0 k� ��*��*14 'Q�1G�"H1  ��     �  �8A��"���E����dE�`(��]��A\�VA[�AA��QXI3�T0 k� ��*��*14 'Q�1G�"H1  ��     �  �8A��#���E����dE�`*��]��A\�VA[�BA��QXI3�T0 k� ��*��*14 'Q�1G�"H1  ��     �  �8A��#���E����dL\\,<�]��A\�VA[�BA��QTI3�T0 k� ��*��*14 'Q�1G�"H1  ��     �  �8A��#���E����dL\X.<�]��A\�VA[�BA��QTI3�T0 k� ��*��*14 'Q�1G�"H1  ��     �  �8A��#���M���dL\X0<�]��A\�VA[�BA��QTI3�T0 k� ��*��*14 'Q�1G�"H1  ��     �  �8A��#���M���cL\T1<�]��A\�VA[�BA��QTI3�T0 k� ��+��+14 'Q�1G�"H1  ��     �  �8A��#���M���cL\T3<�]��A\�VA[�CA��QTI3�T0 k� ��+��+14 'Q�1G�"H1  ��     �  �8A��#���M�ܔcL\P5<�]��A\�VA[�CA��QTI3�T0 k� ��+��+14 'Q�1G�"H1  ��     �  �8A��#λ�M�ܘcL\P6<�]��A\�VA[�CA��QPI3�T0 k� ��+��+14 'Q�1G�"H1  ��     �  �8A��$η�M�ܘcL\L8<�]��A\�VA[�CA��QPI3�T0 k� ��+��+14 'Q�1G�"H1  ��     �  �8A��$ί�M.�ܘcL\L:<�]��A\�VA[�CA��QPJ3�T0 k� ��+��+14 'Q�1G�"H1  ��     �  �8A��$Ϋ�M.�ܘcL\L;<�]��A\�UA[�DA��QPJ3�T0 k� ��+��+14 'Q�1G�"H1  ��     �  �8A��$Σ�M.�ܘcL\H=<�]��A\�UA[�DA��QPJ3�T0 k� ��+��+14 'Q�1G�"H1  ��     �  �8A��$Λ�M.�ܜcL\H><�]��A\�UA[�DA��QLJ3�T0 k� ��,��,14 'Q�1G�"H1  ��     �  �8A��$Η�M.xܜcL\D@<�]��A\�UA[�DA��QLJ3�T0 k� ��,��,14 'Q�1G�"H1  ��     �  �8A��$Ώ�M.tܜcL\DA<�]��A\�UA[�DA��QLJ3�T0 k� �|,��,14 'Q�1G�"H1  ��     �  �8A��$΃�M.hL�cLl@D<�]��A\�TA[�EA��QLJ3�T0 k� �x,�|,14 'Q�1G�"H1  ��     �  �8A��%��M.`L�cLl<F<�]��A\�TA[�EA��QLJ3�T0 k� �t,�x,14 'Q�1G�"H1  ��     �  �8A��%�w�M\L�cLl<G<�]��A\�SA[�EA��QHJ3�T0 k� �t,�x,14 'Q�1G�"H1  ��     �  �8A��%�s�MXL�cLl<I<�]��A\�SA[�EA��QHJ3�T0 k� �p,�t,14 'Q�1G�"H1  ��     �  �8A��%�k�MPL�bLl<I<�]��A\�SA[�EA��QHJ3�T0 k� �p,�t,14 'Q�1G�"H1  ��     �  �8A��%�g�ML��bLl<J<�]��A\�RA[�FA��QHJ3�T0 k� �l-�p-14 'Q�1G�"H1  ��     �  �8A��%�_�MD��bLl<L<�]��A\�RA[�FA��QHJ3�T0 k� �h-�l-14 'Q�1G�"H1  ��     �  �8A��%�[�M@��aLl8M<�]��A\�RA[�FA��QHJ3�T0 k� �h-�l-14 'Q�1G�"H1  ��     �  �8A��%�S�M<��aLl8N<�]��A\�RA[�FA��QHJ3�T0 k� �d-�h-14 'Q�1G�"H1  ��     �  �8A��%�O�M8��aLl8P<�]��A\�QA\ FA��QDJ3�T0 k� �d-�h-14 'Q�1G�"H1  ��     �  �8A��%�G�M0��aLl4Q<|]��A\�QA\ FA��QDJ3�T0 k� �`-�d-14 'Q�1G�"H1  ��     �  �8A��&�C�E�,��`Ll4R<|]��A\�QA\ FA��QDJ3�T0 k� �`-�d-14 'Q�1G�"H1  ��     �  �8A��&�;�E�(��`Ll4S<|]��A\�PA\ GA��QDJ3�T0 k� �\-�`-14 'Q�1G�"H1  ��     �  �8A��&�7�E� ��`Ll0U<x]��A\�PA\ GA��QDJ3�T0 k� �\-�`-14 'Q�1G�"H1  ��     �  �8A�|&�/�E���`Ll0V<x]��A\�PA\ GA��QDJ3�T0 k� �X-�\-14 'Q�1G�"H1  ��     �  �8A�|&�+�E���`Ll0W<x]��A\�PA\ GA��QDJ3�T0 k� �X-�\-14 'Q�1G�"H1  ��    �  �8A�x&�#�E���`Ll0X<t]��A\�OA\ GA��Q@J3�T0 k� �T.�X.14 'Q�1G�"H1  ��     �  �8A�x&��E���`Ll,Y<t]��A\�OA\ GA��Q@J"��T0 k� �T.�X.14 'Q�1G�"H1  ��    �  �8A�t&��E� ��`Ll,Z<t]��A\�OA\ GA��Q@J"��T0 k� �P.�T.14 'Q�1G�"H1  ��     �  �8A�t&��E�  ��`Ll,[<p]��A\�OA\ GA��Q@J"��T0 k� �P.�T.14 'Q�1G�"H1  ��     �  �8A�p&��E�� ��`Ll,\<p]��A\�NA\ HA��Q@J"��T0 k� �L.�P.14 'Q�1G�"H1  ��     �  �8A�p&��D=�!��`Ll(]<p]��A\�NA\ HA��Q@J"��T0 k� �L.�P.14 'Q�1G�"H1  ��     �  �8A�l&��D=�!��`Ll(_<l]��A\�NA\ HA��Q@J"��T0 k� �H.�L.14 'Q�1G�"H1  ��     �  �8A�l'���D=�"��`Ll(`<l]��A\�NA\ HA��Q@J"��T0 k� �H.�L.14 'Q�1G�"H1  ��     �  �8A�l'���D=�"��`Ll(a<l]��A\�MA\ HA��Q<J"��T0 k� �H.�L.14 'Q�1G�"H1  ��     �  �8A�h'���D=�# �`Ll$b<h]��A\�MA\HA��Q<J"��T0 k� �D.�H.14 'Q�1G�"H1  ��     �  �8A�h'��D=�$ �`Ll$c<h]��A\�MA\HA��Q<J"��T0 k� �D.�H.14 'Q�1G�"H1  ��     �  �8A�d'��D=�$ �`Ll$c<h]��A\�MA\HA��Q<J"��T0 k� �@.�D.14 'Q�1G�"H1  ��    �  �8A�d'��D=�% �`Ll$d<d]��A\�MA\HA��Q<J3�T0 k� �@/�D/14 'Q�1G�"H1  ��     �  �8A�d'��D=�& �`Ll e<d]��A\�LA\HA��Q<J3�T0 k� �@/�D/14 'Q�1G�"H1  ��     �  �8A�`'��D=�' �`Ll f<d]��A\�LA\IA��Q<J3�T0 k� �</�@/14 'Q�1G�"H1  ��     �  �8A�`'��D=�' �`Ll g<d]��A\�LA\IA��Q<J3�T0 k� �</�@/14 'Q�1G�"H1  ��     �  �8A�\'� D=�( �`Ll h<`]��A\�LA\IA��Q<J3�T0 k� �8/�</14 'Q�1G�"H1  ��     �  �8A�\'�DM�) �`Ll i<`]��A\�LA\IA��Q<J3�T0 k� �8/�</14 'Q�1G�"H1  ��     �  �8A�\'�DM�* �`Llj<`]��A\�KA\IA��Q8J3�T0 k� �8/�</14 'Q�1G�"H1  ��     �  �8A�X'�DM�*L�`Llk<\]��A\�KA\IA��Q8K3�T0 k� �4/�8/14 'Q�1G�"H1  ��     �  �8A�T'�DM�+L�`Llk<\]�A\�KA\IA��Q8K3�T0 k� �0/�4/14 'Q�1G�"H1  ��     �  �8A�T'�DM�,L�`Lll<\]�A\�KA\IA��Q8K3�T0 k� �0/�4/14 'Q�1G�"H1  ��     �  �8A�P'�DM�-L�`Llm<\]�A\�KA\IA��Q8K3�T0 k� �,/�0/14 'Q�1G�"H1  ��     �  �8A�L'�DM�.L�`Lln<X]�A\�JA\IA��Q8K"s�T0 k� �(/�,/14 'Q�1G�"H1  ��     �  �8A�H'�DM�0L�`L\o<X]�A\�JA\JA��Q8K"s�T0 k� �$/�(/14 'Q�1G�"H1  ��     �  �8A�D'�DM�1L�`L\o<X]�A\�JA\JA��Q8K"s�T0 k� � /�$/14 'Q�1G�"H1  ��     �  �8A�@'�	DM|2L�`L\p<X]�A\�JA\JA��Q8K"s�T0 k� �.� .14 'Q�1G�"H1  ��     �  �8A�@'�
DMt3L�`L\q<X]�A\�JA\JA��Q8K"s�T0 k� �.� .14 'Q�1G�"H1  ��     �  �8A�<'�D]p5L�`L\r<T]�A\�JA\JA��Q8K"s�T0 k� �.�.14 'Q�1G�"H1  ��     �  �8A�8'�D]h6L�`L\r<T]{�A\�IA\JA��Q8K"s�T0 k� �.�.14 'Q�1G�"H1  ��     �  �8A�4'�D]d7L�`Fs<T]{�A\�IA\JA��Q4K"s�T0 k� �.�.14 'Q�1G�"H1  ��     �  �8A�4'�D]`9��`Ft<T]{�A\�IA\JA��Q4K"s�T0 k� �.�.14 'Q�1G�"H1  ��     �  �8A�0&�D]X:��`Fu<P]{�A\�IA\JA��Q4K"s�T0 k� �.�.14 'Q�1G�"H1  ��     �  �8A�,&�D]T;��`Fv<P]{�A\�IA\JA��Q4K"s�T0 k� �.�.14 'Q�1G�"H1  ��     �  �8A�(&�D]L=��`Fv<P]{�A\�IA\JA��Q4K3�T0 k� �.�.14 'Q�1G�"H1  ��     �  �8A�(&�D]H>��`Fw<P]{�A\�IA\JA��Q4K3�T0 k� �.�.14 'Q�1G�"H1  ��     �  �8A�$&�D]@@��`Fx<P]{�A\�HA\JA��Q4K3�T0 k� �.�.14 'Q�1G�"H1  ��     �  �8L= &�D]8A��`E�y<L]{�A\�HA\KA��Q4K3�T0 k� �,�,14 'Q�1G�"H1  ��     �  �8L= &�D]4C��`E�z<L]{�A\�HA\KA��Q4K3�T0 k� �*�*14 'Q�1G�"H1  ��     �  �8L=&�Dm,D\�`E�{<L]w�A\�HA\KA��Q4K3�T0 k� �)�)14 'Q�1G�"H1  ��     �  �8L=&�Dm$F\�`E�|<L]w�A\�HA\KA��Q4K3�T0 k� �(�(14 'Q�1G�"H1  ��     �  �8L=&|Dm G\�`E�}<L]w�A\�HA\KA��Q4K3�T0 k� �'�'14 'Q�1G�"H1  ��     �  �8L=&xDmI\�`E�}<H]w�A\�HA\KA��Q4K3�T0 k� �&�&14 'Q�1G�"H1  ��     �  �8L=&xDmJ\�`E�~<H]w�A\�GA\KA��Q4K3�T0 k� �%�%14 'Q�1G�"H1  ��     �  �8L=&tI�L\�`E� ~<H]w�A\�GA\KA��Q4K3�T0 k� �%�%14 'Q�1G�"H1  ��     �  �8L=&pI�M\�`E�$~<H]w�A\�GA\KA��Q0K3�T0 k� �%�%14 'Q�1G�"H1  ��     �  �8L=&lI�M\�`E�(~<H]w�A\�GA\KA��Q0K3�T0 k� � %�%14 'Q�1G�"H1  ��     �  �8L=&lI�N\�`E�,~<H]w�A\�GA\KA��Q0K3�T0 k� � %�%14 'Q�1G�"H1  ��     �  �8L=&hI�P\�`E�0~<D]w�A\�FA\KA��Q0K3�T0 k� ��%� %14 'Q�1G�"H1  ��     �  �8R	���E1�W@��B��|,���DјB�pEC;�!�r�T0 k� �C��C14 'Q�1G�"H1  ��"    � : SR	���E1�U@��B��|,���DјB�tEC7�!�r�T0 k� �A��A14 'Q�1G�"H1  ��"    � : SR	���E1�TP��B��|,���DјB�xEC7�!�q�T0 k� �@��@14 'Q�1G�"H1  ��"    � : SR	���E1�RP��B��|,���DјB�|EC3�!�q3�T0 k� �>��>14 'Q�1G�"H1  ��"    � : SR	���E1�QP��B��|,���DќB��EC3�!�q3�T0 k� �<��<14 'Q�1G�"H1  ��"    � : SUC	���E1�OP�B�#�|,���DќB��EC/�!�q3�T0 k� �;��;14 'Q�1G�"H1  ��"    � : SUC	���E1�L0w�B�'�|,���DѠBєE�+��r3�T0 k� �7��714 'Q�1G�"H1  ��"    � : SUC	���E!�J0s�B�+�|,���D�BјE�'��r3�T0 k� �7��714 'Q�1G�"H1  ��"    � : TUC	���E!�H0k�B�+�|,���D�	BќE�#��r3�
T0 k� �6��614 'Q�1G�"H1  ��"    � : UUC	���E!�F0g�B�/�|,���D�
BѤE���r3�
T0 k� �5��514 'Q�1G�"H1  ��"    � : VUC	���E!|D0c�B�3�|,���D�BѨE���r3�
T0 k� �3��314 'Q�1G�"H1  ��"    � : WUC�E!xC0[�B�7�|,���D�@�� E���r3�
T0 k� �2��214 'Q�1G�"H1  ��" 	   � : XUC�F�pA0W�B�7�|,���D�@��!E��
A�r3�
T0 k� �1��114 'Q�1G�"H1  ��" 	   � : YUC�F�h>0K�B�?�|,���D�@��"E��
A�r3�	T0 k� �-��-14 'Q�1G�"H1  ��" 	   � : ZUC�F�d< G�B�C�|,���D�@��#E��
A�r3�	T0 k� �+��+14 'Q�1G�"H1  ��" 	   � : [UC�F�`: C�B�G�|,���D��E��$E��
A�r3�	T0 k� �*��*14 'Q�1G�"H1  ��" 	   � : \UC�F�\9 ?�B�K�|,�D��E��$E���
q�r3�	T0 k� �(��(14 'Q�1G�"H1  ��" 	   � : ]ASA��F�X7 7�B�S�|,�D��E��%E���
q�r3�	T0 k� �|&��&14 'Q�1G�"H1  ��" 	   � : ]ASA��F�T5 3�B�W�|,�D��E��%E���
q�r3�	T0 k� �x%�|%14 'Q�1G�"H1  ��" 	   � : ]ASA��F�P4 /�B�[�|,�D��E��&E���
q�r3�	T0 k� �t#�x#14 'Q�1G�"H1  ��" 	   � : ]ASA��F�L2 +�B�_�|,�D��E��'E���
q�r3�	T0 k� �#��#14 'Q�1G�"H1  �" 	   � : eASA��F�H1 +�B�c�|,�D��E��(E���
��r3�	T0 k� �"��"14 'Q�1G�"H1 ��/ 	   � : mC� ��F�@. #�B�o�|,�F�E��)E���
��r3�T0 k� �!��!14 'Q�1G�"H1 ��/ 	   � : uC� ��F�<,��B�s�|,�F�E��)E���
��r3�T0 k� � �� 14 'Q�1G�"H1 ��/ 	   � : }C� ��F�8+��B�{�|,�F�E��*E���
��r3�T0 k� ����14 'Q�1G�"H1 ��/ 	   � : �C� ��F�4)��B��|,�F�E��+E����r3�T0 k� ����14 'Q�1G�"H1 ��/ 	   � : �C� ��F�0(��B���|, ��F�E� +E����s3�T0 k� ����14 'Q�1G�"H1 ��/ 
   � : �C����F�,'��B���|, ��F�E�,E����s3�T0 k� ����14 'Q�1G�"H1 ��/ 
   � : �C����F�(%��B���|, ��F�E�-e����s3�T0 k� ����14 'Q�1G�"H1 ��/ 
   � : �C����F�$$��B���|, ÷F�E�-eҿ��s3�T0 k� ��14 'Q�1G�"H1 ��/ 
   � : �C����F� #��B���|, ǸF�E�.eһ� ��s3�T0 k� ��14 'Q�1G�"H1 ��/ 
   � : �E� ���F�!��B���|,˸F�E�/eҷ� ��s3�T0 k� � �$14 'Q�1G�"H1	 ��/ 
   � : �E� ���F� ��B���|,ϹE� E�/eү� ��s3�T0 k� �,�014 'Q�1G�"H1	 ��/ 
   � : �E�����F���B���|,ӹE�C�0eҫ� ��s3�T0 k� �8�<14 'Q�1G�"H1
 ��/ 
   � : �E�����F���B���|,ۺE� C�1eҧ� ��s3�T0 k� �H�L14 'Q�1G�"H1 ��/ 
   � : �E�����F� �B�ú|,ߺE� C�1eң� a�s3�T0 k� �T�X14 'Q�1G�"H1 ��/ 
   � : �E�����F� �B�Ǻ|,�E� C�2eҟ� a�s3�T0 k� �`�d14 'Q�1G�"H1 ��/ 
   � : �E�����F� �B�Ϻ|,�E�!C�2eқ� a�s3�T0 k� �l�p14 'Q�1G�"H1 ��/ 
   � : �E�����F� �B�׹|,�E�!EB3eқ� a�s3�T0 k� �|��14 'Q�1G�"H1 ��/ 
   � : �E�����F� �B�߹|,��E�$"EB3eҗ� a�s3�T0 k� ���14 'Q�1G�"H1 ��/ 
   � : �E�����F�  �B��|,���E�("EB4eғ���s3�T0 k� ���14 'Q�1G�"H1 ��/ 
   � : �E���ÍF�� �B��|,���E�0#EB4eҏ���s3�T0 k� ���14 'Q�1G�"H1 ��/ 
   � : �E���ǍF�� �B���|,��E�8#EB4eҋ���s3�T0 k� ���14 'Q�1G�"H1 ��/ 
   � : �E���ˍF�� �B���|,��E�<$EB5e҇���s3�T0 k� ���14 'Q�1G�"H1 ��/    � : �E���ύF�� �B��|,�E�D$C�5e҃���s3�T0 k� ����14 'Q�1G�"H1 �/    � : �RR��ӍF�� �B��|,�E�L%C�5e����s3�T0 k� "���14 'Q�1G�"H1 ��/    � : �RR��׎E ��B��|,�E�P%C�5e�{���s3�T0 k� "���14 'Q�1G�"H1 ��/    � : �RR��ߎE ��B�#�|,'�E�`%C�5e�w���s3�T0 k� "���14 'Q�1G�"H1 ��/    � : �RR���E ��B�+�|,/�E�h&C�5e�s��s3�T0 k� "���14 'Q�1G�"H1 ��/    � : �RR���E ��B�3�|,7�E�p&C�5e�o��s3�T0 k� "���14 'Q�1G�"H1 ��/    � : �RR���E �
 �B�;�|,�?�E�t&C�5e�k��s3�T0 k� ����14 'Q�1G�"H1 ��/    � : �RR���E �	 �B�C�|,�C�E�|&C�5e�k��s3�T0 k� ����14 'Q�1G�"H1 ��/    � : �Rb����E� �B�K�|,�K�E��&C�5e�g��s3�T0 k� ����14 'Q�1G�"H1 ��/    � : �Rb����E� �B�S�|,�S�E��&C�5e�c���s3�T0 k� ����14 'Q�1G�"H1 ��/    � : �Rb���E� �B�[�|,�[�E��%C�4e�_���s3�T0 k� ����14 'Q�1G�"H1 ��/    � : �Rb���E� �B�c�|,�_�E��%C�4E�_���s3�T0 k� 2���14 'Q�1G�"H1 ��/    � : �Rb���E� �B�k�|,�g�E��%C�4E�[���s3�T0 k� 2���14 'Q�1G�"H1 ��/    � : �Rb���E�#�B�s�|,�o�E��$C�4E�W���s3�T0 k� 2���14 'Q�1G�"H1 ��/    � : �Rb���E�'�B�w�|,�w�E��$C�3E�S���s3�T0 k� 2���14 'Q�1G�"H1 ��/    � : �Rr��E� '�B��|,��E��$C� 3E�S���r3�T0 k� 2���14 'Q�1G�"H1
 ��/    � : �Rr�#�E��+�BЇ�|,у�E��#E� 3FO���r3�T0 k� ����14 'Q�1G�"H1
 ��/    � : �Rr�'�E��/�BЏ�|,ы�E��#E��3FK�� r3�T0 k� ����14 'Q�1G�"H1	 ��/    � : �Rr�3�E���7�BП�|,ћ�E��!E��2FG��q3�T0 k� ����14 'Q�1G�"H1 ��/    � : �Rr�;�E���;�BЧ�|,ѣ�E��!E��2FG��q3�T0 k� ����14 'Q�1G�"H1 ��/    � : �Rr�?�B����?�BЯ�|,ѫ�E�� E��1FG��p3�T0 k� "���14 'Q�1G�"H1 ��/    � : �Rr�G�B����C�Bз�|,ѳ�E��C��1FC��p3�T0 k� "���14 'Q�1G�"H1 ��/    � : �Rr�K�B����G�Bп�|,ѻ�E��C��1FC��o3�T0 k� "���14 'Q�1G�"H1 ��/    � : �Rr�S�B����K�B�Ƕ|,���E��C��1E�C�� o3�T0 k� "���14 'Q�1G�"H1 ��/    � : �Rr�[�B����O�B�϶|,���E��C��1E�?��$n3�T0 k� "���14 'Q�1G�"H1 ��/    � : �Rr�_�B����S�B�׶|,���E��C��0E�?��,m3�T0 k� ���14 'Q�1G�"H1 ��/    � : �Rr�g�B���T B�۵|,���E��C��0E�?��0m3�T0 k� ���14 'Q�1G�"H1 ��/    � : �Rr�o�B���\B��|,���E� C��0E�?��4l3�T0 k� ���14 'Q�1G�"H1 ��/    � : �Rr�s�B���`B��|,���E�C��0E�?��<k3�T0 k� ���14 'Q�1G�"H1 ��/    � : �Rr�{�B���dB��|,���E�C��/E�?��@j3�T0 k� ���14 'Q�1G�"H1 ��/    � : �Rr���B���lB���|,���E�C�/E�?��Dj3�T0 k� B���14 'Q�1G�"H1  ��/    � : �Rr���E��pI�|,��E�C�/E�< �Li3�T0 k� B���14 'Q�1G�"H1  ,�/    � : �Rr���E��|	I�|,��E�C�/E�<�Xg3�T0 k� B���14 'Q�1G�"H1  ��/    � : �Rr���E#���I�|,��E�C�.E�<�\f3�T0 k� B���14 'Q�1G�"H1 ��/    � : �Rr���E+���I�|,�#�E�C�.P�@�de3�T0 k� ���14 'Q�1G�"H1 ��/    � : �Rr���E/���I'�|,�+�C�C�.P�@�hd3�T0 k� ���14 'Q�1G�"H1 ��/    � : �Rr����E�3���I!+�|,�3�C�C�.P�@�pc3�T0 k� ���14 'Q�1G�"H1 ��/    � : �Rr����E�?���I!7�|,�C�C� Eф-P�@�|a3�T0 k� ���14 'Q�1G�"H1 ��/    � : �Rr��ǰE�G���I!?�|,�K�C� E�|-P�@�`3�T0 k� "���14 'Q�1G�"H1 ��/    � : �Rr��ϱE�K���I!C�|,�S�E� E�t-QD	��_3�T0 k� "���14 'Q�1G�"H1 ��/    � : �Rr��ӲD�S���IG�|,�[�E� E�l-QD	��^3�T0 k� "���14 'Q�1G�"H1 ��/    � : �Rr��۳D�W���IO�|,rc�E� 
E�h-QD
��]3�T0 k� "���14 'Q�1G�"H1 ��/    � 9 �Rr���D�c���IW�|,rs�E� E�X,QD��[3�T0 k� "���14 'Q�1G�"H1 ��)    � 8 �Rr���D�k���I[�|,r{�E� E�P,QD��Z3�T0 k� �|��14 'Q�1G�"H1 ��)    � 7 �Rr����E�s���I!_�|,r��E�EQH,QH��Y3�T0 k� �x!�|!14 'Q�1G�"H1 ��)    � 6 �Rr����E�{���I!c�|,r��E�EQ@,QH��Y3�T0 k� �x"�|"14 'Q�1G�"H1 ��)    � 6 �Rr���E�����I!k�|,r��E�EQ0,QH��W3�T0 k� �t$�x$14 'Q�1G�"H1 ��)    � 6 �Rr���E�����I!o�|,r��E�EQ(+P�H��V3�T0 k� 2p%�t%14 'Q�1G�"H1 ��)    � 6 �Rr���P��	�Is�|,r��E�EQ +P�H��U3�T0 k� 2l%�p%14 'Q�1G�"H1 ��)    � 6 �Rr��#�P��	�Iw�|,r��D3EQ,P�H��T3�T0 k� 2h&�l&14 'Q�1G�"H1 ��)    � 6 �Rr��+�P��	�I{�|,r��D3EA-P�H��S3�T0 k� 2h&�l&14 'Q�1G�"H1 ��)    � 6 �Rr�3�P��	�I{�|,r��D3EA.P�H��R3�T0 k� 2h&�l&14 'Q�1G�"H1 ��)    � 6 �Rr�C�P��	 �I��|,r˦D3 EA/E�H��P3�T0 k� �d&�h&14 'Q�1G�"H1 ��)    � 6 �Rr�G�P!��	 �I!��|,bӥD3 EA0E�H� O3�T0 k� �d&�h&14 'Q�1G�"H1 ��)    � 6 �Rr�O�P!��	 �I!��|,bףD3 E@�1E�D�O3�T0 k� �`&�d&14 'Q�1G�"H1 ��)    � 6 �Rr�W�P!��	 �I!��|,bߢD3�E@�1E�D�N3�T0 k� �`'�d'14 'Q�1G�"H1 ��)    � 6 �Rr�_�P!��	 �I!��|,b�D3�E@�2E�D�M3�T0 k� �`'�d'14 'Q�1G�"H1  ��)    � 6 �Rr�g�P!��	�I!��|,b�D2��E@�2ErD�L3�T0 k� "\(�`(14 'Q�1G�"H1  ��)    � 6 �Rr��o�P!��	�I��|,b�DB��E@�2Er@� K3�T0 k� "X)�\)14 'Q�1G�"H1  .�)    � 6 �Rr��{�P!��	�I��|,b��DB��E@�3Er@�0I3�T0 k� "T*�X*14 'Q�1G�"H1  ��)    � 6 �Rr����P!��	�I��|,b��DB��E@�3Er@	�4H3�T0 k� "P+�T+14 'Q�1G�"H1  ��)    � 6 �Rr����P�� ��I��|,b��DB��E0�4Er@	�<G3�T0 k� �P,�T,14 'Q�1G�"H1  ��)    � 6 �Rr����P�� ��I!��|,c�DB��E0�4Er@	�@G3�T0 k� �P-�T-14 'Q�1G�"H1  ��)    � 6 �Rr����P�� ��I!��|,S�DB� E0�4Er@	�DF3�T0 k� �P.�T.14 'Q�1G�"H1  ��)    � 6 �Rr����P� �� I!��|,S�DB� E0�4Eb@	�LE3�T0 k� �@,�D,14 'Q�1G�"H1  ��)    � 6 �Rr����P� ��"I!��|,S�DB� E0�4Eb@
PE3�T0 k� �4,�8,14 'Q�1G�"H1  ��)    � 6 �Rr����E��0�#I!��|,S�DB� E0�4Eb@
TD3�T0 k� �,,�0,14 'Q�1G�"H1  ��)    � 6 �Rr����E��0�&I��|,��DB�E0�3Eb@
\C3�T0 k� � .�$.14 'Q�1G�"H1  ��)    � 6 �Rr����E��0�(I��|,��DR�E0�3Eb<
`C3�T0 k� �.� .14 'Q�1G�"H1  ��)    � 6 �Rr�s��E�'�0�)I��|,��DR�E0�3Eb<	�hB3�T0 k� �/�/14 'Q�1G�"H1  ��)    � 6 �Rr�s��E�+�0�+I��|,��DR�E0�2Eb< 	�hB3�T0 k� �0�014 'Q�1G�"H1  ��)    � 6 �Rr�s��E�3�0�,I��|,��DR�E �2Eb8!	�lB3�T0 k� �1�114 'Q�1G�"H1  ��)    � 6 �Rr�s��E�7�0�.@a��|,S�DR�E �2ER8"	�pB3�T0 k� �+�+14 'Q�1G�"H1  ��)    � 6 �Rr�s��E�?�0�/@a��|,S�DR�E �1ER8$	�tA3�T0 k� �'�'14 'Q�1G�"H1  ��)    � 6 �Rr�s��E�C�0�0@a��|,S�DR�E �1ER4%
xA3�T0 k� �'�'14 'Q�1G�"H1  �)    � 6 �Rr�t�E�O�0�3@a��|,S#�DR�E �/ER0'
|A3�T0 k� ��%��%14 'Q�1G�"H1 ��/    � 6 �Rr�t�E�W�0�4@���|,S#�DR�E |/G�0(
�A3�T0 k� ��%��%14 'Q�1G�"H1 ��/    � 6 zRr�t�Er_�0�6@���|,S#�DR�E x.G�0)
�A3�T0 k� ��$��$14 'Q�1G�"H1 ��/    � 6 rRr�t�Erc�0�7@���|,S�Eb�	E t.G�,*	�A3�T0 k� ��#��#14 'Q�1G�"H1 ��/    � 6 kRr�t#�Erk�0�8@���|,S�Eb�
E p-G�,+	�A3�T0 k� ��"��"14 'Q�1G�"H1 ��/    � 6 dRr� d'�Ers�0�:@���|,C�Eb|E l-G�(,	�A3�T0 k� ��"��"14 'Q�1G�"H1 ��/    � 6 ]Rr� d/�Erw�0�;A��|,C�EbtE h,G�(-	�@3�T0 k� ��!��!14 'Q�1G�"H1 ��/    � 6 VRr� d3�Er�0�<A��|,C�EblE d,G�(.	�@3�T0 k� �� �� 14 'Q�1G�"H1 ��/    � 6 PRr� d;�Er��0�=A��|,C�ERhE `+G�$/��@3�T0 k� �� �� 14 'Q�1G�"H1 ��/    � 6 JRr� d?�Er��0�>A��|,C�ER`E \*G�$0��@3�T0 k� �|��14 'Q�1G�"H1 ��/    � 6 DRr�!dC�Er��0�@A��|,��ERXE X*G� 1��?3�T0 k� �l�p14 'Q�1G�"H1 ��/    � 6 >Rr�!dK�Er��0�ACᗵ|,��ERPE T)G� 2��?3�T0 k� �`�d14 'Q�1G�"H1 ��/    � 6 8Rr�!dO�Er����BCᗵ|,��ERHE T)G� 2��?3�T0 k� �T�X14 'Q�1G�"H1 ��/    � 6 2                                                                                                                                                                            � � �  �  �  c A�  �J����   �      6 \��|j ]�++ � �� &  � �
   ��A�:     &��B-�    �L��   	           Y Z�8�         ��      ���   0
           �;   � �     ��Z,     7B�Z�U    i�g               c Z�8         ���     ���   8	           Q`8  � �	      �@"     P7Q�A;    ��9            	 Z�8         ���    ��� 0
           `QP   � �	   �-�l     `QP�-�l                    	 Z�8          %�     ���   0

          ~>�  Z Z    .��     ~ng�1V    ���               Z�8          �@�      ���  8	
'	            Bb  ��     B��     Bb��      ��                   
	  ��8              c  ���    		 5            �� �        V�]?�    �� ��]R�      ��             	 c �         0  �  ��@   H

          F�O       j�1��     G<��2�    �c��          	 6 �         �  �  ��@ @ (
           K��        ~��]     K�����     �                "          ��     ��H   (G            ��6N  ~
	  ���L    ��=���    ���p             	     �         	 �   �  ��@   H
	(
           Km        � LӢ     KjU L��     )�+               A �         
 �  �  ��@   0
		H
          �\ ��     � �     �\ �                              ����              �  ��@    0

 3                  ��      �                                                                           �                               ��        ���          ��                                                                 �                          %��  ��        ��?�     %�1�@e�    �I�{                   x                j  �        �                          %    ��       ��@       %  �A           "                                                 �                         �A�Z�A�-���]�1��� L ����?�@ 	 
               
  �    �T� u��_      ���� ���� ���� ����  ����. ����< ����J ����X � �� 0�  �� 0ƀ �( 0�  �� 0ŀ �h 0�  � 0Ā �� 0�  �H 0À �� 0�  �� 0 �( 0�  �� 0�� �h 0�  � 0�� �� 0�  �H 0π �� 0�  �� 0΀ �( 0�  �� 0̀ �h 0�  � 0̀ �� 0�  �H 0ˀ���� ����� ����� � � �[� � \� ä }@ � �m@ � n@ -d �o� .� p� .� q  �d �t� �d u����� � � �t� �  u� �D v  AD �r@ BD  s@ B� s� �� w@ � �w` �$ x� 
�\ U� 
�� V  
�| V  
�\ V� 
�� V� 
�| W  
�< W� 
� W� 
�| W�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����8��  �� �  ������  
�fD
��L���"����D" � j  "  B   J jF�"     
�j,
 ��
��
��"  ""B�j��" 
 �
� �  �  
�  &    ��     ��B       &    ��     ��B       K    ��     ��          � ��   �  � ��        LL     �    ��        MM     �    ��        a�         �    ��  � G      �� � �  ���        � �  ���        �        ��        �        ��        �    ��     ���  �        ��                         ���   	�� ��                                    �                ����              &�B ���%��    �8��                18/41 (43%) ebeau  s   5:02                                                                        2  2     �� �� �k~#1 k�#
K.X K4X K5P K6H �	CB �
CJ �CM � CO � �C< �C< �C $ �C# � C'4 � C(# �kj kr � � � � � . �K) �K9 �J� � �J� � J� � J� �J� �B� � � B� � � !B� � � "B� � �#cV u � $c^ } �%"� � � &"� �'� � �(
� �)"� � � *"� �+"� � �,*�1-"�1 ."�1!/�!0
�* �1*:� �2)��3*<�8 4*LhX 5*KXP  *Rp  *Kj  *Kj  *Kj *<j;*r <*FjF  *GjL  *Gh  *Gr                                                                                                                                                                                                                         �� R              @ 
      N �     \ P E e  ��                     �������������������������������������� ���������	�
��������                                                                                          ��    �>|�� ��������������������������������������������������������   �4, C  $ # ���@��k��ς�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               "    %      �  K
�J      ~�                             ������������������������������������������������������                                                                                                                              	          �  �                  ��      �   j          	 	 
  	 
 
 ��������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� ���������������������                                 .    )    ��  $>�J      �  	                           ������������������������������������������������������                                                                                                                                             �  ���                      �        �          	     ������ ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ������                                                                                                                                                                                                                                                                           
                              	                   �             


           �   }�         wwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwww 0 I =                                  � M�W �\                                                                                                                                                                                                                                                                                    )n)n
  �                                        m      k      `                                                                                                                                                                                                                                                                                                                                                                                                                � � �  � ��  � @��  � (��  � (��  � Z��  �����x�����������M����������w����Ҡ����Ѡ����s4                      � s           �   & AG� �  �                 �                                                                                                                                                                                                                                                                                                                                      0 F I   �                       !��                                                                                                                                                                                                                            Y��   �� � ���      �� @      ��������������������� ��������� �� �� ���������������������������� ��������������� ������  ��������������� �������� � ������������ ��� ��� ���� ������������   ������������� � ������������������ ����� ������� ��� ��������������������������� ��� ���������  �������� ���������� �� ������������������� ��������������������������������������  � ��������������������������� ��� �� ��� ������ � ������������������������������������������������������� � ����� ������ � ������              ���������������������������������������������������f��ff�fff�ff���������l�ff�ffffl��ff˼fllf������l��̼�ʗ���˹�ffjz�fkyl�l��fƨ�����������������������̼��̉������������������������������f���f�fff�ff�ffl�ff�flfl�l��xl�wwl���l̻�����˺��fl����l�xx��w��̻���l�f�f�ƻ�fl�����ffl�ffffffff���f���̚���ffflffflfffffffffflfffff������������������������l���l������f����������������������������l��lf��f�fff�f��l˪���ww��w�����flflffffffff�̼̙��fww��w��fx�̻�llffff�ffff���fl���f�l�l�˶����fffl��fflfll����ff��ff��lfl�lf��l���l�����������l�������l�������ʼ�j˚��̩��ʨ��ɘ���xxxȈ��ɉ�x���̇�̺������www��ww��xw���x��xk�����������wx��������������x����l�ƈ��Ƈ���w��Ɨ��̩z�̩yf̪�f�������������������������������̙i���ɖ�yɌ��ˌȉ̚ə̩���ə��Ɉ����x�̹x�̹�����������ƺ�������������������ˈ������˙������̫��̺�������˪�������������̸��̗�����̇��̇�����������������������̈���xx����x���w���ɉ��̨���k���̛̻�������������l��Ʀl�Ɗl�l���̻�lk��̺�f̩�l��f�ɫ�ˉ�lɊ�˙���ʚ���˙�˫̼���ɬ�̚��̼�����̼���̬������̼�����˻������������f����˺�xfl˙z�f������������y������˪�����˥�l�U��www���������wYuU��UY��x������������W���U�f��Vf������������������������f���ff���m�    7      8   �  %                       @     �  �����J���J      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �f ��        p���� ��   p���� �$     `d     �f ��     �f �$ ^$ �@      ����� ��   ����� �$ ^h   ����  ��   ����  �$ ^$     �                      ��� ���� 
"�������������� x��+&  ��+ &         ��   .���x � ��� �� � ��� �$ ^$  ��     Td���2 9 ���J���� �   Q ��@              ��  yf  y<  �!"wr27Cr#G4r3w72#w4t2"Cwt3wG}�wwwwwtwwww4wwGwwwwww��tw�wwwwwwDw��G��w�w���y������w���wy������w�K���t��{���GwKDDCDDt333wwDDDG�DD�~DDD�DDNDDw�DD�tDD~~DDwGDDDDDGDDDuDDGVDDucDGV3Duc3GV33uc33Vffffffffffffffffffffffgfff~ffg�ff~Nfg��f~N�g���~N������N~�����w�www�www�wwwwwwwwwwwwwwwwwwwwwwwwftDwvdDwvgDwwfDwwftwwvdwwvgwwwfDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD#vd�2eU�3Fff3t�G4��D�D,�CG��}�t�wwt�wtw�wOw�w�wOD�w2?�wCOGww�D��H��GH���I���y���y���t��Os#wt4�w�����2���������(�wy������ww���s4��4��tO��t��}w�B4W�DEFwt3G4wCGGGtt�Ctw��wG�Gtw�TwtfEwJ{�Gwz��w���wt�Gw��wt�Gw�wtw�{�GD���D���D���N���GfgvDDDDDDDDDDDD����������������fwfgDDDDDDDDDDDDww��w��w2��w���w��w���x�wy����w"GC42wsDCwt�Cwt��ws�DGt�T7DfEGtwwwwwwwwwwwwwwwwwwwwt3GwsOGwt��wNNNNNNNNNNNNN���FfwfDDDDDDDDDDDDDvUwGfewwvffwwGw��w��G}��w���w����y���w�w�w��www��wwwwwwwwwww�w4wwwwwwBGDwsG3GwwC7wwtGwwDwGwV333c33333333336333f336g33f~36g�ff~Dfg�Df~DDg�DD~DDD�DDDDDDDDDDD��~wN��wD��gDNwvDD�wDN�wD���N�N�wwwwwwwwwwwwwwwwgwwwvwwwwgwwwvwwwwwfwwwvwwwvwwwwwwwwwwwwwwwwwwwwtDDDdDDDgDDDfDDDftDDvdDDvgDDwfDD�����}���}�}���}}��}}�w~I�D�t�y�wts"�wB2�w22�s#C�s#4�w2t�ws�www�3#�w""7w##'wCC#wDG2w3G~������ww�����y���w�����y��Gwwwwt33Dt343�wVt�wUv�wen�wvW�wv��wt�wtGDw�fuG�dvW��Vg��fw�wGw�D�w��w�t�wt����K���{�K�{�{�t�{�wG~�Gt��y�wD�w�N���N���N���N���NDDNNww~D���fuGwdvWw�Vgw�fwwwGwwD�ww�wwt�wwwwwt��wH��wHIIwIyy�y�Gwwt4wt4CGDwwwGwDwwDDGwG�Gt��w�GwEGwvfTw���w}���}�}�w�w�y��wwI��wwI�wwwwwwtwwwDwwwGw�www�wtw�www�www�www"4w#Gw"4ww#Gww4wGwGwwww{w�{��DDDDDDDNDDD�DDN�DD��DN��D���N����������N����www�ww��ww~�~�w~��~��wgw�wvw��wgN�wv���w�N�w������N�w��Hwy�Iwy�Iwt�ywy�ywt�tws#swt4twwwwwwwswww4wwtOwwt�wwwww4WwwEFw$t747wGDGtw�Cww��ww�DGw�T7wfEGwvfTgFFVGFDeDUgFeI�teI���t���wwwIwwwwwwwwwwwwO�wGN�t4�G7G��tt��ww"4w#Gw"4w#Gww4w��Gw�ww4wws3w��������������������D���DN��DDN��������N������������������������wwwfwwwvwwwvwwwwgwwwvwwwwgwwwvwwwwVtwwUvwwenwwvWwwv�wwtwwtGww�"4w#Gw"4w�#Gt�4w�wG�www��wIwwDt��GO��wO��w�O�t���O���G4w�23wwftDwvdDwvgDwwfDgwftvwvfwfffffffDf��DvDGNwDNN�GfDGfwfGwwwGgwwGfw#w�2G22""##3?3333323232#333333t�3""""33�333�333333323333333333""""3�3838383�38383333323"333#33FfffGwwwGwwwGwwwGwwwGwwwGwwwGwww""""��33�?33�?33�?333333#23323#3ffffwwwwwwwwwwwwwfgvwwwwwwwwwwwwffffwwwwwwwwwwwwfwfgwwwwwwwwwwwwr"""s3?�s3?3s3?�s3?3s323s3#3s333""""3�333�333�333�3333333"333333ffffwfwfwvwvwfwvwvwvwwwwwfwvwgww""""33?�33?�33?333?333333323#333"""'3�37?�37�3373337#33733373337DDDFDDDeDDFVDDefDFVfDeffFVffeffft��wt��wt�x�t�DwwDD7wwwDwDGtwwwwDwwwGwtGwtDDwt�wG��ww�w27�s"$w����������������N��fN�fw�fwwfwww���f��fw�fw~fwwwwwwwwwwwwwwwwwwwffffvffgwffg�vfg~wfgw�vgw~wgww�wwGwwwGwwwtwwwtwwwtwwwtwwwtwwwtwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwwCGwtDDwtGww��ww�Gwt�ww{�w�K��C3#w332t342CC7C3�Gt4O��DtO��wwtO�ww>�Gw7wtwGDwwwwGw�wwtOGwD��ww��ww��wt|}ww|sGw}t4ww4wwtCGwwwwww�ww��wwG��wG��wG���N~��D~��D~�www~�ww�ww�ww�wwwwwwwwwwwwwwtwwtGwtwwwtwwwtwwwtwtwttGwDGwDwGwwwGwwwwwwwwwwtDDDGwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwDDDDwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDDGwwwGwwwGwwwGwwwGwwwGwwwGwww�!"wr27CwsG4C4w74�w7O�rGw�3wHw��Oww�wwO�#wOGwwt24wwDGtGwwwtwwGDDDDDDDNDDDDDDN�DDDDDN��DDDDN���D~ww��wwD�ww�GwwDGww�GwwDGww�GwtwwwwwwwwwwwtwwtGwwGwwDwwDwwwwwwwwtGwtGwwGwwwwwwwwwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGwwwGwwwGwwwGwwwGewwwwwwwwwwwwwwwwwwwwwwwfve3333UUwwwwwwwwwwwwwwwwwwwwU3333UUUUUUUwwwwwwwwwwwwwwwwwwww3333UUUUUUUUGwwwGwwwGwwwGwwwGwwwC333EUUUEUUU���w}���}�}�wC4�w4�wwO�www��wHwwDDDDD�DDDDN��DDDw�DD�tNDNtDD�~DD��G�NtgDD~�DN�G�NvgDD��DDDDNDDD�DDDD����DDDD����DDDD���FDDDg��FwDNtG�DGwDDwwDdwwvtwwgtwww~wwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwewwe3wwwwwwwwwwwewwe3we3Ue3UU3UUUUUUUwvC3e3EU3UvUUUfUUUgUUUTUUUTUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUVwVwl�UUUUUUUUUUUUUUUUUUUUUfwwv�������UUUUUUUUUUUUUUUUUUUUwwww��������EUUUEUUUEUUUEUUUEUUUGwwwl���l���D��wDDNvD��vDDNwD��wDDNvD��vDDNwDDDDDDDDDDDDDDDDD��wDDNvD��vDDNwN�DDN�DDD�DDDNtDD���DDDDDDDDDDDDDDgw�FwwDgwwFwwwgwwwwwwwwwwwwwwwwwGwwwGwwwGwwwGuwwFSwwd5wu4UwSTUwvSUvS5Uc5UU5UUUUUUUUUUUUUUUUUUVUUUUUUUUUUUUUUUgUUglUgl�Wl�U|��UUUTgUVv�fv��l��U��UU�UUSUU5SUSSSl�����UU�UUUUUSSU555SS333300303�UUUUUUUU555SSSS333330000  UUUUUUUUSSSS555533330000    eUUUUUUUU555SSSSS333SP000P   UUUSUUU3SSS%53"532#33" 00"   vEUU�geU�\gfU\��UU3�5R5\5#UU355UUUUUUUUUUUUUvUUU�vUU��vUS��u"\�ǘIww�ywG�2#w�www2#GwtDwGwwtGwtwwDDDD����DDDD����DDDD����DDDG���FDDgw�FwwDvww�gwwFwwwgwwwgwwwwwwwwwwwwwwwwwwuwwwSwwu5wwSUwu5UwcUUu5TUSUTe5UWuUUVEUUUEUUUFUUVGUUgeUUVfUUg�UV|�Vv��g��U|�US��S3�UU3��UU�USSUU53U333533S300300   353S330U30303                                                                        0  0   0  0                 0   0   0   0                         #                   02   "     "     "     "   %3S23"P32#P "P 00"    "   %U\�55S�3S2%33"U02#S"352#33"003feUU�vUU��eU\�geU��v3#��2%\�"5U\D��wDDNvD��vDDNwD���DDDNDDDNDDDDDDDDD���DDDDD���DDDDD���DDDDD���DDDD����DDDD����DDDD����DDDD����DDDg��GgDDDw��gGDGg��Fw~Dvwt�gwtwwwwwwwwwwwwwwwuwwwSwwu5wwcUww5Uv5UUcUUUSUUU5UUUUUUVUUUWUUUfUUV|UV|�Ug��V|�Vg��U|�US��U5�US3�U33UU30U533S330U3c000c3 c  P0  0                                                    �� ������                    ������������                 ������������                 ��� ��� ����      "     "     "     "         "     "     "     "    2   "  #  "     "     "   #3UR33S%32500#U6  36 06  vfTgFDDwFGGGUGGG��w��G}��w���wDgw~GgwwFwwwFwwwvwwwgwwwgwwwgwwvwu5U�cUUGSUUF5UU�UUUwUUUTUUU4eUVUUg�UV|�Ug�UU|�UVl�Sg�U5|�SSlU53US3U300S33053 S00 3  00        6      0   P   P   0      ������������������ ��� �������������������������������������������������������������������                            ���w}�Dw}DDGwG�GtD��wD��wEGwvfTw�O�w���wwO���wGw��w��G}��w���wDDDDD���NDDDD��NDD�D����~DDD����DDDF���FDDDv���gDDDg���gDDGg��FwwwwuwwwswwwSwww5wwv5wwu5wwcUwwcU7eUgVuU|UEVlUFW�Uvf�Ug|�UTl�UWlS������������U30 SS U00 3  S0  ������������                    ������������  9�  	�  �  �  �8888����������������������������3������3���8  "     "     "   3�����������                    vd4wFDDGFG�wW�ww�wt�ww{�w�K���O�G����t�O�t���O��OG�w�Gww�"4w�DDDD���NDDD�����DDDD�D�DDDDD���DDFw��FwDDvw��vwDDgw��gwDDgw��gwwwSUwv5Uwv5Uwu5UwsUUwcUUwcUUwSUUUfUUU|�SU|�5VlVSW�U3f�SS|�Uc|�SS3  00  3   3   0       0          �   9   9                  �������ߨ���������������	������                                37��s��7�w���y������w���wy���DDGw��twDDdw��dwDDgG��gGDDgG��gtw5UUv5UVv5UWu5UWu5UWsUUfsUU|sUU||�53lUS5�U35�SS�U30�S3 �50 �S3                 0   0                                       ��                        8������� 9�� �� ��  9�  �   9       �����������������������߉���8�������y�D�tDDyt�wG��ww��wtTwwvegwDDgt��gtDDgw��gwDDgw��gwDDgw��gwsUU|sUVlCUV�EUW�FUW�tUW�tUW�veW��S0 �30 US0 U30 US  U30 SS  U3                     8  � �� ���       � ��8�����0 �0  0       8������ �0                       ��� ��  �   8                ����������������8��� 8��  �    ����������������������������8�����������������������������������DDgw��gwDDgw��gwDDgw��gwDDgw��gwuuW�svW�sgW�sTW�sWg�sVw�sUG�sUg�SS  U3  SS  U3  SS  U3  SS  U3            9  �  9� �� �0 9� 8�� ��  �0  �   0                ��                           ��������  33                    ywwD�twwysww�wwwC#GwtDwwwwwGwwtwsUW\sUWlsUWUsUW�sUW�sUW�sUW�sUW�                     9   ������� 	�0 ��  ��  �0  �   �   �   sUW�sUW�sUW�sUW�sUW�sUW�sUW�sUW�US  V3  US  US  SS  US  SU  U5  ����   �  �  �  �  	�  9�  9��   0                                                 �  9� ������y�tGw�DDwt�wG��ww�w27�s3$wsUW�sUW�CUW�EUW�FUW�tUW�tUW�veW�SSP U3P SS  U3 SS  U3 0SS  U3  UuU7�uU7UuU7luU7\uU7�uU7�uU7<uU7  53  3#  2%  "U %5 "3U 55" 3S�uU7�uU7�uU7�uU7�uU7�uU7�uU7<uU7 52 3%  25 P#U 55 3U 55  3U                                                              �uWW�ug7�uv7�uE7�vu7�we73tU7<vU7                                 """ "!"! ! """"  " 5uU7�uU7UuU7luU7\uU7�uU7�uU7<uU7ffffwwwwwwwwwwwwwwwwwwwwwwwwwwwwffGwwwtwwwtwwwtwwwwGwwwGwwwGwwwt                                                           wwwwwwwwGwwwGwwwGwwwtS33weUUuuUUwwwtwwwtwwwwwwwwwwww3335UUUUUUUUsvUUsgUUsTUUsWeUsVuUsUGwsUg�sUW�SS U3  SS U3  SR  U#  RS  53     �  �  �  �  �� 
�w ��~����   ��  ��  �p  }`  g`  w       ���˜��̽���ͻ�ۧ�̺�w̚�~�����   ��  ��  �p  }`  g`  wU  �CP ���̌˜��̽���ͻ�ۧ�̺�w̚�~�����#0 ��  ��  �r  }h� gk� wU� �CP �#0 ��" ��"/�r""}h�gk��wU� �CP �����ۻ���������_��UU  SU  U5  ��������ۻݽ�۽�����            ������ۻ�ݻ�ݽ������            ��������������������������˚��̸���̽��̍̽��̽�����̻#0 """ 3""/�"""�(��+��U� �CP ���������J�S�T33����������������#0 """ 3""/3"""��M������ ܪ� UuW�UvW�UgW�UTW�UWg�www�������������www@Gww0$ww0wwswwt        +�  "�" ""/�"""����                                     ��                        ��ݻ����                   �  � �� ���       � ���۽���� ��  �       �ۻ�۽� ��                                          3333UUUUUUUU�uU7�uU7�uU4�uUT�uUd335GUUVwUUWW          �  �  �� �� �� �� ��� ��  ��  �   �                                             9             9� 9���� ��0 ��       ��������3 0               3�����������  3U  55  3U  55  3UE     P ` @  E F  d3333ffffffffffffffffffffffffffff                     �   �   ��� �� ��  ��  ��  �   �   �     �  8�  �� �0 9�  ��  �� �0 �                               ffffffffffffffffffffffffffffffff  T   &    331ff6fff6fP   `   @   E   F   t   tP  v`  ffffffffffffffffffff3333UUUUUUUUSS  U3  SS  U3  SS  ��������U9�0                    ����������0                 ����������2                   ���������*0                   �3������#��0   �   �  �  �  ߃����������                    8888��������  	�  9�  :�  ��  :�88����	��0DD@���DD@���DD@���DD@���ffVfffVfffVfffVfffVfwwgwDDgw��gwuu  sv  sg  sT��sWl�sVw�sUG�sUg�UUUUUUUUUUUU�UU�gw������#*�2��3333!#! ! """"  " ��0���0���0                    	��0��� 8��                    DDGfDDGwDDDwDDDvDDDwDDDGDDDGDDDGS33qU7�aSW�q5W<qUU�aU7�qSW<q5U�qU7�qSW<qUU�EU7�FSW�E333GfffDfffDfffDvffDFffDFffDGffDDwwDDDDDDDDBDB'G trpwG't7w Btr                    3333ffffffffffffffffffffffffffffwwwwDDDDDDDDU3P SSP US  �����ݽ��ݽ���������                     DDvw��vwDDFw��FwDDFw��FwDDFw��FwDDGg��GgDDDg���gDDDg���gDDDv���vDDDF���FDDDG����DDDD����DDDD����v5W�v5W�f5W�f5W�g5W�v5W�FSW�FcW�GcW��cW�DvW��FW�DFg��Gg�DG6���V�DDc<��u<DDv1��F1DDGc��GeDDDe���vS  e!  e0 v2 FS Ge8De8��vS�DFe0�Ge2DDfS��veDDGf���vDDDF���GA   e  V  4  TPdPdc  ds                              A   @!  @ e  !V                         !                                                                DDDD����DDDDN���DDDDDN��DDDDDDN�wE0 GFS DFe0�GfSDGfe��vfDDGf���v          0  S  e3 fe0      &P`  E  De @Te @ V                     FP                           !     P  R  `  @   @                   ffSffe0vffcGfffDvff�GffDDFf���v e   V 0  S e4P fg` fgCffE3FP de  V                       De  VDF             @ B   @ P@  dDDD E e   V             DDDD                     DDDD        ffFevfFfDvGf�GtfDDtf��DvDDDD����3  e3  fe30ffeSffffffffvfffDvff         0   S3 fe33fffeffff T      $         340 fde3                    29�ws��w7y��wwGw��w��G}��w���wDDvf���vDDDD����DDDD����DDDD����ffffffffvfff�GffDDDv����DDDD����ffFfffFfffFfffFfgDFfDDFfDDDvDDDNfU33ffffffffffffffffffgDfftDDGDD3333ffffffffffffffffvfffGfffDfff3333ffffffffffffffffftGvgDDGtDDD4333dfffdfffdfffdfffdfffdfffdfff4333dfffdfffdfffdfffDvffDGffDDff3333ffffffffffffffffftGfgDDGtDDG3333fffffffffffffffffffgffftffgD3333ffffffffffffffffGfffDGffDDvfDDDD����DDDD����DDDDDDDDDDDDDDDDDDDD����DDDD���DDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDDDDDDDDDDDDDDDDDDDDDD�DD�DDDDDDDNDDDDDDDDDDDDDDDDDDDD��DDDDDD�DDDDDDDDDDDDDDDDDDDDDDDDN��DDDDDN�DDDDDDDDDDDDDDDDDDDDD���DDDDD���DDDDDDDDDDDDDDDDDDDDDDDN�DDDDDDD�DDDDDDDDDDDDDDDD"""3334DD4DD4DD4G4q3""""3333DDDDDDDD""""3DD3wwww""""3333DDDDDDDD4DDD"7DG2#tG""""3333DD""G3Dq3|U#7|w#w|�""""3333""4DD3"7\w2#C�C2\wt3""""3333DDDDDDDDtDDDtDGtDq3"""'3337DDD7DDD74DD7"7D72#t77#77#w73w7Cw7s77t34wC4wwwL�wt�<w|U\W�wwEwwwGDwtC3333C32"C2tGt3wGw3wGs3wG34tD3'tD"GtDGwDD3w|wCw|�s7wwt3DwwC33wwC3GwwwDGwwC�w3\wt3wwC4tC3'33"G2"GwwwwtwwwDtG#7tG#wtG3wtGCwtGs7DGt3DDwCDDwwt�\Guwwwuwww|DDww�\GDwtC3333C32"C2t7t3t7w3t7t3t7C4t73't7"GD7GwD74Gw4DG4DD7ww7ww7ww7ww7t2DDDDDDDD����DDDDDDDDDDDD�dDDSNvDN��N�������DDDDDDDDDDDD�nDDSDDDDDDDDDDDDDDwwwwws!wws!wws!wws!wDDDDDDDDDDDDwwwwC4wwB"GwA#GA4���D��������DDDDDDDDDDDDDDDDDDDDwwwwwwwwDDDDwwwwC4wwB"GwA#GA4DN�tN��t���tDDDtDDDtDDDtDDDtDDDt3!7t27ww7ww7ww7ww333wwwe1SNv�dDDDDDDDDDDDDDDwwwwDDDDDDSDD�nDDDDDDDDDDDDDDwwwwDDDDws!wws!wws!wws!wws"wwwww3333wwwwA#A4A#GB"GwC4wwwwww3333wwww�DDDDDDDDDDDDDDDDDDDDDDDwwwwDDDD�DDtDDDtDDDtDDDtDDDtDDDtwwwtDDDD  �  �  �  �  �  	�  	�  � �  �  �  ��  ��  ��  ۰  ۰  ۰  ��  ��  �� �� �� �� �  �  �  �  �  ��  ��  ��  ��    P                             EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDFDDDDDDDDDDDDDDDDDDDDDDDDDDfffffffffffffffdffdDffdffdFffdffDDDDDDDDDDDDDDTDDDEDDDEDDDDDDDDDUUUUU"RUU""UUR"UUU"%URUUU"UUUUUU""""""""$D"""DD"""B"""B"""B"""""DDDDDDDDDDDDDDUTDDTTDDUDDDDDDDDDUUUUUUUUUwuUUuuUUwuUUWuUUUwuUUUUwwwwvgwwvvgwvwfwwwvwwwwwwwwwwwwwffffffffffffffffffffffDfffFfffFfDDDDDDDDDDDDDffDDDFdDDDdDDDDDDDDfffffgfffgwffffvfffwffffffffffffwwwwwwwwwwgwwwgwwwvwwwvgwwwgwwwwffffffffff�fff�fff��fff�fffhffff�����������������������x���w����                                                  �  � y� ���         ���i���}���������������    �������������������            {  �y�  ˙` ̹� ��i`                                                           	���}���l|���̛��̜�ww�����������qqA}����}q���̙��w���w}w���������w��͝��yq�|�qk}�����ww�    �   {   �     � qy� ��     	   	     �     s�ww���͜���}���}��ww����t��twwwww}q�q|����qwqw}ww���q|����{��wiyww|��{  ِ  y`  ��  �   �   �        ww                            wy�� ��  ��   y              ������������{��̙v��י�  �y    �������������������i���v�w�     �̹p�͙ �ٛ ٗ  ��                   �      �                   wwwtwwwCwwt1wwCwt1wCt1��C��1�����������""""�����������!�����!""���������Gw�7w�w���G���7����������wwwwwwwwwwwwwwwwwwwwwwwwGwww'www1���s�wC�t1��C��1���1���1���$��"G�$ww�������������������!,���������!w��www!��wq��wr�ww!�wwq�wwwwww!wwwrwww�Gww�'ww�ww��Gw��w��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDDD3333;���;���;���;���7wwwDDDDDDDD3333����������������wwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333=���=���=���=���7wwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333���G���G���G���GwwwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333<���<���<���<���7wwwDDDDDDDD3333��DG��DG��DG��DGwwwwDDDDDDDD3333�DDG�DDG�DDG�DDGwwwwDDDDDDDD3333DDDGDDDGDDDGDDDGwwwwDDDDwwwwUUWUUWUUWUUW333wwwwwwwwUUwUUwUUwUUw333wwwwwwwwfgwfgwfgwfgw333wwwwwwww�ww�ww�ww�ww333wwwwwwww�ww�ww�ww�ww333wwwwwwwwwwwwwwwwwwww333wwwwDDDD33334DDD4DDD4DDD4DDD7wwwDDDD                         d  eU  Fff t�G �� �D�CG��}������������~���ww�ww�w�I���t�y�t�y�t�y�                                                        w   �   �   �   w   w   w   w   w   w                         f@ UP ff O� �� �� �t4���������}���}}��w}��wywyt���w���t�w�t�y�t�y�                            `   p   @   @   p   ��  ��  �p  wp  wp  wp  wp  wp  w   w   w   w             �� �� �� �w �& wv	�wp�� ɪ��̙�������̰��ɰ����ک��؋�H���TZ�REDZ�4DJ 4D          P c c 1 61   11� 1   61 c 1 P c                 ` P 0c` 65    6  �5 6    65  0` ` P             ��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwtD   �   �   �   w   G   G   D@  D@  f^� fO� wp  wp  �p  ��  ��      �   "   "   R   �D  J�  D�  ��  ��  "   ""  """              �p  �G  ��  ��  ��  �O@ tG� 3##�""37##4pCCwpDGww3Gww��ww��ww w  ww  vdw eUw FVg fd��G��w�����������w}}w}}ww�}www~I�D�t�y�    �@  ��  ��  ��  ��  �O  wp�3##�""37##4pCCwpDGww3Gww��ww��ww��tD}�t}�DN}wtOwwtTwwfewtfewFFVwFDewUgFwI�wwI�wwt��wwy�wwwIwwwt t���{���{���t�G����t�G��w{{���{���w���wt��ww��ww�Gwwtww�Gtw���         �  �� �  ��  �p  �p  �p  wp  �p  �p  wp  wp  wp  Dp         t�O��0� �#G27D3"# t32 wD3 wwC wwt wwt ww ww tG tDDt�G��ww��wtTwwfeGtfegvfT@FFVFFDfVUgFdI�wwI���t���wwwI       t �O �� 4� /� #G 3D t3# t32 wD3 wwC wwt wwt ww ww       O  �  �  �  �  wN ww ts� w2� s"7 s#w s7t wwt ww ww         ww C4p4�pwO�pww�pwH�~t���t���t��wwwDwws3GwCCGw4C7t4t7    7   C~� �p �G` �v` ufp fgp Fwp gwp �wp wwp ww  �G  tG  �           ww C4p4�~wO�yww�ywH��t��t���t�wwwwDwws3GwCCGw4C7t4t7 �� .�� �/	��y��w���w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww            C9  OI  ��p �pw�wt�G wIGwwyGwD�GsDDwDwwwGtDwwwww O�@�����G���O�����Op��wp�B4p�!"pr20Cr#@4r3"72"3443GCwwwwG}� �p �����#�������y�w������������w�y�y�ww�Gwwwwt33Dt343    40� DC� �CV ��V �Ef �E` ffp fgp fwp fgp fgp wGp D�p �p t�p            � C9� 4� O� w� wI�pt�Gpt�w t�wwt�DwwDD7wwwDwDGtwwww �� ��2������������y������w���w�y�y�ww��wy�Gwwwwt33Dt343    40  DCp �Cp ��p �D  ��  f�` ge` gfP fv` fwp wGp D�p �p t�p   �� �� q����y�����w���wy�������y���w��ywwwwwwwwwwwwwwwwwwww  �� �� � ���	��𙈉 ���y�������wy�yww��wwwwwwwwwwwwwwwwwwww             C4  4� O� w�wHw�t���t�� t�wwt�DwwDD7wwwDwDGtwwww�$pq3#pB#3p237p2#ww42"�Gt3wG}�                    �p  �p  wp   O�@�����G���O�����Op��wp�B4p            �  ~�  7p  7   p     �  �  �  �  w  w  w  t����ﻻ���K�{�{�t�{�wG~�Gt��y�wvfT@FFVFFDfVUgFdI�wwI���t���wwwID�  W�  g   wp  wp  �p  ��  ��         O  �  �  �  �  wN ww    �p  �G  ��  ��  ��  �O@ tG�  wwpwvVwfewwvfww��w���}������w    p   g   w   g               �� .�� �/	��y��w���w���wy���    �   �   �   �   �   �         �� �� q����y�����w���wy���                        �      �!"pr20Cr#@4r3"72"3443GCwwwwG}�        ��  ?�  Gp  wp  wp  wp  �G O�' t���ww�ww��w}�w��wp���p����ﻻ�wt��ww��ww�Gwwtww�Gtw��� Dp GGG GG��w��G}��w���w���w            �  ~�  gp  g   p             ~� u~�vV` Vfp fp  w       �   �   �   �   �   �                 ~� |~�}�� ��p �p  w             ~� z~�{�� ��p �p  w           ��  ?�  Gp  wp  wp  wp            ~� r~�s#0 "3p 3p  w    �  ~� #p #  r7  #p  7p  w    �  ~� �p �  }�  �p  �p  w    �  ~� �p 
�  {�  �p  �p  w               �  ~�  7p  7   p               �  ~�  �p  �   p   ��  y�  y�  wp  wp  wp  wp  Dp   �t v w~ ww  ww  t  tG  �                �  ��  �   �               �  ~�  �p  �   p        DD t� G��w�w27�w3$ws2w                        �         �  �  �  w  &  v  �w 
�� ��� �˙���
�������ۼ̻��"� �"% 2"#                        �   �   �   {   '   v   j�  ��� ��� ��� �˹ ̽���ة�����˰����,�T"+ 3"%                         7v` weV "fff"O�p"��p"��p"�p3�}p-��p=��p|� }�  }�  ��  ��  ��  ��  �  �  �  �  �  "              `  eV  fff O�  ��  ��  �  �} �� �� ��  |�  }�  ��    =   }   =   =              �������}�}�}�ww~r�� ∈�������������������}�� }�� ��� ��� ����   �   �   �   �   �   �   �   C""42""#2""#2""#2""#s3342"""3333    p   p   p   p   p   p   p    ��������� ��� }�� ��  ��  ����  ��  ��  ��  ��  ��  ��  ��                          � �� ��    "               wvf wfU 7Of`w��f"�� "�p-�}p���� ��� ����x��	�� �� �� "�        f  U` f` f` �p w���� `  eV  ff  O�  ��  �� ����}�                �  �  ��  �            �  �  �   �  ��  �                     �  �  �   � `  eV  ff  O�  ��  ��  ����}���������������p	���         `  eV  ff  O�  ��  ��  ���}�     �  �  �   �  ��  �   �            ��  ��  �   ��  �   ���������������p	���                    3333UUUU                        wwww                    333333333333333333333   w  G� ws@ ws� ws$7w@wwww"                               ����������� ��� �� ��  �    `  eV  ff  O�  ��  ��  � ��}�            """"                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	   �  	   �  	   �  	   �   ����                                             	�  �	 	  ��  	                                �  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	���                �   	    �   	    �   	    �   	����                                                               
   �  
   �  
   �  
   �   ����                                             
�  �
 
  ��  
                                �  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
���                �   
    �   
    �   
    �   
����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "                "  !"!" "                      ��   �                  �  �  �� �               �  �  �ݻ���������2��������ݻݻ� ��                             "                "  !"!" "                ����	�   	�   	�   	   �  	�  �  	�  �  	�	����    �  	�  �  	� ��              �              � 	����  �            " ""   """! "   "      ""  "!  "       " ""                 ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                     P  U  UePVfUUUU        UP  VeP VfUPVeP UP                                                                                                                                                                                      ����
�   
�   
�   
   �  
�  �  
�  �  
�
����    �  
�  �  
� ��              �              � 
����  �                                                                                                                       �����   �   �      �  �  �  �  �  �����    �  �  �  � ��              �              � ����  �                                                                                                                                                                        �w
���̩ۚ,���+��   �   �   �   �  �  9  D3  D2 T2 DB DB �@ ��  ��  ��  �  "" ""�"!��" ��       �                w�  ��� ��� ��� ˼����ɀ�؊�˽ـ��˰��̰�̻@"���"+H�"$X�"$�@"E� U� E� D� ,˸  ��  ��  ,� "" �"" """�"!���� � �              �         �           �       �                                      "  ."  �"    �          �� ̻� ��� ww� ��� vvw    �   �     �     �  �  �   ��  �   ��  �                �"�!/"�  �                                                                                                                                                                                  "  " �" ��" ��- �ۼ w۽��ݹ����� ��� ��  ˼  ��  ˼  ��  H�  �D  J�  J�  �  �  �  �  
�  �  �  �  ,�  " "" �" �"�   ˰  ��  wp ��ډ�v���r�̸��˰��� ��  ��  ��  ��  ̸  ��  ��  DC  C4@ T4@ T40 T30 T30 S;� H�  ��  ��  ��  ""  "  �""� "�/��        �   �   �      �  �   �   �   �   �              �   �   �   �             ���� �                        " "" """ �"  �   �   �                              � ��                  �  �˰ ��� �wp ���                                                                                                                                                                                  0  �0 ! ..0   �  �  �  b  g   w   
   �   �   �  �  �  	�  
�  	�  �  ̽  ̴ �% ""X ."� �%� �H � 	�� �� �  " """""�  ���   �   �   }   g�� z�� ������ˀ���л�����̰��� ��� ۼ������۸�@���0X�S0�E3 �X� EJ� D+  �"/ �" ����� �  �  � �   ��  �                       �  � ���� ��� ��                      "   "   "  �� ��                   ����������                                �   ���                            "  "  "                                                                                                                                                                    �  ��� ݻ� g�� bm� ggz�'w���������������˛������ˊۼ�����˻������H�DH�@U�DPT�E X�T H�P H�@ Ȥ� ̻� ˘ "�� � ���/�"" �""/���               �   �                                                     �  �                      � �                       ���           �                      �  �  �          ����  �   �             ����                         � "            � "�",�"+� ",                       "  .���"    �     �                     �   �   �  �  �  �     �   �   �   �   �  �  �  ��  �      �   �  �� ���������� �                                                                                    �  �  ��  8�  5I  5U  3U  DT  EZ UJ T� �J� ����+�""""�""//��          ��wɪ�pɪ��ɪ��̙�н��н̽Ѝɚݣ��"�<̲�;���0"�0  ="  ""  "/  /�� ���  �����                               �� �� �� ���          �.���       �  �      �  ��  �  ��  �              �                                   ����  �   �             ����                         � "            � "�",�"+� ",                       "  .���"    �     �                                                                                                                                                                                                            �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                   �   �   ��   ��  �   ��   �                                                                                 �  �  ��  �                                                                    	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  T   C   30  =�  ݰ  ۚ  �  
�� ���  +"  "" ���������                   �                        ���� ��� ����                            ��� ���� ��             �  �˰ ��� �wp ���                                                                                                                                                                 	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��    "  "  "                  �� ��� ��                      "   "   "  �� ��                   ����������                �  �  ��  �   �   �        �  �  �   �   ��  �                            �   ���                            �   �                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                        �          �   � � �  ��� ��  �    "   "   "  �� ��                   ����������                          �  �� ��  �    � ���                                                                                                                                                                                             ���
̻���������ܽz�w� ݸ� ���    �   ��  ��  �̰ �̼ �̻ ��˰"�� �����빚�̻�H��4T�EU UU EUU EUU DTT D@ ˰ 	�� 
�� �  "  ""/""�"/������  ��    �ܻ �۸ ����ܙ:0�38�D33�DC3�TD38@338 3;  �"  "   "   �  � �� � �����    ��                          "   "/  "/� ��  ��                   ""  ."  �"    �   ��  �   �                  �  �  �  �                                       �  �   ��                     �    � �  ��                  ���                              �   ���                            �   �                                                                                                   	�  ɪ� ��� ��� ��� ��� ��� �� ��  "( "" "" B. DN TN UN �� 	�� ڙ� ����� " "� � ���   �                        ��  ��  �̰ �۰ g}� �ת�vw��gx����������3ؼ�D:��I�� ̚P+��P",UP"%U�"�� �� ۰ -   " �" �������� � �   �   �   �   �   �   �   �   �   ��  ��  ��  ��                  Ͱ  ˻  ˻  ۻ  ݻ  ��  ��� ��� ��˰��˰̼˚̽��                                                 �    ���  ��                    ��  ��  ��� ���                                                                                                                                                                                                                     �  �� �� ɪ� ������	��͈��ݙ�3C���3���ع����غ��٫��뺛�ɾ谹���������  �   �                       ��  ��  ̻� ������ڌ))ڌ����������ɛ��ݻ34C0��=���ۍ�ٻ����� �� �� ��  Ⱥ  ɫ  ��  ������������������������        �   �   ��  ��  ��������
��� ������� ���   �   ��  ��  ��  ��  �� �  �           �                    �          �         �   �  �  �   �               �   �                                                                                                                                                                                                                            �  0  � 
0 � : 1 ww 1s p 1q�u1uU �������:0wwwwUUUU��������wwwwUUUU :p �p�p�p
0p
p
0p�p�7p �p :7p 
p �p                                                                                                                  ww   � 0 � 0 � p  q  q  q  q 1q�0�0�0�
 � 
  ��    wwww00����
�������    wwww��������








����                                                                                                                                                                                    D@ D�D D@                     �� ������ 0	�� � ���� ���0	��� ��Ð ��9 
	�
 �� 
�  

              �      �      �      
                                                                                                                                                                                                                                                                                                                                                                                                                                              "" #3 #w #w            """"3333wwwwwwww             ""0 34p w4p w4p  #w #w #w #w #w #w #w #wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww4p w4p w4p w4p w4p w4p w4p w4p  #w #w #3 $D 7w            wwwwwwww3333DDDDwwww            w4p w4p 34p DDp wwp             DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4344DCDCDCDD4CD3DCDDDDDDDDDDDDD443D344434444444443DDDDDDDDDDDDD3D3D44443D444444443DDDDDDDDDDDDDDDDD34DD4CDD4CCD34CC4DCC4DC4DDDDDDDDDDDDDDDDCC3DCCCDCC4D3CCDDDDDDDDD34CD4CCD4CCD34CC4DCC4DCCDDDDDDDDDDDDDDDD3D44D44434CDD4CDDDDDD3DDD3DDD3DDD3DDDDDDD3DDD3DDDDDDC43DC43DCD4DD4CDDDDDDDDDDDDDDDDDDDDDD44DC33DD44DC33DD44DDDDDDDDDC33D4DD4434444D443444DD4C33DDDDD3DCD3D3DDC4DD3DDC4DD3D3D4D3DDDDDD3DDD3DDDCDDD4DDDDDDDDDDDDDDDDDDDCDDD34DC33D3334DCDDDCDDDCDDDDDDDCDDDCDDDCDD3334C33DD34DDCDDDDDDDDDDDDD4DDC4DD3D4C4D33DDC4DDDDDDDDDDD3DDD3DD333DD3DDD3DDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDD4DDCDDDDDDDDDDDDDD333DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC4DDC4DDDCDDD3DDC4DD3DDC4DD3DDD4DDDDDDDC33D3DC43DC43DC43DC43DC4C33DDDDDDC4DD34DDC4DDC4DDC4DDC4DD33DDDDDC33D3DC4DDC4DC3DC3DD3DDD3334DDDDC33D4DC4DDC4D33DDDC44DC4C33DDDDDDC3DD33DC43D3D3D3334DD3DDC34DDDD33343DDD333DDDC4DDC43DC4C33DDDDDC33D3DD43DDD333D3DC43DC4C33DDDDD33343DC4DD3DDC4DD3DDD3DDC34DDDDDC33D3DC43DC4C33D3DC43DC4C33DDDDDC33D3DC43DC4C334DDC44DC4C33DDDDDDDDDDD4DDDDDDDDDDDDDDD4DDDDDDDDDDDDDDDDDDC4DDDDDDC4DDC4DDD4DDCDDDDDD33343334DDDDDDDDDDDDDDDDDDDDDDDDDDDD334DDDDD334DDDDDDDDDDDDDC34D4D3DDD3DD34DD3DDDDDDD3DDDDDDD34DCDCDC3CDCCCDC34DCDDDD34DDDDDD34DD34DD44DC43DC33D3DC43DC4DDDD333DC4C4C4C4C33DC4C4C4C4333DDDDDC33D3DC43DDD3DDD3DDD3DC4C33DDDDD333DC4C4C4C4C4C4C4C4C4C4333DDDDD3334C4D4C4DDC34DC4DDC4D43334DDDD3334C4D4C4DDC34DC4DDC4DD33DDDDDDC33D3DC43DDD3D343DC43DC4C33DDDDD3DC43DC43DC433343DC43DC43DC4DDDDD33DDC4DDC4DDC4DDC4DDC4DD33DDDDDDC34DD3DDD3DDD3D3D3D3D3DC34DDDDD34C4C43DC34DC3DDC34DC43D34C4DDDD33DDC4DDC4DDC4DDC4DDC4D43334DDDD3DC4343433343CC43DC43DC43DC4DDDD3DC434C434C43CC43D343D343DC4DDDD333DC4C4C4C4C33DC4DDC4DD33DDDDDDC33D3DC43DC43DC43CC43D3DC333DDDD333DC4C4C4C4C33DC4C4C4C434C4DDDDC33D3DC43DDDC33DDDC43DC4C33DDDDD33334C4CDC4DDC4DDC4DDC4DD33DDDDDC4C4C4C4C4C4C4C4C4C4C4C4D33DDDDD3DC43DC4CDCDC43DC43DD44DD34DDDDD3DC43DC43DC43CC4333434343DC4DDDD3DC43DC4C43DD34DC43D3DC43DC4DDDD3DD33DD3C4C4D33DDC4DDC4DD33DDDDD33344DC4DD3DDC4DD3DDC4D43334DDDDDCDDD3DDC3DD3334C3DDD3DDDCDDDDDDDCDDDC4DDC3D3334DC3DDC4DDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDC334DDDDDDDDDDDDC34DDD3DC33D3D3DC334DDDD3DDD3DDD334D3D3D3D3D3D3D334DDDDDDDDDDDDDC34D3D3D3DDD3D3DC34DDDDDDD3DDD3DC33D3D3D3D3D3D3DC334DDDDDDDDDDDDC34D3DCD333D3DDDC33DDDDDD34DC4DDC4DD33DDC4DDC4DD33DDDDDDDDDDDDDDC3343D3D3D3DC33DDD3DC34D3DDD3DDD334D3D3D3D3D3D3D3D3DDDDDD3DDDDDDC3DDD3DDD3DDD3DDC34DDDDDDD3DDDDDDD3DDD3DDD3DDD3D3D3DC34D3DDD3DDD3D3D3C4D33DD3C4D3D3DDDDDC3DDD3DDD3DDD3DDD3DDD3DDC34DDDDDDDDDDDDD343D3C443C443C443C44DDDDDDDDDDDD333DC4C4C4C4C4C4C4C4DDDDDDDDDDDDC34D3D3D3D3D3D3DC34DDDDDDDDDDDDD334D3D3D3D3D334D3DDD3DDDDDDDDDDDC3343D3D3D3DC33DDD3DDD3DDDDDDDDDC3C4D34DD3DDD3DDC34DDDDDDDDDDDDDC33D3DDDC34DDD3D334DDDDDDDDDD3DDC33DD3DDD3DDD3DDDC3DDDDDDDDDDDDD3D3D3D3D3D3D3D3DC334DDDDDDDDDDDD3D3D3D3D3D3DC34DD3DDDDDDDDDDDDDD3C443C443C443C44C4CDDDDDDDDDDDDD3DC4C43DD34DC43D3DC4DDDDDDDDDDDD3D3D3D3D3D3DC33DDD3DD34DDDDDDDDD333DDC4DD3DDC4DD333DDDDDDD4DDCDDDCDDD4DDDCDDDCDDDD4DDDDDD4DDDCDDDCDDDD4DDCDDDCDDD4DDDDDDwwwwwtDDwAt!""t��B�DA�DAwwwwDDww(Gw"�w��wD(GD(G(GwwwwDDDDAAA��A�DA�DAwwwwDDGw�w(G�(GD(GD(G�GwwwwwwDDwDt�"H�A$DAGwAGwwwwwDDGw$w"""G���GDDDwwwwwwwwwwwwwDDDDAA""A��A�DA�wA�wwwwwDDGw(Dw!�G��GD(Gt(Gt(GwwwwDDDDAA""A��A�DAA""wwwwDDGw�w""(G���GDDDG�w""�wwwwwwwDDwDt�"H(�A�DAGwAGtwwwwDDGw�w""(G���GDDDGwwwwDDDwwwwwDDGwA�wA�wA�wA�DAAwwwwtDGwt$wt(Gt(GD(G(G(GwwwwtDDwA(GB(GH�GH�wH�wH�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGwwwwwtDDwt(Gt(Gt(Gt(Gt(Gt(GwwwwDDGwA�wA�wA�tA�AAAwwwwwDDwt(GA(G�G(Dw�wwGwwwwwwDDGwA�wA�wA�wA�wA�wA�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwDDGDA�AA!A�A�A�wwwwGDGw��w(GG(AG(AG(AGwwwwDDwwAGwAwAGAAA�wwwwtDDwt(Gt(Gt(Gt(GD(G(GwwwwwDDDtB""A��A�DA�wA�wwwwwDDGw�w"(G�(GD(Gt(Gt(GwwwwDDDDAA""A��A�DA�DAwwwwDDGw�w"(G�(GD(GD(G(GwwwwDDGw�w"(G�(GD(GD(G�GwwwwwDDDtA"""A(��A(DDAB"""wwwwDDGw$w""(G���GDDDwGw"$wwwwwtDDDAB""H��tDDwwtwwtwwwwDDDw(G""(G(��G(DDw(Gww(GwwwwwwtDGwA�wA�wA�wA�wA�wA�wwwwwwtDwt(Gt(Gt(Gt(Gt(Gt(GwwwwwDDwt�(Gt�(Gt�(Gt�(Gt�(Gt�(GwwwwDDGDA(DA(HA(HA(HA(HA(HwwwwGDDw�A(G��(G��(G��(G��(G��(GwwwwtDwwA(GwA�wA(Gt�wAwtwwwwwtDwwAGtGA(G�w(Gw�wwwwwwtDGwA�wA�wA�wA�wA(Gt�wwwwwDDwt(Gt(Gt(Gt(GA(G�wwwwwtDDDAB"""H���tDDDwwtAwwAwwwwDDDw(G"!(G�(G�w(Gw(�wwwwwwwtDDwH!t�t!(�H�DH�wH�wwwwwDDww(Gw�w�$wD�(Gt�(Gt�(GwwwwtDDwA(GA(Gt(Gt(Gt(Gt(GwwwwDDDDAB"""H���tDDDtA"""wwwwDDGw$w"!(G��(GDA(G(G""(GwwwwtDDDAB"""H���tDDDwAwB""wwwwDDGww"(G�!(GD�(G�G"�wwwwwtDGwA�tA�tA�tA�tA�tAwwwwDGww�ww(Gw(Gw(Gw(Dw(GwwwwDDDDAA""A��ADDAB"""wwwwDDDw(G""(G���GDDDw�w"!(GwwwwwtDDwBt!"t(�B�DBB""wwwwDDGww""(G���GDDDw(Gw""�wwwwwDDDDAB"""H���DDDDwwwwwwwwwwwwDDDw(G"(G�(GD(Gt(GH�wwwwwwDDDtB""B��BDDHt""wwwwDDGw�w"!(G��(GDA(G�G""�wwwwwwDDDt!A""A(��A(DDA(DDAwwwwDDwwGw"�w��$wD�(GD�(G(GwwwwwDDwt(Gt(Gt(Gt(Gt(Gt(GA""A��A�DA�wA�wH��wtDGwwwww"(G�(GD(Gt(Gt(Gt��GtDDwwwwwA��A�DA�DAAH���DDDDwwww��GD(GD(G(G�G���wDDGwwwwwAGwAGwH$DHt�""wD��wwDDwwwwwwwwwwwwDDDwG""(G���wDDGwwwwwA�wA�wA�DAA"""H���DDDDwwwwt(Gt(GD(G�G""�G��DwDDGwwwwwA��A�DA�DAA"""H���DDDDwwww��GwDDwwDDDw(G""(G���wDDGwwwwwA��A�DA�wA�wB"�wH��wDDGwwwww��GwDDwwwwwwwwwwwwwwwwwwwwwwwwwwAGtAGtB$DHt�""wD��wwDDwwww�(G�(G�(G(G""(G���wDDGwwwwwA�DA�wA�wA�wB"�wH��wDDGwwwwwD(Gt(Gt(Gt(Gt"(Gt��wtDGwwwwwH�wH�wH�wA(GB"(GH��GtDDwwwwwA�wA�wA�DAB"""H���DDDDwwwwt(Gt(GD(G(G""(G���wDDGwwwwwAA��A�DA�wB"�wH��wDDGwwwww�ww(Dw!�GB(Gt"(Gt��GwDDwwwwwwwwwwwwwDDDw(G""(G���wDDGwwwwwA�A�A�A�B"�"H���DDGDwwww(AG(AG(AG(AG(B(G�H�GGDDwwwwwA�!A��A�HA�tB"�wH��wDDGwwwww(G(G!(G�(GH"(Gt��wwDGwwwwwA�wA�wA�DBB"""t���wDDDwwwwt(Gt(GD(G(G""�G���wDDGwwwwwA""A��A�DA�wB"�wH�GwDDwwwwww""�w��GwDDwwwwwwwwwwwwwwwwwwwwwwA""A��A�DA�wB"�wH��wDDGwwwww!�w�GwA$wA(GB"(GH��GDDDwwwwwt���wDDDtDDDAB"""H���tDDDwwww�!(GD�(G�!(G(G""�w��GwDDwwwwwwwwtwwtwwtwwtwwt"wwt�wwtDwwww(Gww(Gww(Gww(Gww(Gww�GwwDwwwwwwwA�wA�wA�DAB"""H���tDDDwwwwA�wA(Gt�wAwt""wwH�wwtDwwwwt�(GH!(G��w(Gw"�ww�GwwDwwwwwwwA(HA(HA(HBH"""t���wDGDwwww��(G��(G��(G(G""�G���wGDGwwwwwwtwAt�A(GB"�wH�GwtDwwwwww�ww(Gw�wA(Gt"(GwH�GwtDwwwwwwAwtwwAwwAwwAwwB(wwtDwwww(Gw"�ww�Gww�www�www�wwwGwwwwwwwwDt��H!�AB"""H���tDDDwwww�Gww�wwwDDDw(G""(G���wDDGwwwwwH�wH�wH(Dt!t�""wH��wtDDwwwwt�(Gt�(GH(G$w""�w��GwDDwwwwwwt(Gt(Gt(Gt(Gt"(Gt��GtDDwwwwwA(��A$DDA$DDAB"""H���DDDDwwww���wDDGwDDDw(G""(G���GDDDwwwwwwH��wtDDtDDDAB"""H���tDDDwwww�!GD�(GH!(G(G""(G���wDDGwwwwwB"""H���tDDDwwwtwwwtwwwtwwwwwwww(G(DG(Gw(Gw"(Gw��wwDGwwwwwwH���tDDDtDDDAB"""H���tDDDwwww��(GDA(GDA(G$w""�w��GwDDwwwwwwB��B�DBDtt�""wH��wtDDwwww��(GDA(GDA(G(G""�w��GwDDwwwwwwwwwwwwwtwwwAwwt�wwt"wwt�wwwDwwwwA�w(Gw�ww(Gww(Gww�wwwGwwwwwwwH��BDDBDDBH"""t���wDDDwwww��(GDA(GDA(G(G""�G���wDDGwwwwwH"""t���tDDDt�t�""wH��wtDDwwww"(G�!(GD�(G$w""�w��GwDDwwwwwwt(GwDDwwDDwt(Gt"(Gt��GwDDwwwww"""������������������""""���������������������""""������II������""""������IIII""""������DI�I�""""������DI�I�""""�����IIDIIIA""""��������DD""""������IADD�A��""""��������I���I�������I���"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD���4���4���4���4���4���43334DDDD"""������������������""""������������������������""""����������""""��������AD�I�""""��������AA�A�""""��������AI�I�""""����DD�I�""""��������DD""""�������IAA�I�""""�������������A��A��"""$���4���4���4���4���4���4������������������333DDD������������������������3333DDDD��������D�D�����3333DDDDM����D��D����3333DDDDA�A�A�D��M�D�����3333DDDDM�M�M�M��M�D����3333DDDD��A�M�M���M�����3333DDDDMDD�����D��D����3333DDDD��D��A�MD������3333DDDDA��A��A�AMMDDM����3333DDDD���4���4���4���4���4���43334DDDD                                333UUUTDDTDDVfwVfwVww3333UUUUDDDDDDDDffvfvgwfwwww3333UUUUDDDDDDDDffffwvffwvgv3333UUUUDDDDDDDDffvffgwvfwww3333UUUUDDDDDDDDgvffgwfwvwgw3333UUUUDDDDDDDDfvfdgwvdvgwd3334UUU�DDG�DDG�ffg�fwg�gww�WwvWwvWw�Wn�V~�Vw�W~�W��wwfwwwwwwwgvvwwwwwwfwwv~wgw��v~�wwgvg�vw~��g~��w~�ww���g���v����wwwwwwgwwvwvww~wwg��w�D�~DDNdDJDvwwww�ww~��f~��ww�wv~��w��������vgwtwwwtw�wt~��~~��~w�v~~��~���~www�gvg�fwg�g�w�~���~���w�w�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUCT���^���^���U���T���TJ�DEDDDCEDuUUUUUUUUUUUUUUUUUUUUEUUUTUUUEEUUUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUUWUUW�UUW�UUW�UUW�UUW�UUW�UUW�UUW�UUUUUU\��\��\��VffX��X��UUUUUUUU������������ffff��������UUUCUUT4���4�����CCffCE���4���Sqrrr!qr'qr'qq'qqq'qqqrqqqrqqqrCEUUCCUUT4\�44\�44<�CCFf�CH��4��UUUWUUUW������������ffff��������UUW�UUW�������������ffg䈈�䈈��R""R""R""R""R""R""R""R"""""""""""""""""""""""""""""""""""#S"%CC"'EC"$GC")D4"��4"��4"��TqqqrqqqsrqrtGDtqwwwwwwwwwwwwwwwt"T4""T""CE""EG""GD""$I""*��R*��/�"%"�"%"�"#"-"#"/"#"/�"""�"""�"""'�""'�""'�""'�""'�""'�""'�""'�"�"t"""�"""D"""D"""D"""D"""D"""DDDDNN�DDDNDDDGDDDCDDDCDDD�DDD�DDr*���"*�B"""B"""B"""B"""B"""B"""""�"""-�""/�"""�"""�"""-"""-"""/""'�""'�""'�""'�""'��"'��"'��"'�"""D"""N"""D"""D"""�"""�"""t"""~NsDD��DN�CN�NCDDDC�DDC�DDCtDDC~DB"""�"""r"""�"""B"""B"""B"""B"""�"'��"'���'�-�'�-�'�/�'�"�'�"���R""R""R""R""R""Www���DDD""""""""""""""""""""wwww����DDDD"""w"""D"".D""tD"%DNwwww����DDDDDCwDDCDDNSD��'DD"TDGwwww����DDDDB"""B"""B"""R"""""""wwww����DDDD"���"-��"-��"/��""��www�����DDDDUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUTSUUT4UUT4��CC��44�ECEfdTS��43��43!rrr!qr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44S�444�CCFf�ECH�5CH"CCC"%EC"$DC""��""��""��""��""*TCCCECCCGECEJ��N�DDJ�DDI�DDD�DDDN"ECB$T4"ECB"DT""�r""�"""�"""R""""""t"""�"""D"""D"""D"""D"""D"""Dr"""�"""B"""B"""B"""B"""B"""B"""UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUC���4��TT��CEffCE��E4���C44TTCEEC4CCE�EEI��I��DD�DE3D5DD54UUUCEUUEL�̤4�̤4��EFff5H��D���"""D"""E"""E"""N"""$"""$"""$"""Tw#swrqrsqqqrrrrtGttwwwwwwwwwwwwtR"""B"""B"""B"""""""""""""""R"""wq3wwqwwt!wGGwwq'ws3333DDDDwwwwUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUY�UUUUUUUUUUUUUUUUUUUUUUUUUUUE�UUEUUY�UUY���̚��������ffff���������UTT�UCEED4UDSCEED4UdSEE�D�C����qrrrqqr'qqr'qqq'qqq'qqqrqqqrqqqrCEUUCEUUT4\�44\�44<�CCFf�CH��44�"""#"""%"""%"""""""$"""$"""$"""T"T4""T3""CE""EG""GD""$I""*��R*��DDDNN�DDDNDDDGDDDBDDDBDDD�DDD�DDNrDD��DN�BN�NBDDDB�DDB�DDBtDDB~DDBwDDBDDNRD��'DD"TDGwwww����DDDD3333UUUUDDDDDDDDffvjvgw�www�3333UUUUDDDDDDDD�fff�vff�vgvwwf�www�wwgzvwwtwwwewwvtwgw��v~�wgv��vwD��gE��wENwwT^�gT^�v4^��43UUCCEUCCEUE44UTT4UUECCUTT5UT5EUUCTUUTU���E���E���EfffE���C����CEUUCEUUT4\�44\�44��CCFf�CH��44�"""#"""%"""%"""#"""$"""$"""$"""TUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUCT���^���^���U���T�J�D�IDT��DE��wUUTtUUED��D3��5D��D3fffV��������'Qrwq7'ws'ssr'rq'rqqrrqqrqqqrCCUUCCUUT4\�44<�444�CCCf3ECH35CH"""""""""""""""""""$"""$"""$"""TCCCECCCGECEJ��N�DDJ�DDI�DDJ�DDD�3ECB4T4"ECB"DT""�r""�"""�"""R"""DDDNN�DDDNDDDGDDDCDDDBDDD�DDD�DDDBwDDBDDNSD��'DD"TDGwwww����DDDDUUUDDDgvwwwwwww~�y~�zUUUUDDDDgvfgwvvg�~ww�www�wwwUUUUDDDDwgwwwwwwwwww�www�wwgUUUTDDDtwdwtwdwtwtwtwtwtwtwtwww~�t~�t~�u��nUUUUUUUUUDwww4~~N4�tDCN�T4�CCI�TTT�UEEDwwww�w�wN~�nN��~����UUUDUUUSEUUwtwt~twt�twt�~wt�~�tUWUtUWUtUWUtUUUUUU������������""""""UTCEUUCC��uC��uE���E���E""%E""WDCC�UE4UUECE�ECE�EEE�ET4�EE4"DCT"UWUtUWUt���t���t���t���t�%"t�#"t""""""""""""""""""""""""""TD""dD""dN""tD""tG""DG""DG""�FDC�"DJ�"D�"�B""DB""DB""DB""D�""�#"t-""t/�"t/�"t"�"t"�"t"/�t"-�t""""""""""""""""""wwwDDD""Nv""DF""DF"%DE"^D�%�DRwwwwDDDDNr""DB""DB""DB""DB""DB""wwwwDDDD"/�t""�t""�t""�t""/t""/twwwtDDDD �� �������˰̻ "�+ ""  ""  D���J�8�J�D��DUD�UUUEUUTEUUDUUUCUUT3DTC03C3 �30 ˻  ̻  ��  �   �   �                           �"""۲".��""DEB"DUTDCUUT3EUU34UU3EU 33E �3D ��  ��  ��  ��  �� ə �� �� +� ""� """ """ """и�� 
��������N���N뼼D�"�T"" R"" R"� B"� �". ���˰  �  �   �   �                   "     �  �� �� �� ̻ �� �g  �'   f                                                     "   "�  ���
��ת��ڪ��z��wz��w���w���z���
���
���
��� ��� �� ��� ����ɪ�˘̻��˻ ̻� �+  ""  "   ݊� ���М�˻���̼��������������������������̻̼˻�˻�ۻ���Ԋ�X� �E E�E E�EH�UX�UE�ETE�DDE�DD        �   ˰  �˰ ��ː�̻��̻��˹@˻�D��DD��UT�EUT�UUTEUUTUUUPUUUCUUD3UTC3TC3CC3DDC4DD@DDD D�    '   rp  ''  qr  'rp srp w  w'  trp w7 w pqqppqqpp'' pwpp wpw��w��tp��wp��wp�ww�ww �"   "   "                                               ������T�M����˻� �ɚ Ț� 
��  ��  �   �   �      "  "" """�"""�  ��  ̀  �   �   �   �  "�� "˰�����"  " �"/��"/��"/���� ��� ��� ��� �˰ ̻ ""� """ """ ""/��������                     �  
�  �  �  ��  ��  ,� ,� """ """ """"" �""��""���� �  ̻  ��  ��  ��  �   �   �   �               ���������  �        �� �� �� �� ��� "��"+�""""""""""""�""�����        ��  �� ��   �   �   �  �   �   �"  "  "�� �� ���                                  �  �                                                       ��������                ����                         � � ��  ��                      ���                           �  �� ȩ ��� �̽ ��� ���ͼ���"ݻ�"�ۻ"���"����            ����ɪ��̚��̚���ɪۼ̚ۼ˚��˹"�̻"���"+��"+��"�  �� �������������}�wgw�wvr`wwv ��p ��  ��� ��� ��� �˼ ݼ� �ɘ     �� �� ��w@�ww0��C �p wwp rrp' qq'rrrw' 'rt wG     wwpwwwww�������NN��� ���7���'���r�w'wwwrwrwrrqqrqqq           �  �� �� ~w ww �w �� ww qws 'qrtqwG rss '!     wwpwwtww�������NN���p���w���7���r�w'wrrwrwrqrrqqqq                p   r      q  q  wp wp �� ��������� � �"   w   "r  w  qqp w  w  wG' srrprrqrrs'r's rqs rt wp              �   �   �   �  �   �      �   ��  ��        ���                  ����"���   � ��  "" """""""""""""���� ""��  �  �����������      ""  ""� ����� �                                         " � ̻ ��  "" """""""""""""""""""��"������������  �   "   "   "�  �� ��                                   ��� ������   �  �     �  � ��� ��  ���                           " � ̻ ��  "" """""""""""""�+  "   "   "   "�  /���/�����                    �����  ��    """ """ """"""""�"""������                        ���  ���      ,  ""  ""  "" "" �""��"" ����  "   "   "   /��������  �     ""  ""  ""  """��� ���    "   "   ""  ""  ""  ������                      ��  ��  ��                  �������������       �   �               ���    �  �� �� �� ��� ������ݽ�J���˼�ɝ�̹��̻����ͻ���ۻ��""��""-��w ���������������������������                  �  �  �� ��         �� �����ɪ��̚��̚�˼ɪ �� �������������}�wgw�wvr`wwv    �                  ���   �        �   �   �   ��� �������                    ��� ��� ����                              �                 � ���и���݊��    �   �   �   �����������                    ��  ��  ���         DD`tAGDADtDDGVwwe            UUPUVVUeeUeVVVUUeP            6tGc~E^�D�DdDDFgvP        q     qp� ��qw��'��qw�7�   qq   qqp�'�rqw�'� qw        0   3   =   M�  ��  ۸     "   "  �  �  �  �  �  �                      ���       �   �   �   ˰  ̻  ˲  +"  ""          �   �   �   �   �   "      "  "  "  "  "" ""��"" �      ������� �          ����            �   �       �   �                   �   �  �  �""""����������A������""""���������DAA""""�����HDH����H�� � a � l � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l(�(a(����������������� �  � y � � �  � � � ��� ��� � � � � � � � � � � � � ��� ��� � � � � �����y(�(����������������� = l �  � � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����((�l(=����������������    �  � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � �����((�(( ���������������� x X 5 - � � � � � � � � � ������ � � � � � � � � � � � � ������ � � �����(-(5(Xx���������������� w w x � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� � �����(�xww����������������  � w w � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � ��� �����ww�(���������������� �  + � � � � � � � � � � � �� � � ��� � � � � � � � � � � � �� � � ��� �� ����(+((����������������� ` m � W � � � � ��� � � ��� � � ��� � � � � � ��� � � ��� � � ��� � ����(W(�m(`���������������� M   a �B � � ��� � � � � � � � ��� � � � � � ��� � � � � � � � ��� ���	B�(a((M���������������� � 
 � - �C � � � ��� � � � � � ��� � ����� � ��� � � � � � ��� � ���	C�(-(� 
(����������������� � -    �DE � � � ����� ���� ��������� ����� ���� � � ��	E	D�(( (-(����������������� 5 6  X � �F � � � � � ����� � ������� � ��� � ����� � � � � ��	F ��(X((6(5���������������� x �  l � �G � � � � � � � � � � ��������� � ��� � � � � � � � � � ��	G ��l((�x���������������� w w x y�������H���������������������������������H������yxww����������������  � + w�������I�J�K�L�M�N�O � � � � � � ������� � � � � � � ��O�N�M�L�K�J�I������w(+�(���������������� , U 5  � �P���Q�R�S�T�U�V�A�A�A�W�A�A�A�W�A�A�A�A�W�A�A�A�W�A�A�A�V�U�T�S�R�Q���P(�((5(U(,���������������� +  =  U , N�P���X�Y�Z�[�\�]�]�]�^�]�]�]�^�]�]�]�]�^�]�]�]�^�]�]�]�\�[�Z�Y�X���P(N(,(U((=((+���������������� 5      = V U�P���_�`�a�b�U�U�U�c�U�U�U�c�U�U�U�U�c�U�U�U�c�U�U�U�b�a�`�_���P(U(V(=((( ((5���������������� =  U ,     !d�P���e�f�g�h�i�j�k�!�!�i�l�m�n�o�j�k�!�!�i�l�m�i�h�g�f�e���P)d((( ((,(U((=����������������     =  U , N ,�-�p�q�r�s�t�u�
�r�p�r�v�t�s�u�w�
�r�p�p�v�t�s�u�t�s�r�p�p�-(,(N(,(U((=((( ���������������� � � � � � � � � � � � � � � � � � 
 
 
 � � � � � � � � � � � �!x!y!z!{!|!}!y!~ � � � � � � � ����������������� � � � � � � � � � � � � � � � � � � 
 
 � � � � � � � � � � � �!!�!�!�!�!�!�!� � � � � � � � ����������������� ` m � �AA � � � � � � � ��� � � � � � � � � � � � � � � � ��� � � � � � �����(W(�m(`���������������� M  � �AA �@	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	@���(a((M���������������� � 
 � �AA � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � �����(-(� 
(����������������� � - � �!A � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � �� ���(( (-(����������������� 5 69�:�A�  � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���(X((6(5���������������� x � 
�;�>�' � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � ����l((�x���������������� w w x<?3 � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���yxww���������������� + � w w � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ���ww�(+���������������� � W  � � � � � � � � � � �� � �� � � � � � � � � � � � � � �� � �� � � � � � ����((W(�����������������""""������H�H�H�H�""""������HHDDH�H�""""��������H���H�����������fdffaaaDfDDFffff3333DDDDfFffFffFafFafdFfffff3333DDDDfffafffaffaffaDfffffff3333DDDDfafafFaDDFfffff3333DDDDfafDaFfDDffffff3333DDDDFaadDDdffff3333DDDDFfAFffFFFdDDffff3333DDDDffffFfffFfffFfffffffffff3333DDDD""""wwwwqqwADwqwwqw""""wwwwwAqGGGG""""wwwwwqqqAAqA""""wwwwwwqwqAAGA""""wwwwwwwwwwwwwwGwwGww""""wwwwwDAADAG""""wwwwwwGGqqqqD��������������D�����3333DDDDADAI�I��I�D����3333DDDDIIIIIIII�I�I����3333DDDDAA�A�A��ID�����3333DDDDD�I�D��������D�����3333DDDDI��I��I��I���I������3333DDDDIAI�D�DDI����3333DDDD�I�D��I��I���I�����3333DDDD""""�������AD������""""�������AD�I�""""��������AA�A""""��������DAI�A��""""������DI�I�""""�������D�I�I""""������IAD�I����""""�����������������������������I�DD����3333DDDDI�I�DI�II���I�����3333DDDD�I�I�I�ID��I����3333DDDD����������DD����3333DDDD������D���I�����������3333DDDD""""wwwwwqqwqqwqwwwwwwG""""wwwwwqwAAAGA""""wwwwwwqwqDAGAw""""wwwwwqDAwDwwGw""""wwwwwqwqwqwAwAw""""wwwwqqAqAwGwGG""""wwwwwqwADAA""""wwwwDDwGG"""$www4www4www4ww4ww4Dww4UUAUUQUUQUUQUUUDUUUU3333DDDDAADDQUEQUUUDUUUUU3333DDDDAUAUAUAUTEDUUUUU3333DDDDAUAUEEQTEUDUUUU3333DDDDUEUUQQUDUTDUUUU3333DDDDAUAUEDUQEUUDUUUU3333DDDDEAEQEQEQDEUDUUUU3333DDDDADAUDUEUQUUUDUUUU3333DDDDEUAEEQDTEUUUUU3333DDDDEUU4UUU4UUU4UU4DUU4UUU43334DDDD"""���������������""""������MM������""""�������D��""""�������DD��""""������A�A���""""�����MMDMMMM""""���������D�M""""����DD���""""������MDADM�MM��""""������D�M�M"""$���4��4��4�4��4��4������������������333DDD�DD�I�I����3333DDDDADDAII��I���I�����3333DDDD�A��D�DD����3333DDDD�AA�A�A��D�D����3333DDDD�I������D������3333DDDD������DD������3333DDDDI��I��I�I��I��D����3333DDDD�IIDIIID��I����3333DDDD��4��4��4��4�D�4���43334DDDD""""���������������������""""������II������""""������IIII""""������DI�I�""""�����IIDIIIA""""������IADD�A��""""��������I���I�������I���������������������������3333DDDD�DD�M�M����3333DDDDMDMMM�M��M�����3333DDDDM�M�M�M�M�D�����3333DDDDMAMMDMM�MM�M�M�����3333DDDDMDD���������D����3333DDDD�����M�M�DD����3333DDDDM���M���M���M���M�������3333DDDD"""wwwwwwwwqwwwwww""""wwwwwwDqq� �� �k~#1 k�#
K.X K4X K5P K6H �	CB �
CJ �CM � CO � �C< �C< �C $ �C# � C'4 � C(# �kj kr � � � � � . �K) �K9 �J� � �J� � J� � J� �J� �B� � � B� � � !B� � � "B� � �#cV u � $c^ } �%"� � � &"� �'� � �(
� �)"� � � *"� �+"� � �,*�1-"�1 ."�1!/�!0
�* �1*:� �2)��3*<�8 4*LhX 5*KXP  *Rp  *Kj  *Kj  *Kj *<j;*r <*FjF  *GjL  *Gh  *Gr3333DDDD���L��L��L��D�������3333DDDDDL��������DD�����3333DDDD���4���4��4��4D��4���43334DDDD"""wwwwwwqwwDw""""wwwwwwwGGqGqG""""wwwwwwwwGwwGwwGwwGw""""wwwwwwqwwwwDwwwwq""""wwwwqADGAwwqwq""""wwwwwwDG""""wwwwwqwDDwDq""""wwwwwwwGwwGwwwwwqwwwq""""wwwwwwGGqqqqqq"""$www4www4ww4ww4ww4ww4��D�L�L��L���333DDDALAL���D�D����3333DDDD�L��L�D�DD����3333DDDD���������������������������������A�DA�L��L���L�����3333DDDDALL�D�L�����3333DDDD��������������������������������DD�L�L����3333DDDD��4D��4L�4�L4��L4���43334DDDD�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
�<�Z�G�X�Y��U�L��Z�N�K��1�G�S�K� � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � ����������������������������������������
�
�
�
�
�
� � � � � � � � � � � � � � � � � � � � �������������������������������������������=�K�K�S�[��<�K�R�G�T�T�K� � � � � � � �@�9�1�������������������������������������������/�\�M�K�T�_��.�G�\�_�J�U�\� � � � � � �@�9�1�����������������������������������������"��<�Z�K�V�N�G�T��6�K�H�K�G�[� � � � � � �7�=�6�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%��������������������7�=�6� ���������������������������������������СơǡȡɡʡФ����������������� � � � � � �������������������������������������Сˡ̡͡ΡϡФ�����������������@�9�1� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3�T�Y�Z�G�T�Z��;�K�V�R�G�_��������������������-�N�G�T�M�K��1�U�G�R�O�K�����������������������/�J�O�Z��6�O�T�K�Y������������������������1�G�S�K��<�Z�G�Z�Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $������������������������     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %������������������������ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	                                                          	 	 
     	 	 	 	       	    	     	 	 	 	 	                                                       	    	     	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 *                                                        ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7                                                 +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @         	 	                                                 8 9 : ; < = > ? 	 @         	 	 
     	 	 	 	       	    	                                                 
     	 	 	 	       	    	     	 	 	 	 	         ! " # $                                                  ��   	 	 	 	 	         ! " # $ 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %                                                 	 % & ' ( ) 	 	 	 * +  , - . / 0 1 2 %    3 4 5 6 	 	 7 8 9 : ; < = > ? 	 @                                                ����3�4�5�6�	�	�7�8�9�:�;�<�=�>�?�	�@���������	�	�
�����	�	�	�P�                                                ���������	�	�
�����	�	�	�	�������	����	�����	�	�	�	�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                